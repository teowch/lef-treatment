<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.80168">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Curitiba" name="Torneio Regional da 1ª Região (Pré-Mirim/Petiz)" course="LCM" deadline="2024-09-09" entrystartdate="2024-09-02" entrytype="INVITATION" hostclub="Clube Curitibano" hostclub.url="https://clubecuritibano.com.br/" number="38317" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/newInterface/eventos/38317" startmethod="1" timing="AUTOMATIC" touchpad="ONESIDE" masters="F" withdrawuntil="2024-09-11" state="PR" nation="BRA" hytek.courseorder="L">
      <AGEDATE value="2024-01-01" type="YEAR" />
      <POOL name="Parque Aquático do Clube Curitibano" lanemin="1" lanemax="8" />
      <FACILITY city="Curitiba" name="Parque Aquático do Clube Curitibano" nation="BRA" state="PR" street="Avenida Presidente Getúlio Vargas, 2857" street2="Água Verde" zip="80240-040" />
      <POINTTABLE pointtableid="3017" name="AQUA Point Scoring" version="2024" />
      <QUALIFY from="2023-09-14" until="2024-09-13" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-09-14" daytime="09:10" endtime="12:24" number="1" officialmeeting="08:30" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1060" daytime="09:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1814" />
                    <RANKING order="2" place="-1" resultid="1821" />
                    <RANKING order="3" place="-1" resultid="1826" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2326" daytime="09:10" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1062" daytime="09:12" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1063" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1064" daytime="09:12" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1065" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1954" />
                    <RANKING order="2" place="2" resultid="1700" />
                    <RANKING order="3" place="3" resultid="1660" />
                    <RANKING order="4" place="4" resultid="1685" />
                    <RANKING order="5" place="5" resultid="1745" />
                    <RANKING order="6" place="6" resultid="1770" />
                    <RANKING order="7" place="7" resultid="1695" />
                    <RANKING order="8" place="8" resultid="1640" />
                    <RANKING order="9" place="9" resultid="1636" />
                    <RANKING order="10" place="10" resultid="1730" />
                    <RANKING order="11" place="-1" resultid="1650" />
                    <RANKING order="12" place="-1" resultid="1675" />
                    <RANKING order="13" place="-1" resultid="1705" />
                    <RANKING order="14" place="-1" resultid="1790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1516" />
                    <RANKING order="2" place="2" resultid="1576" />
                    <RANKING order="3" place="3" resultid="2077" />
                    <RANKING order="4" place="4" resultid="1157" />
                    <RANKING order="5" place="5" resultid="1710" />
                    <RANKING order="6" place="6" resultid="1521" />
                    <RANKING order="7" place="7" resultid="1665" />
                    <RANKING order="8" place="7" resultid="1912" />
                    <RANKING order="9" place="9" resultid="1621" />
                    <RANKING order="10" place="10" resultid="1581" />
                    <RANKING order="11" place="11" resultid="1551" />
                    <RANKING order="12" place="12" resultid="1968" />
                    <RANKING order="13" place="13" resultid="1785" />
                    <RANKING order="14" place="-1" resultid="1596" />
                    <RANKING order="15" place="-1" resultid="1611" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2327" daytime="09:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2328" daytime="09:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2329" daytime="09:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2330" daytime="09:30" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1067" daytime="09:34" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1068" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1645" />
                    <RANKING order="2" place="2" resultid="2063" />
                    <RANKING order="3" place="3" resultid="1236" />
                    <RANKING order="4" place="4" resultid="1795" />
                    <RANKING order="5" place="5" resultid="1680" />
                    <RANKING order="6" place="6" resultid="1720" />
                    <RANKING order="7" place="7" resultid="1735" />
                    <RANKING order="8" place="8" resultid="1740" />
                    <RANKING order="9" place="9" resultid="1755" />
                    <RANKING order="10" place="10" resultid="1775" />
                    <RANKING order="11" place="11" resultid="1780" />
                    <RANKING order="12" place="12" resultid="1765" />
                    <RANKING order="13" place="-1" resultid="1631" />
                    <RANKING order="14" place="-1" resultid="1690" />
                    <RANKING order="15" place="-1" resultid="1725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1591" />
                    <RANKING order="2" place="2" resultid="1917" />
                    <RANKING order="3" place="3" resultid="1506" />
                    <RANKING order="4" place="4" resultid="1670" />
                    <RANKING order="5" place="5" resultid="1536" />
                    <RANKING order="6" place="6" resultid="1715" />
                    <RANKING order="7" place="7" resultid="1531" />
                    <RANKING order="8" place="8" resultid="2024" />
                    <RANKING order="9" place="9" resultid="1526" />
                    <RANKING order="10" place="10" resultid="1232" />
                    <RANKING order="11" place="11" resultid="1586" />
                    <RANKING order="12" place="12" resultid="1566" />
                    <RANKING order="13" place="13" resultid="1800" />
                    <RANKING order="14" place="14" resultid="1655" />
                    <RANKING order="15" place="15" resultid="1561" />
                    <RANKING order="16" place="16" resultid="2111" />
                    <RANKING order="17" place="-1" resultid="1571" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2331" daytime="09:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2332" daytime="09:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2333" daytime="09:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2334" daytime="09:52" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1070" daytime="09:56" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1071" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2014" />
                    <RANKING order="2" place="2" resultid="1380" />
                    <RANKING order="3" place="3" resultid="1886" />
                    <RANKING order="4" place="4" resultid="1375" />
                    <RANKING order="5" place="5" resultid="1390" />
                    <RANKING order="6" place="6" resultid="1999" />
                    <RANKING order="7" place="7" resultid="1432" />
                    <RANKING order="8" place="8" resultid="1606" />
                    <RANKING order="9" place="9" resultid="1409" />
                    <RANKING order="10" place="-1" resultid="1556" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1305" />
                    <RANKING order="2" place="2" resultid="1360" />
                    <RANKING order="3" place="3" resultid="1395" />
                    <RANKING order="4" place="4" resultid="1340" />
                    <RANKING order="5" place="5" resultid="1750" />
                    <RANKING order="6" place="6" resultid="2106" />
                    <RANKING order="7" place="7" resultid="1345" />
                    <RANKING order="8" place="8" resultid="1385" />
                    <RANKING order="9" place="9" resultid="2009" />
                    <RANKING order="10" place="10" resultid="1197" />
                    <RANKING order="11" place="11" resultid="1335" />
                    <RANKING order="12" place="12" resultid="1926" />
                    <RANKING order="13" place="13" resultid="1989" />
                    <RANKING order="14" place="14" resultid="1975" />
                    <RANKING order="15" place="15" resultid="1501" />
                    <RANKING order="16" place="-1" resultid="1601" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2335" daytime="09:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2336" daytime="10:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2337" daytime="10:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2338" daytime="10:12" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1073" daytime="10:16" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1074" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1437" />
                    <RANKING order="2" place="2" resultid="2043" />
                    <RANKING order="3" place="3" resultid="1462" />
                    <RANKING order="4" place="4" resultid="1447" />
                    <RANKING order="5" place="5" resultid="1832" />
                    <RANKING order="6" place="6" resultid="1252" />
                    <RANKING order="7" place="7" resultid="1616" />
                    <RANKING order="8" place="8" resultid="2058" />
                    <RANKING order="9" place="9" resultid="1476" />
                    <RANKING order="10" place="10" resultid="1400" />
                    <RANKING order="11" place="11" resultid="1903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1285" />
                    <RANKING order="2" place="2" resultid="1325" />
                    <RANKING order="3" place="3" resultid="1350" />
                    <RANKING order="4" place="4" resultid="1937" />
                    <RANKING order="5" place="5" resultid="1295" />
                    <RANKING order="6" place="6" resultid="1355" />
                    <RANKING order="7" place="7" resultid="1310" />
                    <RANKING order="8" place="8" resultid="1320" />
                    <RANKING order="9" place="9" resultid="2004" />
                    <RANKING order="10" place="10" resultid="2068" />
                    <RANKING order="11" place="-1" resultid="1365" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2339" daytime="10:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2340" daytime="10:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2341" daytime="10:26" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1076" daytime="10:30" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1077" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1827" />
                    <RANKING order="2" place="2" resultid="1262" />
                    <RANKING order="3" place="3" resultid="1815" />
                    <RANKING order="4" place="4" resultid="1869" />
                    <RANKING order="5" place="5" resultid="1865" />
                    <RANKING order="6" place="6" resultid="1819" />
                    <RANKING order="7" place="-1" resultid="1822" />
                    <RANKING order="8" place="-1" resultid="1843" />
                    <RANKING order="9" place="-1" resultid="1850" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2342" daytime="10:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2343" daytime="10:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1078" daytime="10:36" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1079" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1271" />
                    <RANKING order="2" place="2" resultid="1857" />
                    <RANKING order="3" place="3" resultid="1847" />
                    <RANKING order="4" place="4" resultid="2141" />
                    <RANKING order="5" place="5" resultid="1861" />
                    <RANKING order="6" place="-1" resultid="1810" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2344" daytime="10:36" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1080" daytime="10:40" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1081" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1684" />
                    <RANKING order="2" place="2" resultid="1172" />
                    <RANKING order="3" place="3" resultid="1220" />
                    <RANKING order="4" place="4" resultid="1769" />
                    <RANKING order="5" place="5" resultid="1964" />
                    <RANKING order="6" place="6" resultid="1635" />
                    <RANKING order="7" place="7" resultid="1744" />
                    <RANKING order="8" place="-1" resultid="1649" />
                    <RANKING order="9" place="-1" resultid="1674" />
                    <RANKING order="10" place="-1" resultid="1704" />
                    <RANKING order="11" place="-1" resultid="1789" />
                    <RANKING order="12" place="-1" resultid="1836" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1994" />
                    <RANKING order="2" place="2" resultid="2129" />
                    <RANKING order="3" place="3" resultid="1620" />
                    <RANKING order="4" place="4" resultid="2134" />
                    <RANKING order="5" place="5" resultid="1162" />
                    <RANKING order="6" place="6" resultid="2124" />
                    <RANKING order="7" place="7" resultid="2082" />
                    <RANKING order="8" place="8" resultid="1267" />
                    <RANKING order="9" place="9" resultid="1959" />
                    <RANKING order="10" place="10" resultid="1179" />
                    <RANKING order="11" place="11" resultid="1550" />
                    <RANKING order="12" place="-1" resultid="1595" />
                    <RANKING order="13" place="-1" resultid="1610" />
                    <RANKING order="14" place="-1" resultid="1626" />
                    <RANKING order="15" place="-1" resultid="1784" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2345" daytime="10:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2346" daytime="10:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2347" daytime="10:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2348" daytime="10:48" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1083" daytime="10:50" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1084" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1739" />
                    <RANKING order="2" place="2" resultid="2062" />
                    <RANKING order="3" place="3" resultid="1754" />
                    <RANKING order="4" place="4" resultid="1908" />
                    <RANKING order="5" place="5" resultid="1719" />
                    <RANKING order="6" place="6" resultid="1774" />
                    <RANKING order="7" place="7" resultid="1779" />
                    <RANKING order="8" place="-1" resultid="1734" />
                    <RANKING order="9" place="-1" resultid="1630" />
                    <RANKING order="10" place="-1" resultid="1724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1535" />
                    <RANKING order="2" place="2" resultid="2023" />
                    <RANKING order="3" place="3" resultid="1176" />
                    <RANKING order="4" place="4" resultid="1560" />
                    <RANKING order="5" place="5" resultid="1951" />
                    <RANKING order="6" place="6" resultid="1565" />
                    <RANKING order="7" place="7" resultid="1211" />
                    <RANKING order="8" place="8" resultid="2096" />
                    <RANKING order="9" place="9" resultid="2101" />
                    <RANKING order="10" place="10" resultid="1714" />
                    <RANKING order="11" place="11" resultid="1799" />
                    <RANKING order="12" place="12" resultid="2038" />
                    <RANKING order="13" place="13" resultid="1183" />
                    <RANKING order="14" place="14" resultid="1546" />
                    <RANKING order="15" place="15" resultid="2019" />
                    <RANKING order="16" place="16" resultid="2087" />
                    <RANKING order="17" place="17" resultid="1541" />
                    <RANKING order="18" place="18" resultid="1654" />
                    <RANKING order="19" place="19" resultid="1570" />
                    <RANKING order="20" place="20" resultid="1231" />
                    <RANKING order="21" place="21" resultid="2110" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2349" daytime="10:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2350" daytime="10:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2351" daytime="10:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2352" daytime="10:56" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1086" daytime="11:00" gender="F" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1087" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1760" />
                    <RANKING order="2" place="2" resultid="1885" />
                    <RANKING order="3" place="3" resultid="2013" />
                    <RANKING order="4" place="4" resultid="1389" />
                    <RANKING order="5" place="5" resultid="2148" />
                    <RANKING order="6" place="6" resultid="1491" />
                    <RANKING order="7" place="7" resultid="1898" />
                    <RANKING order="8" place="8" resultid="1245" />
                    <RANKING order="9" place="9" resultid="1202" />
                    <RANKING order="10" place="10" resultid="1998" />
                    <RANKING order="11" place="11" resultid="2048" />
                    <RANKING order="12" place="12" resultid="1431" />
                    <RANKING order="13" place="13" resultid="1169" />
                    <RANKING order="14" place="14" resultid="2028" />
                    <RANKING order="15" place="15" resultid="1511" />
                    <RANKING order="16" place="16" resultid="1942" />
                    <RANKING order="17" place="17" resultid="1605" />
                    <RANKING order="18" place="18" resultid="1894" />
                    <RANKING order="19" place="19" resultid="1408" />
                    <RANKING order="20" place="20" resultid="1980" />
                    <RANKING order="21" place="21" resultid="1224" />
                    <RANKING order="22" place="22" resultid="2072" />
                    <RANKING order="23" place="-1" resultid="1422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1457" />
                    <RANKING order="2" place="2" resultid="1300" />
                    <RANKING order="3" place="3" resultid="1394" />
                    <RANKING order="4" place="4" resultid="1304" />
                    <RANKING order="5" place="5" resultid="1749" />
                    <RANKING order="6" place="6" resultid="1600" />
                    <RANKING order="7" place="7" resultid="1384" />
                    <RANKING order="8" place="8" resultid="2008" />
                    <RANKING order="9" place="9" resultid="1988" />
                    <RANKING order="10" place="10" resultid="1256" />
                    <RANKING order="11" place="11" resultid="1925" />
                    <RANKING order="12" place="12" resultid="1881" />
                    <RANKING order="13" place="13" resultid="1150" />
                    <RANKING order="14" place="14" resultid="1974" />
                    <RANKING order="15" place="15" resultid="1216" />
                    <RANKING order="16" place="16" resultid="1442" />
                    <RANKING order="17" place="17" resultid="1259" />
                    <RANKING order="18" place="18" resultid="1500" />
                    <RANKING order="19" place="19" resultid="2119" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2353" daytime="11:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2354" daytime="11:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2355" daytime="11:08" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2356" daytime="11:12" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2357" daytime="11:14" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2358" daytime="11:16" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1089" daytime="11:20" gender="M" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1090" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1467" />
                    <RANKING order="2" place="2" resultid="1153" />
                    <RANKING order="3" place="3" resultid="1251" />
                    <RANKING order="4" place="4" resultid="2042" />
                    <RANKING order="5" place="5" resultid="1370" />
                    <RANKING order="6" place="6" resultid="2057" />
                    <RANKING order="7" place="7" resultid="1615" />
                    <RANKING order="8" place="8" resultid="1831" />
                    <RANKING order="9" place="9" resultid="1481" />
                    <RANKING order="10" place="10" resultid="1902" />
                    <RANKING order="11" place="11" resultid="1414" />
                    <RANKING order="12" place="12" resultid="2053" />
                    <RANKING order="13" place="13" resultid="1427" />
                    <RANKING order="14" place="14" resultid="2033" />
                    <RANKING order="15" place="15" resultid="1486" />
                    <RANKING order="16" place="16" resultid="1475" />
                    <RANKING order="17" place="17" resultid="1946" />
                    <RANKING order="18" place="18" resultid="2116" />
                    <RANKING order="19" place="19" resultid="1276" />
                    <RANKING order="20" place="20" resultid="1890" />
                    <RANKING order="21" place="21" resultid="1840" />
                    <RANKING order="22" place="-1" resultid="1928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1324" />
                    <RANKING order="2" place="2" resultid="1315" />
                    <RANKING order="3" place="3" resultid="1330" />
                    <RANKING order="4" place="4" resultid="1349" />
                    <RANKING order="5" place="5" resultid="1496" />
                    <RANKING order="6" place="6" resultid="1290" />
                    <RANKING order="7" place="7" resultid="1936" />
                    <RANKING order="8" place="8" resultid="1309" />
                    <RANKING order="9" place="9" resultid="1189" />
                    <RANKING order="10" place="10" resultid="1206" />
                    <RANKING order="11" place="11" resultid="1249" />
                    <RANKING order="12" place="12" resultid="1192" />
                    <RANKING order="13" place="13" resultid="1280" />
                    <RANKING order="14" place="14" resultid="1240" />
                    <RANKING order="15" place="15" resultid="1319" />
                    <RANKING order="16" place="16" resultid="1932" />
                    <RANKING order="17" place="17" resultid="1404" />
                    <RANKING order="18" place="18" resultid="2091" />
                    <RANKING order="19" place="19" resultid="2138" />
                    <RANKING order="20" place="20" resultid="1452" />
                    <RANKING order="21" place="21" resultid="1227" />
                    <RANKING order="22" place="-1" resultid="1921" />
                    <RANKING order="23" place="-1" resultid="1984" />
                    <RANKING order="24" place="-1" resultid="1364" />
                    <RANKING order="25" place="-1" resultid="1471" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2359" daytime="11:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2360" daytime="11:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2361" daytime="11:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2362" daytime="11:28" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2363" daytime="11:32" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2364" daytime="11:34" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1092" daytime="11:36" gender="F" number="13" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1093" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1953" />
                    <RANKING order="2" place="2" resultid="1699" />
                    <RANKING order="3" place="3" resultid="1659" />
                    <RANKING order="4" place="4" resultid="1694" />
                    <RANKING order="5" place="5" resultid="1963" />
                    <RANKING order="6" place="6" resultid="1639" />
                    <RANKING order="7" place="7" resultid="1729" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1993" />
                    <RANKING order="2" place="2" resultid="1515" />
                    <RANKING order="3" place="3" resultid="2076" />
                    <RANKING order="4" place="4" resultid="1709" />
                    <RANKING order="5" place="5" resultid="1575" />
                    <RANKING order="6" place="6" resultid="1520" />
                    <RANKING order="7" place="7" resultid="1664" />
                    <RANKING order="8" place="8" resultid="2128" />
                    <RANKING order="9" place="9" resultid="1156" />
                    <RANKING order="10" place="10" resultid="1958" />
                    <RANKING order="11" place="11" resultid="2081" />
                    <RANKING order="12" place="12" resultid="2133" />
                    <RANKING order="13" place="13" resultid="1266" />
                    <RANKING order="14" place="14" resultid="2123" />
                    <RANKING order="15" place="15" resultid="1580" />
                    <RANKING order="16" place="16" resultid="1161" />
                    <RANKING order="17" place="-1" resultid="1625" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2365" daytime="11:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2366" daytime="11:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2367" daytime="11:42" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1095" daytime="11:44" gender="M" number="14" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1096" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1644" />
                    <RANKING order="2" place="2" resultid="1689" />
                    <RANKING order="3" place="3" resultid="1794" />
                    <RANKING order="4" place="4" resultid="1679" />
                    <RANKING order="5" place="5" resultid="1907" />
                    <RANKING order="6" place="6" resultid="1764" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1505" />
                    <RANKING order="2" place="2" resultid="1590" />
                    <RANKING order="3" place="3" resultid="1525" />
                    <RANKING order="4" place="4" resultid="1530" />
                    <RANKING order="5" place="5" resultid="1916" />
                    <RANKING order="6" place="6" resultid="1669" />
                    <RANKING order="7" place="7" resultid="1585" />
                    <RANKING order="8" place="8" resultid="2018" />
                    <RANKING order="9" place="9" resultid="1175" />
                    <RANKING order="10" place="10" resultid="1950" />
                    <RANKING order="11" place="11" resultid="1210" />
                    <RANKING order="12" place="12" resultid="2037" />
                    <RANKING order="13" place="13" resultid="1545" />
                    <RANKING order="14" place="14" resultid="2095" />
                    <RANKING order="15" place="15" resultid="2086" />
                    <RANKING order="16" place="16" resultid="2100" />
                    <RANKING order="17" place="17" resultid="1540" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2368" daytime="11:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2369" daytime="11:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2370" daytime="11:48" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1098" daytime="11:52" gender="F" number="15" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1099" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1759" />
                    <RANKING order="2" place="2" resultid="1379" />
                    <RANKING order="3" place="3" resultid="1374" />
                    <RANKING order="4" place="4" resultid="1490" />
                    <RANKING order="5" place="5" resultid="1897" />
                    <RANKING order="6" place="6" resultid="2147" />
                    <RANKING order="7" place="7" resultid="1555" />
                    <RANKING order="8" place="8" resultid="1244" />
                    <RANKING order="9" place="9" resultid="1201" />
                    <RANKING order="10" place="10" resultid="1510" />
                    <RANKING order="11" place="11" resultid="1941" />
                    <RANKING order="12" place="12" resultid="1979" />
                    <RANKING order="13" place="13" resultid="1893" />
                    <RANKING order="14" place="-1" resultid="2047" />
                    <RANKING order="15" place="-1" resultid="1421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1456" />
                    <RANKING order="2" place="2" resultid="2105" />
                    <RANKING order="3" place="3" resultid="1299" />
                    <RANKING order="4" place="4" resultid="1359" />
                    <RANKING order="5" place="5" resultid="1339" />
                    <RANKING order="6" place="6" resultid="1334" />
                    <RANKING order="7" place="7" resultid="1196" />
                    <RANKING order="8" place="8" resultid="1255" />
                    <RANKING order="9" place="9" resultid="1880" />
                    <RANKING order="10" place="10" resultid="1215" />
                    <RANKING order="11" place="11" resultid="1441" />
                    <RANKING order="12" place="-1" resultid="1344" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2371" daytime="11:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2372" daytime="11:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2373" daytime="11:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2374" daytime="11:58" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1101" daytime="12:00" gender="M" number="16" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1102" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1152" />
                    <RANKING order="2" place="2" resultid="1369" />
                    <RANKING order="3" place="3" resultid="1466" />
                    <RANKING order="4" place="4" resultid="1461" />
                    <RANKING order="5" place="5" resultid="1399" />
                    <RANKING order="6" place="6" resultid="1413" />
                    <RANKING order="7" place="7" resultid="1446" />
                    <RANKING order="8" place="8" resultid="1436" />
                    <RANKING order="9" place="9" resultid="1426" />
                    <RANKING order="10" place="10" resultid="1485" />
                    <RANKING order="11" place="11" resultid="1945" />
                    <RANKING order="12" place="12" resultid="2032" />
                    <RANKING order="13" place="13" resultid="2052" />
                    <RANKING order="14" place="14" resultid="1275" />
                    <RANKING order="15" place="15" resultid="2115" />
                    <RANKING order="16" place="-1" resultid="1480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1284" />
                    <RANKING order="2" place="2" resultid="1354" />
                    <RANKING order="3" place="3" resultid="1294" />
                    <RANKING order="4" place="4" resultid="1314" />
                    <RANKING order="5" place="5" resultid="2003" />
                    <RANKING order="6" place="6" resultid="1495" />
                    <RANKING order="7" place="7" resultid="1248" />
                    <RANKING order="8" place="8" resultid="1983" />
                    <RANKING order="9" place="9" resultid="1289" />
                    <RANKING order="10" place="10" resultid="1329" />
                    <RANKING order="11" place="11" resultid="1205" />
                    <RANKING order="12" place="12" resultid="2067" />
                    <RANKING order="13" place="13" resultid="1188" />
                    <RANKING order="14" place="14" resultid="1451" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2375" daytime="12:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2376" daytime="12:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2377" daytime="12:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2378" daytime="12:06" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-09-14" daytime="15:40" endtime="19:38" number="2" officialmeeting="15:00" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1104" daytime="15:40" gender="F" number="17" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1105" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1264" />
                    <RANKING order="2" place="2" resultid="1817" />
                    <RANKING order="3" place="3" resultid="1829" />
                    <RANKING order="4" place="4" resultid="1871" />
                    <RANKING order="5" place="5" resultid="1867" />
                    <RANKING order="6" place="-1" resultid="1808" />
                    <RANKING order="7" place="-1" resultid="1824" />
                    <RANKING order="8" place="-1" resultid="1845" />
                    <RANKING order="9" place="-1" resultid="1852" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2379" daytime="15:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2380" daytime="15:42" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1106" daytime="15:46" gender="M" number="18" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1107" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1273" />
                    <RANKING order="2" place="2" resultid="1877" />
                    <RANKING order="3" place="3" resultid="1812" />
                    <RANKING order="4" place="4" resultid="1863" />
                    <RANKING order="5" place="-1" resultid="1805" />
                    <RANKING order="6" place="-1" resultid="1855" />
                    <RANKING order="7" place="-1" resultid="1859" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2381" daytime="15:46" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1108" daytime="15:48" gender="F" number="19" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1109" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1956" />
                    <RANKING order="2" place="2" resultid="1687" />
                    <RANKING order="3" place="3" resultid="1662" />
                    <RANKING order="4" place="4" resultid="1702" />
                    <RANKING order="5" place="5" resultid="1966" />
                    <RANKING order="6" place="6" resultid="1642" />
                    <RANKING order="7" place="7" resultid="1697" />
                    <RANKING order="8" place="8" resultid="1637" />
                    <RANKING order="9" place="9" resultid="1747" />
                    <RANKING order="10" place="10" resultid="1732" />
                    <RANKING order="11" place="-1" resultid="1772" />
                    <RANKING order="12" place="-1" resultid="1677" />
                    <RANKING order="13" place="-1" resultid="1707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1110" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1996" />
                    <RANKING order="2" place="2" resultid="1518" />
                    <RANKING order="3" place="3" resultid="2079" />
                    <RANKING order="4" place="4" resultid="1578" />
                    <RANKING order="5" place="5" resultid="1712" />
                    <RANKING order="6" place="6" resultid="1523" />
                    <RANKING order="7" place="7" resultid="1623" />
                    <RANKING order="8" place="8" resultid="1972" />
                    <RANKING order="9" place="9" resultid="1961" />
                    <RANKING order="10" place="10" resultid="1667" />
                    <RANKING order="11" place="-1" resultid="1583" />
                    <RANKING order="12" place="-1" resultid="1613" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2382" daytime="15:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2383" daytime="15:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2384" daytime="16:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2385" daytime="16:06" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1111" daytime="16:12" gender="M" number="20" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1112" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1646" />
                    <RANKING order="2" place="2" resultid="2064" />
                    <RANKING order="3" place="3" resultid="1797" />
                    <RANKING order="4" place="4" resultid="1681" />
                    <RANKING order="5" place="5" resultid="1722" />
                    <RANKING order="6" place="6" resultid="1757" />
                    <RANKING order="7" place="7" resultid="1737" />
                    <RANKING order="8" place="-1" resultid="1632" />
                    <RANKING order="9" place="-1" resultid="1692" />
                    <RANKING order="10" place="-1" resultid="1726" />
                    <RANKING order="11" place="-1" resultid="1741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1538" />
                    <RANKING order="2" place="2" resultid="1507" />
                    <RANKING order="3" place="3" resultid="1527" />
                    <RANKING order="4" place="4" resultid="1671" />
                    <RANKING order="5" place="5" resultid="1533" />
                    <RANKING order="6" place="6" resultid="1592" />
                    <RANKING order="7" place="7" resultid="1587" />
                    <RANKING order="8" place="8" resultid="1717" />
                    <RANKING order="9" place="9" resultid="2040" />
                    <RANKING order="10" place="10" resultid="1568" />
                    <RANKING order="11" place="11" resultid="2020" />
                    <RANKING order="12" place="12" resultid="2097" />
                    <RANKING order="13" place="13" resultid="1562" />
                    <RANKING order="14" place="14" resultid="1801" />
                    <RANKING order="15" place="15" resultid="2088" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2386" daytime="16:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2387" daytime="16:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2388" daytime="16:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2389" daytime="16:32" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1114" daytime="16:36" gender="F" number="21" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1115" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1888" />
                    <RANKING order="2" place="2" resultid="2015" />
                    <RANKING order="3" place="3" resultid="1761" />
                    <RANKING order="4" place="4" resultid="1381" />
                    <RANKING order="5" place="5" resultid="1391" />
                    <RANKING order="6" place="6" resultid="1424" />
                    <RANKING order="7" place="7" resultid="2001" />
                    <RANKING order="8" place="8" resultid="1434" />
                    <RANKING order="9" place="9" resultid="1419" />
                    <RANKING order="10" place="10" resultid="1377" />
                    <RANKING order="11" place="11" resultid="1493" />
                    <RANKING order="12" place="12" resultid="1513" />
                    <RANKING order="13" place="13" resultid="1558" />
                    <RANKING order="14" place="14" resultid="2050" />
                    <RANKING order="15" place="15" resultid="1607" />
                    <RANKING order="16" place="16" resultid="1410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1307" />
                    <RANKING order="2" place="2" resultid="1459" />
                    <RANKING order="3" place="3" resultid="1397" />
                    <RANKING order="4" place="4" resultid="1302" />
                    <RANKING order="5" place="5" resultid="1341" />
                    <RANKING order="6" place="6" resultid="1751" />
                    <RANKING order="7" place="7" resultid="1387" />
                    <RANKING order="8" place="8" resultid="1361" />
                    <RANKING order="9" place="9" resultid="1257" />
                    <RANKING order="10" place="10" resultid="2011" />
                    <RANKING order="11" place="11" resultid="1443" />
                    <RANKING order="12" place="-1" resultid="1346" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2390" daytime="16:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2391" daytime="16:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2392" daytime="16:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2393" daytime="17:02" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1117" daytime="17:10" gender="M" number="22" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1118" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1438" />
                    <RANKING order="2" place="2" resultid="1469" />
                    <RANKING order="3" place="3" resultid="2060" />
                    <RANKING order="4" place="4" resultid="1463" />
                    <RANKING order="5" place="5" resultid="1372" />
                    <RANKING order="6" place="6" resultid="1448" />
                    <RANKING order="7" place="7" resultid="2044" />
                    <RANKING order="8" place="8" resultid="1833" />
                    <RANKING order="9" place="9" resultid="1618" />
                    <RANKING order="10" place="10" resultid="1488" />
                    <RANKING order="11" place="11" resultid="1428" />
                    <RANKING order="12" place="12" resultid="1477" />
                    <RANKING order="13" place="13" resultid="2035" />
                    <RANKING order="14" place="14" resultid="1401" />
                    <RANKING order="15" place="15" resultid="1948" />
                    <RANKING order="16" place="-1" resultid="1416" />
                    <RANKING order="17" place="-1" resultid="1483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1332" />
                    <RANKING order="2" place="2" resultid="1326" />
                    <RANKING order="3" place="3" resultid="1317" />
                    <RANKING order="4" place="4" resultid="1351" />
                    <RANKING order="5" place="5" resultid="1985" />
                    <RANKING order="6" place="6" resultid="1497" />
                    <RANKING order="7" place="7" resultid="1356" />
                    <RANKING order="8" place="8" resultid="1292" />
                    <RANKING order="9" place="9" resultid="1312" />
                    <RANKING order="10" place="10" resultid="2069" />
                    <RANKING order="11" place="-1" resultid="1287" />
                    <RANKING order="12" place="-1" resultid="1297" />
                    <RANKING order="13" place="-1" resultid="1321" />
                    <RANKING order="14" place="-1" resultid="1366" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2394" daytime="17:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2395" daytime="17:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2396" daytime="17:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2397" daytime="17:34" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1120" daytime="17:40" gender="F" number="23" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1121" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1263" />
                    <RANKING order="2" place="2" resultid="1828" />
                    <RANKING order="3" place="3" resultid="1816" />
                    <RANKING order="4" place="4" resultid="1866" />
                    <RANKING order="5" place="5" resultid="1870" />
                    <RANKING order="6" place="-1" resultid="1807" />
                    <RANKING order="7" place="-1" resultid="1823" />
                    <RANKING order="8" place="-1" resultid="1844" />
                    <RANKING order="9" place="-1" resultid="1851" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2398" daytime="17:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2399" daytime="17:42" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1122" daytime="17:46" gender="M" number="24" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1123" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1272" />
                    <RANKING order="2" place="2" resultid="1876" />
                    <RANKING order="3" place="3" resultid="2142" />
                    <RANKING order="4" place="4" resultid="1811" />
                    <RANKING order="5" place="5" resultid="1862" />
                    <RANKING order="6" place="6" resultid="1858" />
                    <RANKING order="7" place="-1" resultid="1804" />
                    <RANKING order="8" place="-1" resultid="1848" />
                    <RANKING order="9" place="-1" resultid="1854" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2400" daytime="17:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2401" daytime="17:48" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1124" daytime="17:50" gender="F" number="25" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1125" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1686" />
                    <RANKING order="2" place="2" resultid="1965" />
                    <RANKING order="3" place="3" resultid="1701" />
                    <RANKING order="4" place="4" resultid="1838" />
                    <RANKING order="5" place="5" resultid="1222" />
                    <RANKING order="6" place="6" resultid="1696" />
                    <RANKING order="7" place="7" resultid="1641" />
                    <RANKING order="8" place="8" resultid="1731" />
                    <RANKING order="9" place="-1" resultid="1652" />
                    <RANKING order="10" place="-1" resultid="1676" />
                    <RANKING order="11" place="-1" resultid="1792" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2078" />
                    <RANKING order="2" place="2" resultid="2131" />
                    <RANKING order="3" place="3" resultid="2084" />
                    <RANKING order="4" place="4" resultid="2136" />
                    <RANKING order="5" place="5" resultid="1159" />
                    <RANKING order="6" place="6" resultid="1666" />
                    <RANKING order="7" place="7" resultid="1622" />
                    <RANKING order="8" place="8" resultid="1522" />
                    <RANKING order="9" place="9" resultid="1914" />
                    <RANKING order="10" place="10" resultid="1164" />
                    <RANKING order="11" place="11" resultid="1181" />
                    <RANKING order="12" place="12" resultid="1969" />
                    <RANKING order="13" place="13" resultid="2126" />
                    <RANKING order="14" place="14" resultid="1269" />
                    <RANKING order="15" place="15" resultid="1553" />
                    <RANKING order="16" place="-1" resultid="1598" />
                    <RANKING order="17" place="-1" resultid="1612" />
                    <RANKING order="18" place="-1" resultid="1628" />
                    <RANKING order="19" place="-1" resultid="1787" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2402" daytime="17:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2403" daytime="17:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2404" daytime="17:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2405" daytime="18:00" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1127" daytime="18:02" gender="M" number="26" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1128" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1237" />
                    <RANKING order="2" place="2" resultid="1796" />
                    <RANKING order="3" place="3" resultid="1691" />
                    <RANKING order="4" place="4" resultid="1873" />
                    <RANKING order="5" place="5" resultid="1909" />
                    <RANKING order="6" place="6" resultid="1721" />
                    <RANKING order="7" place="7" resultid="1736" />
                    <RANKING order="8" place="8" resultid="1756" />
                    <RANKING order="9" place="9" resultid="2144" />
                    <RANKING order="10" place="10" resultid="2155" />
                    <RANKING order="11" place="11" resultid="1776" />
                    <RANKING order="12" place="12" resultid="1781" />
                    <RANKING order="13" place="13" resultid="2152" />
                    <RANKING order="14" place="14" resultid="2161" />
                    <RANKING order="15" place="15" resultid="1766" />
                    <RANKING order="16" place="16" resultid="2158" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1918" />
                    <RANKING order="2" place="2" resultid="1532" />
                    <RANKING order="3" place="3" resultid="1716" />
                    <RANKING order="4" place="4" resultid="1166" />
                    <RANKING order="5" place="5" resultid="1567" />
                    <RANKING order="6" place="6" resultid="1537" />
                    <RANKING order="7" place="7" resultid="1212" />
                    <RANKING order="8" place="8" resultid="2025" />
                    <RANKING order="9" place="9" resultid="2102" />
                    <RANKING order="10" place="10" resultid="2039" />
                    <RANKING order="11" place="11" resultid="1233" />
                    <RANKING order="12" place="12" resultid="1656" />
                    <RANKING order="13" place="13" resultid="1547" />
                    <RANKING order="14" place="14" resultid="1542" />
                    <RANKING order="15" place="15" resultid="1184" />
                    <RANKING order="16" place="16" resultid="1572" />
                    <RANKING order="17" place="17" resultid="2112" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2406" daytime="18:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2407" daytime="18:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2408" daytime="18:08" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2409" daytime="18:12" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2410" daytime="18:14" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1130" daytime="18:16" gender="F" number="27" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1131" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1418" />
                    <RANKING order="2" place="2" resultid="1423" />
                    <RANKING order="3" place="3" resultid="1376" />
                    <RANKING order="4" place="4" resultid="1887" />
                    <RANKING order="5" place="5" resultid="2000" />
                    <RANKING order="6" place="6" resultid="1899" />
                    <RANKING order="7" place="7" resultid="1246" />
                    <RANKING order="8" place="8" resultid="1433" />
                    <RANKING order="9" place="9" resultid="2049" />
                    <RANKING order="10" place="10" resultid="1203" />
                    <RANKING order="11" place="11" resultid="2029" />
                    <RANKING order="12" place="12" resultid="1512" />
                    <RANKING order="13" place="13" resultid="2149" />
                    <RANKING order="14" place="14" resultid="1895" />
                    <RANKING order="15" place="15" resultid="2073" />
                    <RANKING order="16" place="-1" resultid="1492" />
                    <RANKING order="17" place="-1" resultid="1557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1132" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1458" />
                    <RANKING order="2" place="2" resultid="1602" />
                    <RANKING order="3" place="3" resultid="1301" />
                    <RANKING order="4" place="4" resultid="1306" />
                    <RANKING order="5" place="5" resultid="1396" />
                    <RANKING order="6" place="6" resultid="1386" />
                    <RANKING order="7" place="7" resultid="2010" />
                    <RANKING order="8" place="8" resultid="1990" />
                    <RANKING order="9" place="9" resultid="1198" />
                    <RANKING order="10" place="10" resultid="2107" />
                    <RANKING order="11" place="11" resultid="1882" />
                    <RANKING order="12" place="12" resultid="1976" />
                    <RANKING order="13" place="13" resultid="1217" />
                    <RANKING order="14" place="14" resultid="1336" />
                    <RANKING order="15" place="15" resultid="1502" />
                    <RANKING order="16" place="16" resultid="1260" />
                    <RANKING order="17" place="-1" resultid="2120" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2411" daytime="18:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2412" daytime="18:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2413" daytime="18:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2414" daytime="18:28" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2415" daytime="18:32" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1133" daytime="18:34" gender="M" number="28" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1134" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1154" />
                    <RANKING order="2" place="2" resultid="1468" />
                    <RANKING order="3" place="3" resultid="1617" />
                    <RANKING order="4" place="4" resultid="1371" />
                    <RANKING order="5" place="5" resultid="2059" />
                    <RANKING order="6" place="6" resultid="1904" />
                    <RANKING order="7" place="7" resultid="2034" />
                    <RANKING order="8" place="8" resultid="1487" />
                    <RANKING order="9" place="9" resultid="2054" />
                    <RANKING order="10" place="10" resultid="1277" />
                    <RANKING order="11" place="11" resultid="1947" />
                    <RANKING order="12" place="12" resultid="1929" />
                    <RANKING order="13" place="-1" resultid="1415" />
                    <RANKING order="14" place="-1" resultid="1482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1938" />
                    <RANKING order="2" place="2" resultid="1286" />
                    <RANKING order="3" place="3" resultid="1207" />
                    <RANKING order="4" place="4" resultid="1331" />
                    <RANKING order="5" place="5" resultid="1316" />
                    <RANKING order="6" place="6" resultid="1311" />
                    <RANKING order="7" place="7" resultid="1291" />
                    <RANKING order="8" place="8" resultid="2005" />
                    <RANKING order="9" place="9" resultid="1193" />
                    <RANKING order="10" place="10" resultid="2092" />
                    <RANKING order="11" place="11" resultid="1241" />
                    <RANKING order="12" place="12" resultid="1922" />
                    <RANKING order="13" place="13" resultid="1190" />
                    <RANKING order="14" place="14" resultid="1933" />
                    <RANKING order="15" place="15" resultid="1405" />
                    <RANKING order="16" place="16" resultid="1453" />
                    <RANKING order="17" place="17" resultid="1228" />
                    <RANKING order="18" place="-1" resultid="2139" />
                    <RANKING order="19" place="-1" resultid="1296" />
                    <RANKING order="20" place="-1" resultid="1472" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2416" daytime="18:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2417" daytime="18:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2418" daytime="18:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2419" daytime="18:46" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2420" daytime="18:50" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1136" daytime="18:54" gender="F" number="29" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1137" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1955" />
                    <RANKING order="2" place="2" resultid="1661" />
                    <RANKING order="3" place="3" resultid="1173" />
                    <RANKING order="4" place="4" resultid="1221" />
                    <RANKING order="5" place="5" resultid="1771" />
                    <RANKING order="6" place="6" resultid="1837" />
                    <RANKING order="7" place="7" resultid="1746" />
                    <RANKING order="8" place="-1" resultid="1651" />
                    <RANKING order="9" place="-1" resultid="1706" />
                    <RANKING order="10" place="-1" resultid="1791" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1995" />
                    <RANKING order="2" place="2" resultid="1517" />
                    <RANKING order="3" place="3" resultid="1711" />
                    <RANKING order="4" place="4" resultid="1577" />
                    <RANKING order="5" place="5" resultid="1158" />
                    <RANKING order="6" place="6" resultid="2130" />
                    <RANKING order="7" place="7" resultid="1163" />
                    <RANKING order="8" place="8" resultid="2135" />
                    <RANKING order="9" place="9" resultid="1960" />
                    <RANKING order="10" place="10" resultid="1180" />
                    <RANKING order="11" place="11" resultid="2083" />
                    <RANKING order="12" place="12" resultid="1971" />
                    <RANKING order="13" place="13" resultid="1913" />
                    <RANKING order="14" place="14" resultid="1552" />
                    <RANKING order="15" place="15" resultid="2125" />
                    <RANKING order="16" place="16" resultid="1268" />
                    <RANKING order="17" place="-1" resultid="1582" />
                    <RANKING order="18" place="-1" resultid="1597" />
                    <RANKING order="19" place="-1" resultid="1627" />
                    <RANKING order="20" place="-1" resultid="1786" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2421" daytime="18:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2422" daytime="18:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2423" daytime="18:58" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2424" daytime="19:00" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1139" daytime="19:02" gender="M" number="30" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1140" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1647" />
                    <RANKING order="2" place="2" resultid="2065" />
                    <RANKING order="3" place="3" resultid="1238" />
                    <RANKING order="4" place="4" resultid="1682" />
                    <RANKING order="5" place="5" resultid="1874" />
                    <RANKING order="6" place="6" resultid="2145" />
                    <RANKING order="7" place="7" resultid="1910" />
                    <RANKING order="8" place="8" resultid="2153" />
                    <RANKING order="9" place="9" resultid="1767" />
                    <RANKING order="10" place="10" resultid="2159" />
                    <RANKING order="11" place="11" resultid="1777" />
                    <RANKING order="12" place="12" resultid="1782" />
                    <RANKING order="13" place="13" resultid="2156" />
                    <RANKING order="14" place="14" resultid="2162" />
                    <RANKING order="15" place="-1" resultid="1633" />
                    <RANKING order="16" place="-1" resultid="1727" />
                    <RANKING order="17" place="-1" resultid="1742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1141" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1593" />
                    <RANKING order="2" place="2" resultid="1919" />
                    <RANKING order="3" place="3" resultid="1508" />
                    <RANKING order="4" place="4" resultid="1672" />
                    <RANKING order="5" place="5" resultid="2026" />
                    <RANKING order="6" place="6" resultid="1528" />
                    <RANKING order="7" place="7" resultid="1177" />
                    <RANKING order="8" place="8" resultid="1167" />
                    <RANKING order="9" place="9" resultid="1588" />
                    <RANKING order="10" place="10" resultid="1213" />
                    <RANKING order="11" place="11" resultid="2098" />
                    <RANKING order="12" place="12" resultid="2089" />
                    <RANKING order="13" place="13" resultid="2103" />
                    <RANKING order="14" place="14" resultid="2021" />
                    <RANKING order="15" place="15" resultid="1234" />
                    <RANKING order="16" place="16" resultid="1657" />
                    <RANKING order="17" place="17" resultid="1802" />
                    <RANKING order="18" place="18" resultid="1563" />
                    <RANKING order="19" place="19" resultid="1548" />
                    <RANKING order="20" place="20" resultid="1543" />
                    <RANKING order="21" place="21" resultid="1185" />
                    <RANKING order="22" place="22" resultid="1573" />
                    <RANKING order="23" place="23" resultid="2113" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2425" daytime="19:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2426" daytime="19:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2427" daytime="19:08" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2428" daytime="19:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2429" daytime="19:12" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1142" daytime="19:14" gender="F" number="31" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1143" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1392" />
                    <RANKING order="2" place="2" resultid="1382" />
                    <RANKING order="3" place="3" resultid="1762" />
                    <RANKING order="4" place="4" resultid="1170" />
                    <RANKING order="5" place="5" resultid="1900" />
                    <RANKING order="6" place="6" resultid="2150" />
                    <RANKING order="7" place="7" resultid="2030" />
                    <RANKING order="8" place="8" resultid="1608" />
                    <RANKING order="9" place="9" resultid="2074" />
                    <RANKING order="10" place="10" resultid="1943" />
                    <RANKING order="11" place="11" resultid="1225" />
                    <RANKING order="12" place="-1" resultid="2016" />
                    <RANKING order="13" place="-1" resultid="1411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1144" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1337" />
                    <RANKING order="2" place="2" resultid="2108" />
                    <RANKING order="3" place="3" resultid="1362" />
                    <RANKING order="4" place="4" resultid="1752" />
                    <RANKING order="5" place="5" resultid="1991" />
                    <RANKING order="6" place="6" resultid="1603" />
                    <RANKING order="7" place="7" resultid="1218" />
                    <RANKING order="8" place="8" resultid="1503" />
                    <RANKING order="9" place="9" resultid="1342" />
                    <RANKING order="10" place="10" resultid="1199" />
                    <RANKING order="11" place="11" resultid="1444" />
                    <RANKING order="12" place="12" resultid="1977" />
                    <RANKING order="13" place="13" resultid="2121" />
                    <RANKING order="14" place="-1" resultid="1347" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2430" daytime="19:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2431" daytime="19:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2432" daytime="19:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2433" daytime="19:20" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1145" daytime="19:24" gender="M" number="32" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1146" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1834" />
                    <RANKING order="2" place="2" resultid="2045" />
                    <RANKING order="3" place="3" resultid="1449" />
                    <RANKING order="4" place="4" resultid="1253" />
                    <RANKING order="5" place="5" resultid="1439" />
                    <RANKING order="6" place="6" resultid="2055" />
                    <RANKING order="7" place="7" resultid="1478" />
                    <RANKING order="8" place="8" resultid="1464" />
                    <RANKING order="9" place="9" resultid="1278" />
                    <RANKING order="10" place="10" resultid="1429" />
                    <RANKING order="11" place="11" resultid="2117" />
                    <RANKING order="12" place="12" resultid="1905" />
                    <RANKING order="13" place="13" resultid="1930" />
                    <RANKING order="14" place="-1" resultid="1402" />
                    <RANKING order="15" place="-1" resultid="1891" />
                    <RANKING order="16" place="-1" resultid="1841" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1327" />
                    <RANKING order="2" place="2" resultid="1986" />
                    <RANKING order="3" place="3" resultid="1352" />
                    <RANKING order="4" place="4" resultid="1208" />
                    <RANKING order="5" place="5" resultid="1194" />
                    <RANKING order="6" place="6" resultid="1357" />
                    <RANKING order="7" place="7" resultid="1939" />
                    <RANKING order="8" place="8" resultid="2070" />
                    <RANKING order="9" place="9" resultid="1923" />
                    <RANKING order="10" place="10" resultid="1281" />
                    <RANKING order="11" place="11" resultid="1229" />
                    <RANKING order="12" place="12" resultid="1454" />
                    <RANKING order="13" place="13" resultid="2093" />
                    <RANKING order="14" place="-1" resultid="2006" />
                    <RANKING order="15" place="-1" resultid="1406" />
                    <RANKING order="16" place="-1" resultid="1322" />
                    <RANKING order="17" place="-1" resultid="1367" />
                    <RANKING order="18" place="-1" resultid="1473" />
                    <RANKING order="19" place="-1" resultid="1498" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2434" daytime="19:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2435" daytime="19:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2436" daytime="19:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2437" daytime="19:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2438" daytime="19:32" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="1883" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Frederico" lastname="Massad Andrade" birthdate="2012-03-22" gender="M" nation="BRA" license="416948" athleteid="1931" externalid="416948">
              <RESULTS>
                <RESULT eventid="1089" points="182" swimtime="00:01:22.61" resultid="1932" heatid="2360" lane="2" />
                <RESULT eventid="1133" points="133" swimtime="00:01:41.07" resultid="1933" heatid="2418" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Samuel" lastname="Melo Lima" birthdate="2015-10-30" gender="M" nation="BRA" license="406933" swrid="5725994" athleteid="1906" externalid="406933">
              <RESULTS>
                <RESULT eventid="1095" points="27" swimtime="00:01:13.72" resultid="1907" heatid="2368" lane="7" />
                <RESULT eventid="1083" points="69" swimtime="00:01:03.09" resultid="1908" heatid="2350" lane="7" entrytime="00:01:02.06" entrycourse="LCM" />
                <RESULT eventid="1127" points="82" swimtime="00:00:54.01" resultid="1909" heatid="2409" lane="8" entrytime="00:00:55.81" entrycourse="LCM" />
                <RESULT eventid="1139" points="85" swimtime="00:00:47.52" resultid="1910" heatid="2426" lane="2" entrytime="00:00:50.19" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Borges Duarte" birthdate="2014-02-10" gender="F" nation="BRA" license="408688" swrid="5725985" athleteid="1911" externalid="408688">
              <RESULTS>
                <RESULT eventid="1064" points="170" swimtime="00:03:23.44" resultid="1912" heatid="2328" lane="1" />
                <RESULT eventid="1136" points="175" swimtime="00:00:42.18" resultid="1913" heatid="2422" lane="3" entrytime="00:00:43.25" entrycourse="LCM" />
                <RESULT eventid="1124" points="153" swimtime="00:00:50.17" resultid="1914" heatid="2404" lane="6" entrytime="00:00:50.47" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Paes Schemiko" birthdate="2013-02-25" gender="F" nation="BRA" license="406918" swrid="5725995" athleteid="1896" externalid="406918">
              <RESULTS>
                <RESULT eventid="1098" points="237" swimtime="00:00:39.47" resultid="1897" heatid="2373" lane="4" entrytime="00:00:42.23" entrycourse="LCM" />
                <RESULT eventid="1086" points="292" swimtime="00:01:17.88" resultid="1898" heatid="2353" lane="5" />
                <RESULT eventid="1130" points="243" swimtime="00:01:31.85" resultid="1899" heatid="2411" lane="3" />
                <RESULT eventid="1142" points="260" swimtime="00:00:45.68" resultid="1900" heatid="2431" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Henrique Ballatka" birthdate="2013-08-26" gender="M" nation="BRA" license="405839" swrid="5697229" athleteid="1889" externalid="405839">
              <RESULTS>
                <RESULT eventid="1089" points="91" swimtime="00:01:44.06" resultid="1890" heatid="2360" lane="7" />
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada.  (Horário: 19:18)" eventid="1145" status="DSQ" swimtime="00:00:55.65" resultid="1891" heatid="2435" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Manoel Forte" birthdate="2013-01-13" gender="M" nation="BRA" license="414859" swrid="5755340" athleteid="1927" externalid="414859">
              <RESULTS>
                <RESULT comment="SW 10.7 - Puxou a corda da raia &quot;lane rope&quot;.  (Horário: 11:36)" eventid="1089" status="DSQ" swimtime="00:02:00.20" resultid="1928" heatid="2359" lane="2" />
                <RESULT eventid="1133" points="83" swimtime="00:01:58.15" resultid="1929" heatid="2419" lane="8" />
                <RESULT eventid="1145" points="64" swimtime="00:01:04.69" resultid="1930" heatid="2434" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Ribeiro Melo" birthdate="2013-02-25" gender="M" nation="BRA" license="406921" swrid="5717293" athleteid="1901" externalid="406921">
              <RESULTS>
                <RESULT eventid="1089" points="198" swimtime="00:01:20.32" resultid="1902" heatid="2363" lane="1" entrytime="00:01:20.96" entrycourse="LCM" />
                <RESULT eventid="1073" points="163" swimtime="00:03:28.37" resultid="1903" heatid="2339" lane="3" entrytime="00:03:31.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="152" swimtime="00:01:36.68" resultid="1904" heatid="2418" lane="6" />
                <RESULT eventid="1145" points="91" swimtime="00:00:57.57" resultid="1905" heatid="2436" lane="3" entrytime="00:00:53.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Schneider Yazbek" birthdate="2013-03-07" gender="F" nation="BRA" license="378329" swrid="5588907" athleteid="1884" externalid="378329">
              <RESULTS>
                <RESULT eventid="1086" points="343" swimtime="00:01:13.80" resultid="1885" heatid="2357" lane="4" entrytime="00:01:16.37" entrycourse="LCM" />
                <RESULT eventid="1070" points="312" swimtime="00:03:05.77" resultid="1886" heatid="2338" lane="1" entrytime="00:03:04.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="250" swimtime="00:01:30.96" resultid="1887" heatid="2412" lane="2" />
                <RESULT eventid="1114" points="381" swimtime="00:05:24.58" resultid="1888" heatid="2392" lane="4" entrytime="00:05:44.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.33" />
                    <SPLIT distance="200" swimtime="00:02:42.04" />
                    <SPLIT distance="300" swimtime="00:04:06.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="De Ormeno" birthdate="2014-04-02" gender="M" nation="BRA" license="408702" swrid="5740009" athleteid="1915" externalid="408702">
              <RESULTS>
                <RESULT eventid="1095" points="151" swimtime="00:00:41.79" resultid="1916" heatid="2369" lane="5" entrytime="00:00:44.96" entrycourse="LCM" />
                <RESULT eventid="1067" points="220" swimtime="00:02:48.89" resultid="1917" heatid="2332" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="208" swimtime="00:00:39.71" resultid="1918" heatid="2410" lane="4" entrytime="00:00:40.16" entrycourse="LCM" />
                <RESULT eventid="1139" points="229" swimtime="00:00:34.17" resultid="1919" heatid="2429" lane="3" entrytime="00:00:34.47" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benicio" lastname="Alves" birthdate="2012-04-26" gender="M" nation="BRA" license="370588" swrid="5740005" athleteid="1920" externalid="370588">
              <RESULTS>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 11:42)" eventid="1089" status="DSQ" swimtime="00:00:00.00" resultid="1921" heatid="2361" lane="6" entrytime="00:01:27.75" entrycourse="LCM" />
                <RESULT eventid="1133" points="165" swimtime="00:01:34.00" resultid="1922" heatid="2416" lane="5" />
                <RESULT eventid="1145" points="117" swimtime="00:00:52.98" resultid="1923" heatid="2435" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Siqueira Lopes" birthdate="2012-04-28" gender="F" nation="BRA" license="414671" swrid="5755342" athleteid="1924" externalid="414671">
              <RESULTS>
                <RESULT eventid="1086" points="298" swimtime="00:01:17.40" resultid="1925" heatid="2354" lane="7" />
                <RESULT eventid="1070" points="256" swimtime="00:03:18.57" resultid="1926" heatid="2335" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Zanatta Duda" birthdate="2013-08-28" gender="F" nation="BRA" license="406914" swrid="5717306" athleteid="1892" externalid="406914">
              <RESULTS>
                <RESULT eventid="1098" points="62" swimtime="00:01:01.72" resultid="1893" heatid="2372" lane="8" />
                <RESULT eventid="1086" points="177" swimtime="00:01:32.07" resultid="1894" heatid="2355" lane="4" entrytime="00:01:39.14" entrycourse="LCM" />
                <RESULT eventid="1130" points="155" swimtime="00:01:46.53" resultid="1895" heatid="2414" lane="8" entrytime="00:01:48.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="263" nation="BRA" region="PR" clubid="1282" swrid="75436" name="Clube Curitibano" shortname="Curitibano">
          <ATHLETES>
            <ATHLETE firstname="Lucas" lastname="Azevedo Alanis" birthdate="2013-12-07" gender="M" nation="BRA" license="376991" swrid="5588540" athleteid="1474" externalid="376991">
              <RESULTS>
                <RESULT eventid="1089" points="159" swimtime="00:01:26.46" resultid="1475" heatid="2361" lane="1" entrytime="00:01:30.72" entrycourse="LCM" />
                <RESULT eventid="1073" points="172" swimtime="00:03:24.89" resultid="1476" heatid="2340" lane="8" entrytime="00:03:22.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="185" swimtime="00:06:26.22" resultid="1477" heatid="2395" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.81" />
                    <SPLIT distance="200" swimtime="00:03:11.50" />
                    <SPLIT distance="300" swimtime="00:04:50.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="151" swimtime="00:00:48.63" resultid="1478" heatid="2437" lane="2" entrytime="00:00:50.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Francia Soares" birthdate="2014-06-01" gender="F" nation="BRA" license="391011" swrid="5602540" athleteid="1549" externalid="391011">
              <RESULTS>
                <RESULT eventid="1080" points="83" swimtime="00:01:06.68" resultid="1550" heatid="2346" lane="8" entrytime="00:01:21.02" entrycourse="LCM" />
                <RESULT eventid="1064" points="144" swimtime="00:03:35.06" resultid="1551" heatid="2329" lane="4" entrytime="00:03:37.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="173" swimtime="00:00:42.32" resultid="1552" heatid="2422" lane="4" entrytime="00:00:42.89" entrycourse="LCM" />
                <RESULT eventid="1124" points="95" swimtime="00:00:58.85" resultid="1553" heatid="2402" lane="4" entrytime="00:01:01.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Hallage Papp" birthdate="2012-07-02" gender="M" nation="BRA" license="377042" swrid="5588736" athleteid="1470" externalid="377042">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="1471" heatid="2362" lane="2" entrytime="00:01:23.78" entrycourse="LCM" />
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="1472" heatid="2418" lane="7" />
                <RESULT eventid="1145" status="DNS" swimtime="00:00:00.00" resultid="1473" heatid="2436" lane="2" entrytime="00:00:54.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Brandt Macedo" birthdate="2013-04-19" gender="M" nation="BRA" license="414421" swrid="5755329" athleteid="1839" externalid="414421">
              <RESULTS>
                <RESULT eventid="1089" points="63" swimtime="00:01:57.26" resultid="1840" heatid="2360" lane="8" />
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 19:15)" eventid="1145" status="DSQ" swimtime="00:01:05.24" resultid="1841" heatid="2434" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Schmidt Wozniaki" birthdate="2012-07-07" gender="M" nation="BRA" license="376963" swrid="5588905" athleteid="1403" externalid="376963">
              <RESULTS>
                <RESULT eventid="1089" points="170" swimtime="00:01:24.44" resultid="1404" heatid="2359" lane="4" />
                <RESULT eventid="1133" points="104" swimtime="00:01:49.61" resultid="1405" heatid="2417" lane="7" />
                <RESULT comment="SW 7.1 - A cabeça não rompeu a superfície antes que as mãos se virassem para dentro na parte mais ampla do segundo movimento após o início ou a virada.&#10;&#10;&#10;&#10;&#10;&#10;&#10;  (Horário: 19:23), Após a saída." eventid="1145" status="DSQ" swimtime="00:00:51.22" resultid="1406" heatid="2437" lane="8" entrytime="00:00:52.03" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Della Villa Yang" birthdate="2015-02-27" gender="F" nation="BRA" license="393283" swrid="5616442" athleteid="1658" externalid="393283">
              <RESULTS>
                <RESULT eventid="1092" points="112" swimtime="00:00:50.61" resultid="1659" heatid="2366" lane="6" entrytime="00:00:51.17" entrycourse="LCM" />
                <RESULT eventid="1064" points="180" swimtime="00:03:19.79" resultid="1660" heatid="2330" lane="7" entrytime="00:03:33.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="210" swimtime="00:00:39.68" resultid="1661" heatid="2423" lane="7" entrytime="00:00:41.98" entrycourse="LCM" />
                <RESULT eventid="1108" points="183" swimtime="00:03:41.87" resultid="1662" heatid="2385" lane="2" entrytime="00:03:52.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:51.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gael" lastname="Stramandinoli Zanicotti" birthdate="2015-03-21" gender="M" nation="BRA" license="406954" swrid="5717298" athleteid="1763" externalid="406954">
              <RESULTS>
                <RESULT eventid="1095" points="18" swimtime="00:01:24.47" resultid="1764" heatid="2368" lane="5" entrytime="00:01:25.97" entrycourse="LCM" />
                <RESULT eventid="1067" points="51" swimtime="00:04:33.82" resultid="1765" heatid="2332" lane="8" />
                <RESULT eventid="1127" points="44" swimtime="00:01:06.61" resultid="1766" heatid="2408" lane="1" entrytime="00:01:01.23" entrycourse="LCM" />
                <RESULT eventid="1139" points="52" swimtime="00:00:55.71" resultid="1767" heatid="2426" lane="1" entrytime="00:00:56.59" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="De Lima Cavalcanti" birthdate="2014-10-07" gender="M" nation="BRA" license="385884" swrid="5684550" athleteid="1713" externalid="385884">
              <RESULTS>
                <RESULT eventid="1083" points="117" swimtime="00:00:52.96" resultid="1714" heatid="2349" lane="1" />
                <RESULT eventid="1067" points="195" swimtime="00:02:55.83" resultid="1715" heatid="2334" lane="2" entrytime="00:03:02.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="191" swimtime="00:00:40.88" resultid="1716" heatid="2410" lane="5" entrytime="00:00:40.63" entrycourse="LCM" />
                <RESULT eventid="1111" points="151" swimtime="00:03:33.62" resultid="1717" heatid="2387" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Tallao Benke" birthdate="2012-01-02" gender="F" nation="BRA" license="376984" swrid="5588931" athleteid="1455" externalid="376984">
              <RESULTS>
                <RESULT eventid="1098" points="410" swimtime="00:00:32.88" resultid="1456" heatid="2374" lane="5" entrytime="00:00:33.98" entrycourse="LCM" />
                <RESULT eventid="1086" points="495" swimtime="00:01:05.36" resultid="1457" heatid="2354" lane="2" />
                <RESULT eventid="1130" points="438" swimtime="00:01:15.45" resultid="1458" heatid="2415" lane="4" entrytime="00:01:16.06" entrycourse="LCM" />
                <RESULT eventid="1114" points="464" swimtime="00:05:03.87" resultid="1459" heatid="2393" lane="4" entrytime="00:05:06.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.09" />
                    <SPLIT distance="200" swimtime="00:02:29.07" />
                    <SPLIT distance="300" swimtime="00:03:49.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joana" lastname="Asinelli Casagrande" birthdate="2013-10-26" gender="F" nation="BRA" license="376970" swrid="5588536" athleteid="1417" externalid="376970">
              <RESULTS>
                <RESULT eventid="1130" points="298" swimtime="00:01:25.75" resultid="1418" heatid="2414" lane="4" entrytime="00:01:28.72" entrycourse="LCM" />
                <RESULT eventid="1114" points="271" swimtime="00:06:03.64" resultid="1419" heatid="2391" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.85" />
                    <SPLIT distance="200" swimtime="00:03:02.40" />
                    <SPLIT distance="300" swimtime="00:04:36.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Henrique Tiboni Araujo" birthdate="2013-06-11" gender="M" nation="BRA" license="376968" swrid="5588747" athleteid="1412" externalid="376968">
              <RESULTS>
                <RESULT eventid="1101" points="172" swimtime="00:00:40.01" resultid="1413" heatid="2376" lane="5" entrytime="00:00:49.38" entrycourse="LCM" />
                <RESULT eventid="1089" points="197" swimtime="00:01:20.52" resultid="1414" heatid="2361" lane="7" entrytime="00:01:28.29" entrycourse="LCM" />
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="1415" heatid="2419" lane="2" entrytime="00:01:41.79" entrycourse="LCM" />
                <RESULT eventid="1117" status="DNS" swimtime="00:00:00.00" resultid="1416" heatid="2394" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Pacheco" birthdate="2012-10-13" gender="F" nation="BRA" license="376981" swrid="5602566" athleteid="1440" externalid="376981">
              <RESULTS>
                <RESULT eventid="1098" points="56" swimtime="00:01:03.76" resultid="1441" heatid="2372" lane="2" />
                <RESULT eventid="1086" points="219" swimtime="00:01:25.77" resultid="1442" heatid="2356" lane="1" entrytime="00:01:32.88" entrycourse="LCM" />
                <RESULT eventid="1114" points="197" swimtime="00:06:44.29" resultid="1443" heatid="2392" lane="1" entrytime="00:07:04.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.92" />
                    <SPLIT distance="200" swimtime="00:03:18.76" />
                    <SPLIT distance="300" swimtime="00:05:02.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="176" swimtime="00:00:52.01" resultid="1444" heatid="2432" lane="7" entrytime="00:00:54.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Da Cunha Souza" birthdate="2015-05-30" gender="F" nation="BRA" license="400016" swrid="5652883" athleteid="1698" externalid="400016">
              <RESULTS>
                <RESULT eventid="1092" points="125" swimtime="00:00:48.83" resultid="1699" heatid="2366" lane="2" entrytime="00:00:52.13" entrycourse="LCM" />
                <RESULT eventid="1064" points="182" swimtime="00:03:18.98" resultid="1700" heatid="2329" lane="3" entrytime="00:03:44.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="172" swimtime="00:00:48.21" resultid="1701" heatid="2405" lane="3" entrytime="00:00:45.72" entrycourse="LCM" />
                <RESULT eventid="1108" points="157" swimtime="00:03:53.74" resultid="1702" heatid="2384" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Viera Correa" birthdate="2012-03-07" gender="M" nation="BRA" license="369269" swrid="5602590" athleteid="1313" externalid="369269">
              <RESULTS>
                <RESULT eventid="1101" points="226" swimtime="00:00:36.52" resultid="1314" heatid="2376" lane="1" />
                <RESULT eventid="1089" points="340" swimtime="00:01:07.09" resultid="1315" heatid="2364" lane="3" entrytime="00:01:09.41" entrycourse="LCM" />
                <RESULT eventid="1133" points="226" swimtime="00:01:24.66" resultid="1316" heatid="2420" lane="6" entrytime="00:01:23.38" entrycourse="LCM" />
                <RESULT eventid="1117" points="314" swimtime="00:05:23.71" resultid="1317" heatid="2397" lane="3" entrytime="00:05:31.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.64" />
                    <SPLIT distance="200" swimtime="00:02:37.48" />
                    <SPLIT distance="300" swimtime="00:04:02.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Guimaraes Mesquita" birthdate="2015-10-05" gender="F" nation="BRA" license="393263" swrid="5616444" athleteid="1648" externalid="393263">
              <RESULTS>
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="1649" heatid="2346" lane="7" entrytime="00:01:10.17" entrycourse="LCM" />
                <RESULT eventid="1064" status="DNS" swimtime="00:00:00.00" resultid="1650" heatid="2328" lane="7" />
                <RESULT eventid="1136" status="DNS" swimtime="00:00:00.00" resultid="1651" heatid="2421" lane="6" entrytime="00:00:56.88" entrycourse="LCM" />
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="1652" heatid="2402" lane="3" entrytime="00:01:03.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Almeida Jorge" birthdate="2015-05-27" gender="M" nation="BRA" license="406836" swrid="5717242" athleteid="1753" externalid="406836">
              <RESULTS>
                <RESULT eventid="1083" points="76" swimtime="00:01:01.16" resultid="1754" heatid="2350" lane="1" entrytime="00:01:02.73" entrycourse="LCM" />
                <RESULT eventid="1067" points="63" swimtime="00:04:15.48" resultid="1755" heatid="2331" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:06.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="65" swimtime="00:00:58.52" resultid="1756" heatid="2408" lane="3" entrytime="00:00:56.88" entrycourse="LCM" />
                <RESULT eventid="1111" points="73" swimtime="00:04:31.84" resultid="1757" heatid="2386" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:14.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Cipriani Presiazniuk" birthdate="2012-07-03" gender="M" nation="BRA" license="369267" swrid="5588594" athleteid="1308" externalid="369267">
              <RESULTS>
                <RESULT eventid="1089" points="278" swimtime="00:01:11.77" resultid="1309" heatid="2363" lane="3" entrytime="00:01:16.43" entrycourse="LCM" />
                <RESULT eventid="1073" points="221" swimtime="00:03:08.36" resultid="1310" heatid="2340" lane="7" entrytime="00:03:13.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="211" swimtime="00:01:26.61" resultid="1311" heatid="2419" lane="4" entrytime="00:01:30.49" entrycourse="LCM" />
                <RESULT eventid="1117" points="253" swimtime="00:05:47.89" resultid="1312" heatid="2395" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.67" />
                    <SPLIT distance="200" swimtime="00:02:54.19" />
                    <SPLIT distance="300" swimtime="00:04:24.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Caron Braga" birthdate="2016-02-01" gender="F" nation="BRA" license="415256" swrid="5755333" athleteid="1864" externalid="415256">
              <RESULTS>
                <RESULT eventid="1076" points="65" swimtime="00:01:06.76" resultid="1865" heatid="2342" lane="5" />
                <RESULT eventid="1120" points="71" swimtime="00:00:56.92" resultid="1866" heatid="2398" lane="4" entrytime="00:01:08.36" entrycourse="LCM" />
                <RESULT eventid="1104" points="54" swimtime="00:01:16.95" resultid="1867" heatid="2380" lane="7" entrytime="00:01:11.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Marie Silva" birthdate="2014-08-24" gender="F" nation="BRA" license="391025" swrid="5602556" athleteid="1594" externalid="391025">
              <RESULTS>
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="1595" heatid="2347" lane="1" entrytime="00:01:00.06" entrycourse="LCM" />
                <RESULT eventid="1064" status="DNS" swimtime="00:00:00.00" resultid="1596" heatid="2330" lane="2" entrytime="00:03:22.07" entrycourse="LCM" />
                <RESULT eventid="1136" status="DNS" swimtime="00:00:00.00" resultid="1597" heatid="2421" lane="7" />
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="1598" heatid="2402" lane="6" entrytime="00:01:04.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Miranda Carvalho" birthdate="2015-07-07" gender="F" nation="BRA" license="410200" swrid="5740015" athleteid="1788" externalid="410200">
              <RESULTS>
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="1789" heatid="2346" lane="2" entrytime="00:01:09.01" entrycourse="LCM" />
                <RESULT eventid="1064" status="DNS" swimtime="00:00:00.00" resultid="1790" heatid="2327" lane="3" />
                <RESULT eventid="1136" status="DNS" swimtime="00:00:00.00" resultid="1791" heatid="2421" lane="3" entrytime="00:00:56.54" entrycourse="LCM" />
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="1792" heatid="2402" lane="5" entrytime="00:01:02.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Caron Braga" birthdate="2016-02-01" gender="F" nation="BRA" license="415257" swrid="5755332" athleteid="1868" externalid="415257">
              <RESULTS>
                <RESULT eventid="1076" points="77" swimtime="00:01:02.88" resultid="1869" heatid="2342" lane="3" />
                <RESULT eventid="1120" points="49" swimtime="00:01:04.19" resultid="1870" heatid="2398" lane="5" entrytime="00:01:09.32" entrycourse="LCM" />
                <RESULT eventid="1104" points="66" swimtime="00:01:12.01" resultid="1871" heatid="2380" lane="1" entrytime="00:01:18.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Felipe Canalli" birthdate="2015-12-23" gender="M" nation="BRA" license="406749" swrid="5717261" athleteid="1738" externalid="406749">
              <RESULTS>
                <RESULT eventid="1083" points="144" swimtime="00:00:49.41" resultid="1739" heatid="2352" lane="1" entrytime="00:00:51.04" entrycourse="LCM" />
                <RESULT eventid="1067" points="66" swimtime="00:04:11.92" resultid="1740" heatid="2331" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:58.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" status="DNS" swimtime="00:00:00.00" resultid="1741" heatid="2387" lane="4" entrytime="00:04:49.80" entrycourse="LCM" />
                <RESULT eventid="1139" status="DNS" swimtime="00:00:00.00" resultid="1742" heatid="2425" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Fernandes  Dos Reis" birthdate="2012-09-18" gender="M" nation="BRA" license="369279" swrid="5588696" athleteid="1353" externalid="369279">
              <RESULTS>
                <RESULT eventid="1101" points="250" swimtime="00:00:35.31" resultid="1354" heatid="2378" lane="5" entrytime="00:00:34.87" entrycourse="LCM" />
                <RESULT eventid="1073" points="235" swimtime="00:03:04.61" resultid="1355" heatid="2341" lane="6" entrytime="00:03:03.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="267" swimtime="00:05:41.39" resultid="1356" heatid="2397" lane="2" entrytime="00:05:39.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.22" />
                    <SPLIT distance="200" swimtime="00:02:44.56" />
                    <SPLIT distance="300" swimtime="00:04:13.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="157" swimtime="00:00:48.04" resultid="1357" heatid="2436" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="De Fortes" birthdate="2015-06-01" gender="M" nation="BRA" license="399680" swrid="5652884" athleteid="1688" externalid="399680">
              <RESULTS>
                <RESULT eventid="1095" points="98" swimtime="00:00:48.24" resultid="1689" heatid="2369" lane="3" entrytime="00:00:47.21" entrycourse="LCM" />
                <RESULT eventid="1067" status="DNS" swimtime="00:00:00.00" resultid="1690" heatid="2333" lane="3" entrytime="00:03:49.34" entrycourse="LCM" />
                <RESULT eventid="1127" points="113" swimtime="00:00:48.69" resultid="1691" heatid="2409" lane="2" entrytime="00:00:50.38" entrycourse="LCM" />
                <RESULT eventid="1111" status="DNS" swimtime="00:00:00.00" resultid="1692" heatid="2388" lane="2" entrytime="00:04:19.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Cavalcanti Breginski" birthdate="2016-04-06" gender="F" nation="BRA" license="415012" swrid="5755334" athleteid="1849" externalid="415012">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="1850" heatid="2343" lane="6" entrytime="00:01:05.62" entrycourse="LCM" />
                <RESULT eventid="1120" status="DNS" swimtime="00:00:00.00" resultid="1851" heatid="2399" lane="7" entrytime="00:01:07.28" entrycourse="LCM" />
                <RESULT eventid="1104" status="DNS" swimtime="00:00:00.00" resultid="1852" heatid="2379" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Antunes Saboia" birthdate="2012-06-28" gender="M" nation="BRA" license="369278" swrid="5602511" athleteid="1348" externalid="369278">
              <RESULTS>
                <RESULT eventid="1089" points="301" swimtime="00:01:09.88" resultid="1349" heatid="2364" lane="2" entrytime="00:01:10.67" entrycourse="LCM" />
                <RESULT eventid="1073" points="261" swimtime="00:02:58.18" resultid="1350" heatid="2341" lane="3" entrytime="00:02:57.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="300" swimtime="00:05:28.39" resultid="1351" heatid="2394" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.89" />
                    <SPLIT distance="200" swimtime="00:02:43.04" />
                    <SPLIT distance="300" swimtime="00:04:07.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="246" swimtime="00:00:41.39" resultid="1352" heatid="2438" lane="3" entrytime="00:00:41.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Rossi Mattioli" birthdate="2013-05-08" gender="F" nation="BRA" license="376988" swrid="5588892" athleteid="1489" externalid="376988">
              <RESULTS>
                <RESULT eventid="1098" points="244" swimtime="00:00:39.09" resultid="1490" heatid="2373" lane="2" entrytime="00:00:47.70" entrycourse="LCM" />
                <RESULT eventid="1086" points="297" swimtime="00:01:17.44" resultid="1491" heatid="2357" lane="7" entrytime="00:01:20.58" entrycourse="LCM" />
                <RESULT comment="SW 6.5 - Não terminou a prova enquanto estava de costas.&#10;&#10;&#10;&#10;&#10;&#10;&#10;  (Horário: 18:13)" eventid="1130" status="DSQ" swimtime="00:01:36.84" resultid="1492" heatid="2411" lane="4" />
                <RESULT eventid="1114" points="245" swimtime="00:06:15.90" resultid="1493" heatid="2392" lane="2" entrytime="00:06:16.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.04" />
                    <SPLIT distance="200" swimtime="00:03:06.62" />
                    <SPLIT distance="300" swimtime="00:04:44.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Afonso Fowler" birthdate="2014-01-22" gender="M" nation="BRA" license="393264" swrid="5661338" athleteid="1653" externalid="393264">
              <RESULTS>
                <RESULT eventid="1083" points="83" swimtime="00:00:59.32" resultid="1654" heatid="2349" lane="5" entrytime="00:01:10.86" entrycourse="LCM" />
                <RESULT eventid="1067" points="106" swimtime="00:03:35.44" resultid="1655" heatid="2331" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="100" swimtime="00:00:50.66" resultid="1656" heatid="2409" lane="3" entrytime="00:00:49.09" entrycourse="LCM" />
                <RESULT eventid="1139" points="131" swimtime="00:00:41.09" resultid="1657" heatid="2428" lane="3" entrytime="00:00:37.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Della Villa Yang" birthdate="2012-10-08" gender="F" nation="BRA" license="369276" swrid="5588653" athleteid="1338" externalid="369276">
              <RESULTS>
                <RESULT eventid="1098" points="269" swimtime="00:00:37.84" resultid="1339" heatid="2374" lane="3" entrytime="00:00:36.96" entrycourse="LCM" />
                <RESULT eventid="1070" points="346" swimtime="00:02:59.54" resultid="1340" heatid="2338" lane="3" entrytime="00:02:57.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="418" swimtime="00:05:14.61" resultid="1341" heatid="2393" lane="3" entrytime="00:05:11.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.54" />
                    <SPLIT distance="200" swimtime="00:02:35.16" />
                    <SPLIT distance="300" swimtime="00:03:56.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="214" swimtime="00:00:48.70" resultid="1342" heatid="2431" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Nishimura Ramina" birthdate="2013-11-25" gender="M" nation="BRA" license="376989" swrid="5588831" athleteid="1484" externalid="376989">
              <RESULTS>
                <RESULT eventid="1101" points="110" swimtime="00:00:46.40" resultid="1485" heatid="2376" lane="3" entrytime="00:00:58.19" entrycourse="LCM" />
                <RESULT eventid="1089" points="166" swimtime="00:01:25.10" resultid="1486" heatid="2360" lane="5" entrytime="00:01:39.12" entrycourse="LCM" />
                <RESULT eventid="1133" points="145" swimtime="00:01:38.05" resultid="1487" heatid="2417" lane="2" />
                <RESULT eventid="1117" points="192" swimtime="00:06:20.90" resultid="1488" heatid="2396" lane="3" entrytime="00:06:27.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.65" />
                    <SPLIT distance="200" swimtime="00:03:05.52" />
                    <SPLIT distance="300" swimtime="00:04:45.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Livia Bittencourt" birthdate="2015-11-23" gender="F" nation="BRA" license="393260" swrid="5616446" athleteid="1634" externalid="393260">
              <RESULTS>
                <RESULT eventid="1080" points="92" swimtime="00:01:04.57" resultid="1635" heatid="2346" lane="6" entrytime="00:01:08.05" entrycourse="LCM" />
                <RESULT eventid="1064" points="86" swimtime="00:04:15.03" resultid="1636" heatid="2328" lane="6" />
                <RESULT eventid="1108" points="104" swimtime="00:04:27.78" resultid="1637" heatid="2382" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:12.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Magalhaes Dabul" birthdate="2014-01-05" gender="M" nation="BRA" license="391023" swrid="5602555" athleteid="1584" externalid="391023">
              <RESULTS>
                <RESULT eventid="1095" points="131" swimtime="00:00:43.77" resultid="1585" heatid="2370" lane="2" entrytime="00:00:42.17" entrycourse="LCM" />
                <RESULT eventid="1067" points="136" swimtime="00:03:17.88" resultid="1586" heatid="2333" lane="7" entrytime="00:04:02.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="153" swimtime="00:03:33.10" resultid="1587" heatid="2389" lane="7" entrytime="00:03:44.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="166" swimtime="00:00:38.03" resultid="1588" heatid="2428" lane="2" entrytime="00:00:38.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Hyczy Sarraff" birthdate="2016-12-22" gender="M" nation="BRA" license="415013" athleteid="1853" externalid="415013">
              <RESULTS>
                <RESULT eventid="1122" status="DNS" swimtime="00:00:00.00" resultid="1854" heatid="2400" lane="5" />
                <RESULT eventid="1106" status="DNS" swimtime="00:00:00.00" resultid="1855" heatid="2381" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Andrade Vosgerau" birthdate="2016-02-16" gender="F" nation="BRA" license="415010" swrid="5755328" athleteid="1842" externalid="415010">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="1843" heatid="2343" lane="7" entrytime="00:01:11.06" entrycourse="LCM" />
                <RESULT eventid="1120" status="DNS" swimtime="00:00:00.00" resultid="1844" heatid="2398" lane="3" />
                <RESULT eventid="1104" status="DNS" swimtime="00:00:00.00" resultid="1845" heatid="2379" lane="4" entrytime="00:01:15.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Jarenko Gomes" birthdate="2014-05-17" gender="F" nation="BRA" license="407692" swrid="5725992" athleteid="1783" externalid="407692">
              <RESULTS>
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="1784" heatid="2347" lane="8" entrytime="00:01:01.64" entrycourse="LCM" />
                <RESULT eventid="1064" points="105" swimtime="00:03:59.04" resultid="1785" heatid="2327" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" status="DNS" swimtime="00:00:00.00" resultid="1786" heatid="2421" lane="5" entrytime="00:00:51.11" entrycourse="LCM" />
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="1787" heatid="2403" lane="1" entrytime="00:00:57.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Paulo Celles" birthdate="2016-09-07" gender="M" nation="BRA" license="411996" swrid="5740017" athleteid="1803" externalid="411996">
              <RESULTS>
                <RESULT eventid="1122" status="DNS" swimtime="00:00:00.00" resultid="1804" heatid="2401" lane="2" entrytime="00:01:08.21" entrycourse="LCM" />
                <RESULT eventid="1106" status="DNS" swimtime="00:00:00.00" resultid="1805" heatid="2381" lane="3" entrytime="00:01:21.96" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Ribas Luz" birthdate="2015-02-05" gender="F" nation="BRA" license="406743" swrid="5717291" athleteid="1728" externalid="406743">
              <RESULTS>
                <RESULT eventid="1092" points="54" swimtime="00:01:04.30" resultid="1729" heatid="2365" lane="1" />
                <RESULT eventid="1064" points="85" swimtime="00:04:15.96" resultid="1730" heatid="2327" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:01.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="99" swimtime="00:00:57.98" resultid="1731" heatid="2404" lane="1" entrytime="00:00:53.10" entrycourse="LCM" />
                <RESULT eventid="1108" points="86" swimtime="00:04:45.49" resultid="1732" heatid="2384" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:15.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Sieczkowski Pacheco" birthdate="2015-11-20" gender="F" nation="BRA" license="393261" swrid="5616450" athleteid="1638" externalid="393261">
              <RESULTS>
                <RESULT eventid="1092" points="71" swimtime="00:00:58.84" resultid="1639" heatid="2365" lane="6" entrytime="00:00:56.60" entrycourse="LCM" />
                <RESULT eventid="1064" points="98" swimtime="00:04:03.97" resultid="1640" heatid="2329" lane="2" entrytime="00:03:54.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:54.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="101" swimtime="00:00:57.63" resultid="1641" heatid="2404" lane="8" entrytime="00:00:53.26" entrycourse="LCM" />
                <RESULT eventid="1108" points="123" swimtime="00:04:13.34" resultid="1642" heatid="2384" lane="4" entrytime="00:04:13.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:59.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="De Macedo Martynychen" birthdate="2015-06-12" gender="F" nation="BRA" license="399681" swrid="5652885" athleteid="1693" externalid="399681">
              <RESULTS>
                <RESULT eventid="1092" points="110" swimtime="00:00:50.87" resultid="1694" heatid="2365" lane="3" entrytime="00:00:56.52" entrycourse="LCM" />
                <RESULT eventid="1064" points="102" swimtime="00:04:01.05" resultid="1695" heatid="2328" lane="4" entrytime="00:04:13.92" entrycourse="LCM" />
                <RESULT eventid="1124" points="104" swimtime="00:00:57.01" resultid="1696" heatid="2403" lane="5" entrytime="00:00:56.76" entrycourse="LCM" />
                <RESULT eventid="1108" points="117" swimtime="00:04:17.73" resultid="1697" heatid="2383" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:04.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enrico" lastname="Calixto Rauen" birthdate="2016-06-25" gender="M" nation="BRA" license="415011" swrid="5755330" athleteid="1846" externalid="415011">
              <RESULTS>
                <RESULT eventid="1078" points="52" swimtime="00:01:03.06" resultid="1847" heatid="2344" lane="7" />
                <RESULT eventid="1122" status="DNS" swimtime="00:00:00.00" resultid="1848" heatid="2401" lane="3" entrytime="00:01:02.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Vanzo Assumpcao" birthdate="2012-05-15" gender="M" nation="BRA" license="369258" swrid="5588942" athleteid="1283" externalid="369258">
              <RESULTS>
                <RESULT eventid="1101" points="359" swimtime="00:00:31.33" resultid="1284" heatid="2378" lane="4" entrytime="00:00:32.62" entrycourse="LCM" />
                <RESULT eventid="1073" points="311" swimtime="00:02:48.14" resultid="1285" heatid="2341" lane="4" entrytime="00:02:49.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="302" swimtime="00:01:16.89" resultid="1286" heatid="2420" lane="4" entrytime="00:01:19.28" entrycourse="LCM" />
                <RESULT eventid="1117" status="DNS" swimtime="00:00:00.00" resultid="1287" heatid="2395" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Toscani Kim" birthdate="2013-02-15" gender="F" nation="BRA" license="372683" swrid="5588939" athleteid="1378" externalid="372683">
              <RESULTS>
                <RESULT eventid="1098" points="256" swimtime="00:00:38.46" resultid="1379" heatid="2373" lane="5" entrytime="00:00:42.62" entrycourse="LCM" />
                <RESULT eventid="1070" points="320" swimtime="00:03:04.38" resultid="1380" heatid="2337" lane="5" entrytime="00:03:06.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="313" swimtime="00:05:46.60" resultid="1381" heatid="2392" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.02" />
                    <SPLIT distance="200" swimtime="00:02:49.06" />
                    <SPLIT distance="300" swimtime="00:04:18.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="302" swimtime="00:00:43.42" resultid="1382" heatid="2433" lane="5" entrytime="00:00:43.19" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcela" lastname="Tallao Benke" birthdate="2014-10-07" gender="F" nation="BRA" license="382075" swrid="5602586" athleteid="1514" externalid="382075">
              <RESULTS>
                <RESULT eventid="1092" points="234" swimtime="00:00:39.60" resultid="1515" heatid="2367" lane="5" entrytime="00:00:39.97" entrycourse="LCM" />
                <RESULT eventid="1064" points="277" swimtime="00:02:52.96" resultid="1516" heatid="2330" lane="4" entrytime="00:02:55.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="321" swimtime="00:00:34.47" resultid="1517" heatid="2424" lane="5" entrytime="00:00:34.88" entrycourse="LCM" />
                <RESULT eventid="1108" points="286" swimtime="00:03:11.39" resultid="1518" heatid="2385" lane="4" entrytime="00:03:15.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Gois Nogueira" birthdate="2014-03-11" gender="F" nation="BRA" license="393258" swrid="5616443" athleteid="1624" externalid="393258">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="1625" heatid="2365" lane="2" entrytime="00:00:56.96" entrycourse="LCM" />
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="1626" heatid="2348" lane="1" entrytime="00:00:53.22" entrycourse="LCM" />
                <RESULT eventid="1136" status="DNS" swimtime="00:00:00.00" resultid="1627" heatid="2423" lane="1" entrytime="00:00:42.10" entrycourse="LCM" />
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="1628" heatid="2404" lane="2" entrytime="00:00:50.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Menezes" birthdate="2015-07-28" gender="F" nation="BRA" license="412898" swrid="5755339" athleteid="1835" externalid="412898">
              <RESULTS>
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="1836" heatid="2345" lane="5" />
                <RESULT eventid="1136" points="125" swimtime="00:00:47.18" resultid="1837" heatid="2422" lane="7" entrytime="00:00:47.17" entrycourse="LCM" />
                <RESULT eventid="1124" points="124" swimtime="00:00:53.74" resultid="1838" heatid="2403" lane="6" entrytime="00:00:57.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="De Moraes" birthdate="2014-09-18" gender="M" nation="BRA" license="391024" swrid="5602529" athleteid="1589" externalid="391024">
              <RESULTS>
                <RESULT eventid="1095" points="171" swimtime="00:00:40.08" resultid="1590" heatid="2370" lane="3" entrytime="00:00:40.53" entrycourse="LCM" />
                <RESULT eventid="1067" points="224" swimtime="00:02:47.77" resultid="1591" heatid="2334" lane="5" entrytime="00:02:57.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="159" swimtime="00:03:30.13" resultid="1592" heatid="2389" lane="6" entrytime="00:03:29.31" entrycourse="LCM" />
                <RESULT eventid="1139" points="264" swimtime="00:00:32.57" resultid="1593" heatid="2429" lane="5" entrytime="00:00:33.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Da Cunha Souza" birthdate="2013-09-17" gender="M" nation="BRA" license="376975" swrid="5588618" athleteid="1425" externalid="376975">
              <RESULTS>
                <RESULT eventid="1101" points="126" swimtime="00:00:44.32" resultid="1426" heatid="2376" lane="4" entrytime="00:00:44.64" entrycourse="LCM" />
                <RESULT eventid="1089" points="193" swimtime="00:01:21.05" resultid="1427" heatid="2362" lane="5" entrytime="00:01:22.34" entrycourse="LCM" />
                <RESULT eventid="1117" points="186" swimtime="00:06:25.40" resultid="1428" heatid="2396" lane="6" entrytime="00:06:34.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.38" />
                    <SPLIT distance="200" swimtime="00:03:12.40" />
                    <SPLIT distance="300" swimtime="00:04:50.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="126" swimtime="00:00:51.70" resultid="1429" heatid="2436" lane="7" entrytime="00:00:55.89" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Coelho Ghignone" birthdate="2015-01-05" gender="M" nation="BRA" license="410201" swrid="5740006" athleteid="1793" externalid="410201">
              <RESULTS>
                <RESULT eventid="1095" points="75" swimtime="00:00:52.62" resultid="1794" heatid="2369" lane="1" entrytime="00:00:56.47" entrycourse="LCM" />
                <RESULT eventid="1067" points="119" swimtime="00:03:27.00" resultid="1795" heatid="2332" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="125" swimtime="00:00:47.05" resultid="1796" heatid="2410" lane="8" entrytime="00:00:46.72" entrycourse="LCM" />
                <RESULT eventid="1111" points="110" swimtime="00:03:57.46" resultid="1797" heatid="2387" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:54.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Cury Abreu" birthdate="2013-05-17" gender="F" nation="BRA" license="376974" swrid="5588614" athleteid="1420" externalid="376974">
              <RESULTS>
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="1421" heatid="2373" lane="8" entrytime="00:00:50.10" entrycourse="LCM" />
                <RESULT eventid="1086" status="DNS" swimtime="00:00:00.00" resultid="1422" heatid="2357" lane="5" entrytime="00:01:17.65" entrycourse="LCM" />
                <RESULT eventid="1130" points="273" swimtime="00:01:28.34" resultid="1423" heatid="2415" lane="8" entrytime="00:01:28.64" entrycourse="LCM" />
                <RESULT eventid="1114" points="284" swimtime="00:05:58.09" resultid="1424" heatid="2390" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.84" />
                    <SPLIT distance="200" swimtime="00:02:55.95" />
                    <SPLIT distance="300" swimtime="00:04:29.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alan" lastname="Batista Grise" birthdate="2014-03-27" gender="M" nation="BRA" license="391007" swrid="5602513" athleteid="1539" externalid="391007">
              <RESULTS>
                <RESULT eventid="1095" points="40" swimtime="00:01:04.87" resultid="1540" heatid="2368" lane="6" />
                <RESULT eventid="1083" points="87" swimtime="00:00:58.47" resultid="1541" heatid="2350" lane="5" entrytime="00:01:00.33" entrycourse="LCM" />
                <RESULT eventid="1127" points="83" swimtime="00:00:53.98" resultid="1542" heatid="2408" lane="4" entrytime="00:00:56.30" entrycourse="LCM" />
                <RESULT eventid="1139" points="99" swimtime="00:00:45.07" resultid="1543" heatid="2426" lane="6" entrytime="00:00:48.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Cavalca Petraglia" birthdate="2015-08-06" gender="M" nation="BRA" license="397275" swrid="5641757" athleteid="1678" externalid="397275">
              <RESULTS>
                <RESULT eventid="1095" points="70" swimtime="00:00:54.01" resultid="1679" heatid="2369" lane="2" entrytime="00:00:54.37" entrycourse="LCM" />
                <RESULT eventid="1067" points="94" swimtime="00:03:43.67" resultid="1680" heatid="2331" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="96" swimtime="00:04:08.35" resultid="1681" heatid="2388" lane="7" entrytime="00:04:19.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:03.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="100" swimtime="00:00:45.02" resultid="1682" heatid="2427" lane="1" entrytime="00:00:45.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Salomao" birthdate="2012-05-07" gender="M" nation="BRA" license="369261" swrid="5602581" athleteid="1293" externalid="369261">
              <RESULTS>
                <RESULT eventid="1101" points="233" swimtime="00:00:36.14" resultid="1294" heatid="2378" lane="1" entrytime="00:00:37.73" entrycourse="LCM" />
                <RESULT eventid="1073" points="246" swimtime="00:03:01.91" resultid="1295" heatid="2339" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="1296" heatid="2416" lane="4" />
                <RESULT eventid="1117" status="DNS" swimtime="00:00:00.00" resultid="1297" heatid="2397" lane="5" entrytime="00:05:28.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Taborda Ribas" birthdate="2015-12-30" gender="M" nation="BRA" license="406748" swrid="5717299" athleteid="1733" externalid="406748">
              <RESULTS>
                <RESULT comment="SW 7.4 - Movimentos das pernas não simultâneos.  (Horário: 11:08)" eventid="1083" status="DSQ" swimtime="00:01:09.95" resultid="1734" heatid="2349" lane="7" />
                <RESULT eventid="1067" points="71" swimtime="00:04:05.32" resultid="1735" heatid="2332" lane="5" entrytime="00:04:09.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="66" swimtime="00:00:58.26" resultid="1736" heatid="2408" lane="6" entrytime="00:00:57.77" entrycourse="LCM" />
                <RESULT eventid="1111" points="62" swimtime="00:04:47.56" resultid="1737" heatid="2387" lane="5" entrytime="00:04:58.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:15.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maya" lastname="Assahida Moreria" birthdate="2014-02-24" gender="F" nation="BRA" license="391020" swrid="5602512" athleteid="1574" externalid="391020">
              <RESULTS>
                <RESULT eventid="1092" points="161" swimtime="00:00:44.88" resultid="1575" heatid="2367" lane="7" entrytime="00:00:46.48" entrycourse="LCM" />
                <RESULT eventid="1064" points="238" swimtime="00:03:01.91" resultid="1576" heatid="2330" lane="5" entrytime="00:03:15.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="262" swimtime="00:00:36.86" resultid="1577" heatid="2423" lane="6" entrytime="00:00:41.12" entrycourse="LCM" />
                <RESULT eventid="1108" points="208" swimtime="00:03:32.63" resultid="1578" heatid="2385" lane="3" entrytime="00:03:44.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enrico" lastname="Gubert Camargo" birthdate="2016-02-12" gender="M" nation="BRA" license="417119" athleteid="1875" externalid="417119">
              <RESULTS>
                <RESULT eventid="1122" points="57" swimtime="00:00:54.19" resultid="1876" heatid="2400" lane="4" />
                <RESULT eventid="1106" points="60" swimtime="00:01:05.99" resultid="1877" heatid="2381" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Crescente Rastelli" birthdate="2015-01-21" gender="M" nation="BRA" license="416673" athleteid="1872" externalid="416673">
              <RESULTS>
                <RESULT eventid="1127" points="92" swimtime="00:00:52.09" resultid="1873" heatid="2406" lane="3" />
                <RESULT eventid="1139" points="99" swimtime="00:00:45.14" resultid="1874" heatid="2425" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Ruschka Druszcz" birthdate="2016-05-09" gender="F" nation="BRA" license="412025" swrid="5740018" athleteid="1825" externalid="412025">
              <RESULTS>
                <RESULT eventid="1060" status="DNS" swimtime="00:00:00.00" resultid="1826" heatid="2326" lane="5" />
                <RESULT eventid="1076" points="89" swimtime="00:00:59.98" resultid="1827" heatid="2343" lane="5" entrytime="00:01:00.99" entrycourse="LCM" />
                <RESULT eventid="1120" points="87" swimtime="00:00:53.15" resultid="1828" heatid="2399" lane="5" entrytime="00:00:52.02" entrycourse="LCM" />
                <RESULT eventid="1104" points="105" swimtime="00:01:01.80" resultid="1829" heatid="2380" lane="3" entrytime="00:01:06.26" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Szpak Zraik" birthdate="2015-04-10" gender="M" nation="BRA" license="393259" swrid="5616451" athleteid="1629" externalid="393259">
              <RESULTS>
                <RESULT eventid="1083" status="DNS" swimtime="00:00:00.00" resultid="1630" heatid="2352" lane="3" entrytime="00:00:48.23" entrycourse="LCM" />
                <RESULT eventid="1067" status="DNS" swimtime="00:00:00.00" resultid="1631" heatid="2333" lane="4" entrytime="00:03:40.19" entrycourse="LCM" />
                <RESULT eventid="1111" status="DNS" swimtime="00:00:00.00" resultid="1632" heatid="2389" lane="8" entrytime="00:04:01.60" entrycourse="LCM" />
                <RESULT eventid="1139" status="DNS" swimtime="00:00:00.00" resultid="1633" heatid="2427" lane="5" entrytime="00:00:40.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enrico" lastname="Hallage Bianchini" birthdate="2014-02-27" gender="M" nation="BRA" license="397164" swrid="5661348" athleteid="1668" externalid="397164">
              <RESULTS>
                <RESULT eventid="1095" points="142" swimtime="00:00:42.62" resultid="1669" heatid="2369" lane="4" entrytime="00:00:43.86" entrycourse="LCM" />
                <RESULT eventid="1067" points="202" swimtime="00:02:53.57" resultid="1670" heatid="2333" lane="6" entrytime="00:03:56.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="165" swimtime="00:03:27.49" resultid="1671" heatid="2389" lane="1" entrytime="00:03:49.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="213" swimtime="00:00:35.01" resultid="1672" heatid="2429" lane="2" entrytime="00:00:35.44" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Portes Fabiane" birthdate="2012-12-28" gender="M" nation="BRA" license="376983" swrid="5588864" athleteid="1450" externalid="376983">
              <RESULTS>
                <RESULT eventid="1101" points="54" swimtime="00:00:58.91" resultid="1451" heatid="2375" lane="4" />
                <RESULT eventid="1089" points="111" swimtime="00:01:37.40" resultid="1452" heatid="2360" lane="6" entrytime="00:01:48.01" entrycourse="LCM" />
                <RESULT eventid="1133" points="96" swimtime="00:01:52.45" resultid="1453" heatid="2419" lane="1" entrytime="00:01:59.49" entrycourse="LCM" />
                <RESULT eventid="1145" points="80" swimtime="00:00:59.99" resultid="1454" heatid="2436" lane="1" entrytime="00:01:02.03" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Alice Palhano" birthdate="2016-04-06" gender="F" nation="BRA" license="412015" swrid="5740004" athleteid="1818" externalid="412015">
              <RESULTS>
                <RESULT eventid="1076" points="48" swimtime="00:01:13.62" resultid="1819" heatid="2342" lane="4" entrytime="00:01:13.51" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olavo" lastname="Valduga Artigas" birthdate="2012-06-26" gender="M" nation="BRA" license="369270" swrid="5588941" athleteid="1318" externalid="369270">
              <RESULTS>
                <RESULT eventid="1089" points="186" swimtime="00:01:21.97" resultid="1319" heatid="2362" lane="8" entrytime="00:01:25.88" entrycourse="LCM" />
                <RESULT eventid="1073" points="198" swimtime="00:03:15.54" resultid="1320" heatid="2341" lane="8" entrytime="00:03:09.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" status="DNS" swimtime="00:00:00.00" resultid="1321" heatid="2396" lane="8" />
                <RESULT eventid="1145" status="DNS" swimtime="00:00:00.00" resultid="1322" heatid="2438" lane="8" entrytime="00:00:45.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Baptistella" birthdate="2013-01-23" gender="M" nation="BRA" license="391152" swrid="5602545" athleteid="1614" externalid="391152">
              <RESULTS>
                <RESULT eventid="1089" points="242" swimtime="00:01:15.10" resultid="1615" heatid="2362" lane="7" entrytime="00:01:24.28" entrycourse="LCM" />
                <RESULT eventid="1073" points="214" swimtime="00:03:10.45" resultid="1616" heatid="2340" lane="2" entrytime="00:03:11.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="212" swimtime="00:01:26.41" resultid="1617" heatid="2419" lane="5" entrytime="00:01:30.64" entrycourse="LCM" />
                <RESULT eventid="1117" points="232" swimtime="00:05:58.14" resultid="1618" heatid="2395" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Morais Shibata" birthdate="2014-02-09" gender="M" nation="BRA" license="391018" swrid="5602561" athleteid="1564" externalid="391018">
              <RESULTS>
                <RESULT eventid="1083" points="132" swimtime="00:00:50.84" resultid="1565" heatid="2351" lane="4" entrytime="00:00:52.29" entrycourse="LCM" />
                <RESULT eventid="1067" points="136" swimtime="00:03:18.16" resultid="1566" heatid="2333" lane="2" entrytime="00:03:57.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="151" swimtime="00:00:44.14" resultid="1567" heatid="2410" lane="1" entrytime="00:00:45.33" entrycourse="LCM" />
                <RESULT eventid="1111" points="139" swimtime="00:03:40.01" resultid="1568" heatid="2388" lane="6" entrytime="00:04:17.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Mayer Paludetto" birthdate="2012-10-30" gender="F" nation="BRA" license="369264" swrid="5588811" athleteid="1303" externalid="369264">
              <RESULTS>
                <RESULT eventid="1086" points="444" swimtime="00:01:07.77" resultid="1304" heatid="2358" lane="2" entrytime="00:01:13.49" entrycourse="LCM" />
                <RESULT eventid="1070" points="413" swimtime="00:02:49.34" resultid="1305" heatid="2338" lane="4" entrytime="00:02:50.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="347" swimtime="00:01:21.55" resultid="1306" heatid="2413" lane="6" />
                <RESULT eventid="1114" points="465" swimtime="00:05:03.81" resultid="1307" heatid="2393" lane="2" entrytime="00:05:16.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                    <SPLIT distance="200" swimtime="00:02:32.00" />
                    <SPLIT distance="300" swimtime="00:03:49.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Garcia" birthdate="2015-10-26" gender="M" nation="BRA" license="406967" swrid="5717271" athleteid="1778" externalid="406967">
              <RESULTS>
                <RESULT eventid="1083" points="22" swimtime="00:01:32.25" resultid="1779" heatid="2349" lane="3" entrytime="00:01:27.24" entrycourse="LCM" />
                <RESULT eventid="1067" points="52" swimtime="00:04:32.76" resultid="1780" heatid="2332" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:15.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="46" swimtime="00:01:05.64" resultid="1781" heatid="2407" lane="4" entrytime="00:01:03.30" entrycourse="LCM" />
                <RESULT eventid="1139" points="34" swimtime="00:01:04.38" resultid="1782" heatid="2425" lane="4" entrytime="00:01:08.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Cabrini Vieira" birthdate="2012-02-11" gender="F" nation="BRA" license="376961" swrid="5588571" athleteid="1393" externalid="376961">
              <RESULTS>
                <RESULT eventid="1086" points="446" swimtime="00:01:07.65" resultid="1394" heatid="2353" lane="4" />
                <RESULT eventid="1070" points="358" swimtime="00:02:57.48" resultid="1395" heatid="2338" lane="6" entrytime="00:02:59.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="331" swimtime="00:01:22.87" resultid="1396" heatid="2415" lane="5" entrytime="00:01:17.59" entrycourse="LCM" />
                <RESULT eventid="1114" points="434" swimtime="00:05:10.67" resultid="1397" heatid="2393" lane="5" entrytime="00:05:09.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.56" />
                    <SPLIT distance="200" swimtime="00:02:34.15" />
                    <SPLIT distance="300" swimtime="00:03:55.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Alzamora Calado" birthdate="2013-04-26" gender="F" nation="BRA" license="376960" swrid="5588522" athleteid="1388" externalid="376960">
              <RESULTS>
                <RESULT eventid="1086" points="336" swimtime="00:01:14.35" resultid="1389" heatid="2358" lane="8" entrytime="00:01:16.15" entrycourse="LCM" />
                <RESULT eventid="1070" points="289" swimtime="00:03:10.63" resultid="1390" heatid="2337" lane="1" entrytime="00:03:17.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="304" swimtime="00:05:49.71" resultid="1391" heatid="2390" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.10" />
                    <SPLIT distance="200" swimtime="00:02:52.67" />
                    <SPLIT distance="300" swimtime="00:04:24.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="310" swimtime="00:00:43.05" resultid="1392" heatid="2433" lane="8" entrytime="00:00:46.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luigi" lastname="Antoniuk Paganini" birthdate="2014-11-13" gender="M" nation="BRA" license="382127" swrid="5602509" athleteid="1529" externalid="382127">
              <RESULTS>
                <RESULT eventid="1095" points="153" swimtime="00:00:41.63" resultid="1530" heatid="2370" lane="7" entrytime="00:00:42.45" entrycourse="LCM" />
                <RESULT eventid="1067" points="186" swimtime="00:02:58.63" resultid="1531" heatid="2334" lane="8" entrytime="00:03:23.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="208" swimtime="00:00:39.73" resultid="1532" heatid="2410" lane="3" entrytime="00:00:40.90" entrycourse="LCM" />
                <RESULT eventid="1111" points="163" swimtime="00:03:28.33" resultid="1533" heatid="2388" lane="3" entrytime="00:04:15.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Albuquerque" birthdate="2012-11-16" gender="F" nation="BRA" license="369281" swrid="5602506" athleteid="1358" externalid="369281">
              <RESULTS>
                <RESULT eventid="1098" points="273" swimtime="00:00:37.64" resultid="1359" heatid="2374" lane="8" entrytime="00:00:41.49" entrycourse="LCM" />
                <RESULT eventid="1070" points="368" swimtime="00:02:55.95" resultid="1360" heatid="2338" lane="2" entrytime="00:02:59.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="369" swimtime="00:05:28.09" resultid="1361" heatid="2393" lane="8" entrytime="00:05:39.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.39" />
                    <SPLIT distance="200" swimtime="00:02:42.63" />
                    <SPLIT distance="300" swimtime="00:04:07.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="305" swimtime="00:00:43.28" resultid="1362" heatid="2431" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Moreira Pasqual" birthdate="2014-07-09" gender="M" nation="BRA" license="382125" swrid="5602562" athleteid="1524" externalid="382125">
              <RESULTS>
                <RESULT eventid="1095" points="164" swimtime="00:00:40.68" resultid="1525" heatid="2370" lane="6" entrytime="00:00:40.70" entrycourse="LCM" />
                <RESULT eventid="1067" points="175" swimtime="00:03:02.30" resultid="1526" heatid="2333" lane="5" entrytime="00:03:42.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="171" swimtime="00:03:25.24" resultid="1527" heatid="2388" lane="4" entrytime="00:04:12.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="201" swimtime="00:00:35.69" resultid="1528" heatid="2429" lane="8" entrytime="00:00:36.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Steven" lastname="Matheussi Viana E Silva" birthdate="2012-05-03" gender="M" nation="BRA" license="376986" swrid="5588810" athleteid="1494" externalid="376986">
              <RESULTS>
                <RESULT eventid="1101" points="213" swimtime="00:00:37.26" resultid="1495" heatid="2378" lane="2" entrytime="00:00:37.30" entrycourse="LCM" />
                <RESULT eventid="1089" points="294" swimtime="00:01:10.45" resultid="1496" heatid="2359" lane="3" />
                <RESULT eventid="1117" points="282" swimtime="00:05:35.54" resultid="1497" heatid="2396" lane="4" entrytime="00:05:56.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.83" />
                    <SPLIT distance="200" swimtime="00:02:47.49" />
                    <SPLIT distance="300" swimtime="00:04:13.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" status="DNS" swimtime="00:00:00.00" resultid="1498" heatid="2438" lane="6" entrytime="00:00:41.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Pens Correa" birthdate="2015-11-27" gender="M" nation="BRA" license="393262" swrid="5616449" athleteid="1643" externalid="393262">
              <RESULTS>
                <RESULT eventid="1095" points="183" swimtime="00:00:39.20" resultid="1644" heatid="2370" lane="5" entrytime="00:00:38.70" entrycourse="LCM" />
                <RESULT eventid="1067" points="203" swimtime="00:02:53.54" resultid="1645" heatid="2334" lane="3" entrytime="00:03:01.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="213" swimtime="00:03:10.62" resultid="1646" heatid="2389" lane="3" entrytime="00:03:27.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="213" swimtime="00:00:34.99" resultid="1647" heatid="2429" lane="6" entrytime="00:00:34.96" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Xavier Jardim" birthdate="2012-01-23" gender="M" nation="BRA" license="369259" swrid="5641781" athleteid="1288" externalid="369259">
              <RESULTS>
                <RESULT eventid="1101" points="192" swimtime="00:00:38.57" resultid="1289" heatid="2377" lane="4" entrytime="00:00:39.71" entrycourse="LCM" />
                <RESULT eventid="1089" points="286" swimtime="00:01:11.10" resultid="1290" heatid="2364" lane="7" entrytime="00:01:10.67" entrycourse="LCM" />
                <RESULT eventid="1133" points="208" swimtime="00:01:27.07" resultid="1291" heatid="2420" lane="2" entrytime="00:01:24.67" entrycourse="LCM" />
                <RESULT eventid="1117" points="265" swimtime="00:05:42.28" resultid="1292" heatid="2395" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.96" />
                    <SPLIT distance="200" swimtime="00:02:50.65" />
                    <SPLIT distance="300" swimtime="00:04:19.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Guimaraes Mesquita" birthdate="2013-12-30" gender="F" nation="BRA" license="391027" swrid="5602544" athleteid="1604" externalid="391027">
              <RESULTS>
                <RESULT eventid="1086" points="189" swimtime="00:01:30.05" resultid="1605" heatid="2356" lane="7" entrytime="00:01:31.04" entrycourse="LCM" />
                <RESULT eventid="1070" points="182" swimtime="00:03:42.36" resultid="1606" heatid="2336" lane="6" entrytime="00:03:38.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:57.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="194" swimtime="00:06:45.92" resultid="1607" heatid="2391" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.65" />
                    <SPLIT distance="200" swimtime="00:03:23.87" />
                    <SPLIT distance="300" swimtime="00:05:08.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="148" swimtime="00:00:55.04" resultid="1608" heatid="2432" lane="2" entrytime="00:00:54.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Pisani Ferreira" birthdate="2014-01-26" gender="M" nation="BRA" license="391017" swrid="5602570" athleteid="1559" externalid="391017">
              <RESULTS>
                <RESULT eventid="1083" points="151" swimtime="00:00:48.63" resultid="1560" heatid="2352" lane="7" entrytime="00:00:50.61" entrycourse="LCM" />
                <RESULT eventid="1067" points="102" swimtime="00:03:37.99" resultid="1561" heatid="2333" lane="8" entrytime="00:04:05.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="116" swimtime="00:03:53.54" resultid="1562" heatid="2388" lane="1" entrytime="00:04:27.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:59.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="129" swimtime="00:00:41.32" resultid="1563" heatid="2427" lane="4" entrytime="00:00:40.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Zagonel Krempel" birthdate="2015-07-27" gender="F" nation="BRA" license="406962" swrid="5717305" athleteid="1768" externalid="406962">
              <RESULTS>
                <RESULT eventid="1080" points="94" swimtime="00:01:03.95" resultid="1769" heatid="2346" lane="5" entrytime="00:01:02.90" entrycourse="LCM" />
                <RESULT eventid="1064" points="114" swimtime="00:03:52.08" resultid="1770" heatid="2327" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="128" swimtime="00:00:46.77" resultid="1771" heatid="2422" lane="1" entrytime="00:00:47.52" entrycourse="LCM" />
                <RESULT comment="SW 8.3 - Movimento alternado das pernas ou pés.  (Horário: 15:54), (Medley Individual, Borboleta)." eventid="1108" status="DSQ" swimtime="00:04:19.90" resultid="1772" heatid="2382" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:11.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Cabrera Cirino Dos Santos" birthdate="2013-03-30" gender="M" nation="BRA" license="376990" swrid="5588570" athleteid="1479" externalid="376990">
              <RESULTS>
                <RESULT comment="SW 8.3 - Movimento alternado das pernas ou pés.  (Horário: 12:16)" eventid="1101" status="DSQ" swimtime="00:00:42.99" resultid="1480" heatid="2377" lane="8" entrytime="00:00:43.87" entrycourse="LCM" />
                <RESULT eventid="1089" points="218" swimtime="00:01:17.76" resultid="1481" heatid="2363" lane="8" entrytime="00:01:20.98" entrycourse="LCM" />
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="1482" heatid="2418" lane="8" />
                <RESULT eventid="1117" status="DNS" swimtime="00:00:00.00" resultid="1483" heatid="2396" lane="5" entrytime="00:06:00.28" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Szpak De Vasconcelos" birthdate="2012-06-29" gender="M" nation="BRA" license="369271" swrid="5588928" athleteid="1323" externalid="369271">
              <RESULTS>
                <RESULT eventid="1089" points="341" swimtime="00:01:07.07" resultid="1324" heatid="2364" lane="4" entrytime="00:01:06.90" entrycourse="LCM" />
                <RESULT eventid="1073" points="304" swimtime="00:02:49.42" resultid="1325" heatid="2341" lane="5" entrytime="00:02:50.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="322" swimtime="00:05:20.85" resultid="1326" heatid="2395" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.58" />
                    <SPLIT distance="200" swimtime="00:02:38.17" />
                    <SPLIT distance="300" swimtime="00:04:00.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="325" swimtime="00:00:37.72" resultid="1327" heatid="2438" lane="4" entrytime="00:00:38.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Toscani Kim" birthdate="2015-10-02" gender="F" nation="BRA" license="397276" swrid="5641778" athleteid="1683" externalid="397276">
              <RESULTS>
                <RESULT eventid="1080" points="183" swimtime="00:00:51.34" resultid="1684" heatid="2348" lane="6" entrytime="00:00:50.80" entrycourse="LCM" />
                <RESULT eventid="1064" points="171" swimtime="00:03:23.27" resultid="1685" heatid="2330" lane="8" entrytime="00:03:36.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="200" swimtime="00:00:45.88" resultid="1686" heatid="2404" lane="7" entrytime="00:00:51.48" entrycourse="LCM" />
                <RESULT eventid="1108" points="195" swimtime="00:03:37.37" resultid="1687" heatid="2385" lane="1" entrytime="00:03:54.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Kraemer Geremia" birthdate="2013-08-16" gender="M" nation="BRA" license="377041" swrid="5588762" athleteid="1465" externalid="377041">
              <RESULTS>
                <RESULT eventid="1101" points="203" swimtime="00:00:37.84" resultid="1466" heatid="2378" lane="8" entrytime="00:00:39.11" entrycourse="LCM" />
                <RESULT eventid="1089" points="283" swimtime="00:01:11.30" resultid="1467" heatid="2364" lane="1" entrytime="00:01:14.54" entrycourse="LCM" />
                <RESULT eventid="1133" points="215" swimtime="00:01:26.08" resultid="1468" heatid="2417" lane="3" />
                <RESULT eventid="1117" points="257" swimtime="00:05:45.79" resultid="1469" heatid="2396" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.41" />
                    <SPLIT distance="200" swimtime="00:02:53.60" />
                    <SPLIT distance="300" swimtime="00:04:22.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Saporiti Salvi" birthdate="2013-06-28" gender="M" nation="BRA" license="377032" swrid="5588896" athleteid="1460" externalid="377032">
              <RESULTS>
                <RESULT eventid="1101" points="186" swimtime="00:00:38.99" resultid="1461" heatid="2377" lane="1" entrytime="00:00:43.63" entrycourse="LCM" />
                <RESULT eventid="1073" points="224" swimtime="00:03:07.49" resultid="1462" heatid="2340" lane="4" entrytime="00:03:10.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="244" swimtime="00:05:51.95" resultid="1463" heatid="2396" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:57.23" />
                    <SPLIT distance="300" swimtime="00:04:27.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="138" swimtime="00:00:50.11" resultid="1464" heatid="2437" lane="1" entrytime="00:00:51.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Bernardi Pedrosa" birthdate="2013-03-09" gender="F" nation="BRA" license="376977" swrid="5588551" athleteid="1430" externalid="376977">
              <RESULTS>
                <RESULT eventid="1086" points="265" swimtime="00:01:20.41" resultid="1431" heatid="2357" lane="1" entrytime="00:01:21.00" entrycourse="LCM" />
                <RESULT eventid="1070" points="233" swimtime="00:03:24.82" resultid="1432" heatid="2336" lane="5" entrytime="00:03:29.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="230" swimtime="00:01:33.46" resultid="1433" heatid="2414" lane="5" entrytime="00:01:31.64" entrycourse="LCM" />
                <RESULT eventid="1114" points="271" swimtime="00:06:03.53" resultid="1434" heatid="2391" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.83" />
                    <SPLIT distance="200" swimtime="00:03:01.96" />
                    <SPLIT distance="300" swimtime="00:04:36.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cecilia Carvalho" birthdate="2014-10-30" gender="F" nation="BRA" license="391021" swrid="5602525" athleteid="1579" externalid="391021">
              <RESULTS>
                <RESULT eventid="1092" points="74" swimtime="00:00:58.05" resultid="1580" heatid="2365" lane="7" entrytime="00:00:57.32" entrycourse="LCM" />
                <RESULT eventid="1064" points="151" swimtime="00:03:31.51" resultid="1581" heatid="2328" lane="5" entrytime="00:04:17.55" entrycourse="LCM" />
                <RESULT eventid="1136" status="DNS" swimtime="00:00:00.00" resultid="1582" heatid="2422" lane="6" entrytime="00:00:44.16" entrycourse="LCM" />
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="1583" heatid="2384" lane="6" entrytime="00:04:54.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Hadad" birthdate="2015-09-09" gender="M" nation="BRA" license="406740" swrid="5717272" athleteid="1718" externalid="406740">
              <RESULTS>
                <RESULT eventid="1083" points="56" swimtime="00:01:07.82" resultid="1719" heatid="2350" lane="8" entrytime="00:01:05.79" entrycourse="LCM" />
                <RESULT eventid="1067" points="80" swimtime="00:03:56.07" resultid="1720" heatid="2333" lane="1" entrytime="00:04:04.02" entrycourse="LCM" />
                <RESULT eventid="1127" points="73" swimtime="00:00:56.11" resultid="1721" heatid="2408" lane="7" entrytime="00:00:59.70" entrycourse="LCM" />
                <RESULT eventid="1111" points="74" swimtime="00:04:30.84" resultid="1722" heatid="2387" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Albuquerque" birthdate="2012-08-17" gender="F" nation="BRA" license="369275" swrid="5602507" athleteid="1333" externalid="369275">
              <RESULTS>
                <RESULT eventid="1098" points="264" swimtime="00:00:38.05" resultid="1334" heatid="2374" lane="6" entrytime="00:00:38.73" entrycourse="LCM" />
                <RESULT eventid="1070" points="274" swimtime="00:03:13.95" resultid="1335" heatid="2337" lane="3" entrytime="00:03:06.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="189" swimtime="00:01:39.84" resultid="1336" heatid="2413" lane="2" />
                <RESULT eventid="1142" points="437" swimtime="00:00:38.41" resultid="1337" heatid="2433" lane="4" entrytime="00:00:39.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Shwetz Clivatti" birthdate="2015-03-05" gender="M" nation="BRA" license="406963" swrid="5717297" athleteid="1773" externalid="406963">
              <RESULTS>
                <RESULT eventid="1083" points="46" swimtime="00:01:12.33" resultid="1774" heatid="2349" lane="4" entrytime="00:01:09.43" entrycourse="LCM" />
                <RESULT eventid="1067" points="55" swimtime="00:04:27.70" resultid="1775" heatid="2331" lane="7" />
                <RESULT eventid="1127" points="56" swimtime="00:01:01.35" resultid="1776" heatid="2408" lane="8" entrytime="00:01:02.66" entrycourse="LCM" />
                <RESULT eventid="1139" points="47" swimtime="00:00:57.86" resultid="1777" heatid="2426" lane="7" entrytime="00:00:55.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Vianna Almeida" birthdate="2014-12-16" gender="M" nation="BRA" license="410292" swrid="5740019" athleteid="1798" externalid="410292">
              <RESULTS>
                <RESULT eventid="1083" points="114" swimtime="00:00:53.38" resultid="1799" heatid="2351" lane="2" entrytime="00:00:54.16" entrycourse="LCM" />
                <RESULT eventid="1067" points="112" swimtime="00:03:31.46" resultid="1800" heatid="2332" lane="4" entrytime="00:04:07.62" entrycourse="LCM" />
                <RESULT eventid="1111" points="102" swimtime="00:04:03.77" resultid="1801" heatid="2387" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:03.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="131" swimtime="00:00:41.17" resultid="1802" heatid="2427" lane="2" entrytime="00:00:43.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Petraglia" birthdate="2012-03-28" gender="M" nation="BRA" license="369282" swrid="5602569" athleteid="1363" externalid="369282">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="1364" heatid="2364" lane="8" entrytime="00:01:15.62" entrycourse="LCM" />
                <RESULT eventid="1073" status="DNS" swimtime="00:00:00.00" resultid="1365" heatid="2340" lane="1" entrytime="00:03:15.85" entrycourse="LCM" />
                <RESULT eventid="1117" status="DNS" swimtime="00:00:00.00" resultid="1366" heatid="2397" lane="6" entrytime="00:05:35.54" entrycourse="LCM" />
                <RESULT eventid="1145" status="DNS" swimtime="00:00:00.00" resultid="1367" heatid="2438" lane="1" entrytime="00:00:45.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Pisani Ferreira" birthdate="2012-08-06" gender="F" nation="BRA" license="376985" swrid="5588862" athleteid="1499" externalid="376985">
              <RESULTS>
                <RESULT eventid="1086" points="199" swimtime="00:01:28.50" resultid="1500" heatid="2356" lane="2" entrytime="00:01:30.94" entrycourse="LCM" />
                <RESULT eventid="1070" points="180" swimtime="00:03:43.04" resultid="1501" heatid="2336" lane="2" entrytime="00:03:39.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="148" swimtime="00:01:48.30" resultid="1502" heatid="2412" lane="6" />
                <RESULT eventid="1142" points="222" swimtime="00:00:48.10" resultid="1503" heatid="2432" lane="3" entrytime="00:00:47.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giuliana" lastname="Sovierzoski Ferreira" birthdate="2015-01-20" gender="F" nation="BRA" license="397168" swrid="5641776" athleteid="1673" externalid="397168">
              <RESULTS>
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="1674" heatid="2348" lane="7" entrytime="00:00:53.15" entrycourse="LCM" />
                <RESULT eventid="1064" status="DNS" swimtime="00:00:00.00" resultid="1675" heatid="2328" lane="2" />
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="1676" heatid="2403" lane="8" entrytime="00:00:59.15" entrycourse="LCM" />
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="1677" heatid="2384" lane="3" entrytime="00:04:45.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Stramandinoli Zanicotti" birthdate="2013-06-18" gender="F" nation="BRA" license="376967" swrid="5588924" athleteid="1407" externalid="376967">
              <RESULTS>
                <RESULT eventid="1086" points="162" swimtime="00:01:34.82" resultid="1408" heatid="2355" lane="2" entrytime="00:01:53.85" entrycourse="LCM" />
                <RESULT eventid="1070" points="146" swimtime="00:03:59.25" resultid="1409" heatid="2336" lane="1" entrytime="00:04:05.23" entrycourse="LCM" />
                <RESULT eventid="1114" points="137" swimtime="00:07:35.81" resultid="1410" heatid="2390" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.20" />
                    <SPLIT distance="200" swimtime="00:03:44.42" />
                    <SPLIT distance="300" swimtime="00:05:41.36" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada.  (Horário: 19:21)" eventid="1142" status="DSQ" swimtime="00:00:55.63" resultid="1411" heatid="2432" lane="8" entrytime="00:00:57.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Rampazzo" birthdate="2013-02-18" gender="M" nation="BRA" license="400269" swrid="5748679" athleteid="1830" externalid="400269">
              <RESULTS>
                <RESULT eventid="1089" points="232" swimtime="00:01:16.16" resultid="1831" heatid="2359" lane="5" />
                <RESULT eventid="1073" points="221" swimtime="00:03:08.54" resultid="1832" heatid="2340" lane="3" entrytime="00:03:11.32" entrycourse="LCM" />
                <RESULT eventid="1117" points="232" swimtime="00:05:57.90" resultid="1833" heatid="2395" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.24" />
                    <SPLIT distance="200" swimtime="00:02:52.99" />
                    <SPLIT distance="300" swimtime="00:04:27.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="217" swimtime="00:00:43.13" resultid="1834" heatid="2435" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Saber" birthdate="2014-06-04" gender="F" nation="BRA" license="392141" swrid="5602554" athleteid="1619" externalid="392141">
              <RESULTS>
                <RESULT eventid="1080" points="195" swimtime="00:00:50.23" resultid="1620" heatid="2348" lane="5" entrytime="00:00:49.34" entrycourse="LCM" />
                <RESULT eventid="1064" points="168" swimtime="00:03:24.12" resultid="1621" heatid="2329" lane="7" entrytime="00:03:55.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="160" swimtime="00:00:49.39" resultid="1622" heatid="2404" lane="5" entrytime="00:00:48.94" entrycourse="LCM" />
                <RESULT eventid="1108" points="164" swimtime="00:03:50.09" resultid="1623" heatid="2385" lane="7" entrytime="00:03:53.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:54.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Alice Silva Gomes Xavier" birthdate="2013-02-25" gender="F" nation="BRA" license="371040" swrid="5717241" athleteid="1758" externalid="371040">
              <RESULTS>
                <RESULT eventid="1098" points="260" swimtime="00:00:38.24" resultid="1759" heatid="2374" lane="7" entrytime="00:00:40.07" entrycourse="LCM" />
                <RESULT eventid="1086" points="344" swimtime="00:01:13.76" resultid="1760" heatid="2358" lane="3" entrytime="00:01:12.56" entrycourse="LCM" />
                <RESULT eventid="1114" points="332" swimtime="00:05:39.60" resultid="1761" heatid="2391" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.47" />
                    <SPLIT distance="200" swimtime="00:02:45.59" />
                    <SPLIT distance="300" swimtime="00:04:13.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="300" swimtime="00:00:43.52" resultid="1762" heatid="2433" lane="6" entrytime="00:00:43.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Bittencourt Ribas" birthdate="2013-02-01" gender="F" nation="BRA" license="372682" swrid="5588555" athleteid="1373" externalid="372682">
              <RESULTS>
                <RESULT eventid="1098" points="251" swimtime="00:00:38.71" resultid="1374" heatid="2374" lane="2" entrytime="00:00:39.54" entrycourse="LCM" />
                <RESULT eventid="1070" points="292" swimtime="00:03:09.99" resultid="1375" heatid="2337" lane="4" entrytime="00:03:06.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="263" swimtime="00:01:29.44" resultid="1376" heatid="2415" lane="1" entrytime="00:01:25.97" entrycourse="LCM" />
                <RESULT eventid="1114" points="261" swimtime="00:06:08.05" resultid="1377" heatid="2391" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.15" />
                    <SPLIT distance="200" swimtime="00:03:03.31" />
                    <SPLIT distance="300" swimtime="00:04:38.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Antunes Luzzi" birthdate="2014-02-14" gender="M" nation="BRA" license="391019" swrid="5602510" athleteid="1569" externalid="391019">
              <RESULTS>
                <RESULT eventid="1083" points="74" swimtime="00:01:01.81" resultid="1570" heatid="2350" lane="3" entrytime="00:01:00.39" entrycourse="LCM" />
                <RESULT eventid="1067" status="DNS" swimtime="00:00:00.00" resultid="1571" heatid="2332" lane="7" />
                <RESULT eventid="1127" points="59" swimtime="00:01:00.28" resultid="1572" heatid="2408" lane="2" entrytime="00:00:58.95" entrycourse="LCM" />
                <RESULT eventid="1139" points="91" swimtime="00:00:46.37" resultid="1573" heatid="2426" lane="5" entrytime="00:00:48.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Simioni Albuquerque" birthdate="2014-12-23" gender="F" nation="BRA" license="401980" swrid="5661355" athleteid="1708" externalid="401980">
              <RESULTS>
                <RESULT eventid="1092" points="218" swimtime="00:00:40.58" resultid="1709" heatid="2367" lane="3" entrytime="00:00:42.95" entrycourse="LCM" />
                <RESULT eventid="1064" points="173" swimtime="00:03:22.14" resultid="1710" heatid="2327" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="288" swimtime="00:00:35.74" resultid="1711" heatid="2424" lane="2" entrytime="00:00:38.39" entrycourse="LCM" />
                <RESULT eventid="1108" points="192" swimtime="00:03:38.60" resultid="1712" heatid="2383" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Artigas Pinheiro" birthdate="2013-07-31" gender="F" nation="BRA" license="377153" swrid="5588534" athleteid="1509" externalid="377153">
              <RESULTS>
                <RESULT eventid="1098" points="127" swimtime="00:00:48.53" resultid="1510" heatid="2372" lane="4" entrytime="00:00:50.21" entrycourse="LCM" />
                <RESULT eventid="1086" points="240" swimtime="00:01:23.18" resultid="1511" heatid="2356" lane="4" entrytime="00:01:23.99" entrycourse="LCM" />
                <RESULT eventid="1130" points="198" swimtime="00:01:38.29" resultid="1512" heatid="2414" lane="2" entrytime="00:01:34.78" entrycourse="LCM" />
                <RESULT eventid="1114" points="229" swimtime="00:06:24.34" resultid="1513" heatid="2391" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.46" />
                    <SPLIT distance="200" swimtime="00:03:09.90" />
                    <SPLIT distance="300" swimtime="00:04:50.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Vian" birthdate="2014-03-25" gender="F" nation="BRA" license="393919" swrid="5641779" athleteid="1663" externalid="393919">
              <RESULTS>
                <RESULT eventid="1092" points="134" swimtime="00:00:47.69" resultid="1664" heatid="2366" lane="4" entrytime="00:00:48.00" entrycourse="LCM" />
                <RESULT eventid="1064" points="170" swimtime="00:03:23.44" resultid="1665" heatid="2328" lane="8" />
                <RESULT eventid="1124" points="171" swimtime="00:00:48.36" resultid="1666" heatid="2405" lane="6" entrytime="00:00:45.73" entrycourse="LCM" />
                <RESULT eventid="1108" points="148" swimtime="00:03:58.02" resultid="1667" heatid="2382" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Clara Prado Biscaia" birthdate="2013-10-24" gender="F" nation="BRA" license="391015" swrid="5602526" athleteid="1554" externalid="391015">
              <RESULTS>
                <RESULT eventid="1098" points="172" swimtime="00:00:43.90" resultid="1555" heatid="2373" lane="3" entrytime="00:00:43.95" entrycourse="LCM" />
                <RESULT comment="SW 6.5 - Não terminou a prova enquanto estava de costas.&#10;&#10;&#10;&#10;&#10;&#10;&#10;  (Horário: 10:13), Na volta dos 100m (Medley Individual, Costas)." eventid="1070" status="DSQ" swimtime="00:03:31.45" resultid="1556" heatid="2336" lane="7" entrytime="00:03:40.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 6.4 - A virada não foi iniciada após a conclusão do movimento de braço, após sair da posição de costas.  (Horário: 18:20), Na volta dos 50m." eventid="1130" status="DSQ" swimtime="00:01:46.96" resultid="1557" heatid="2413" lane="5" />
                <RESULT eventid="1114" points="215" swimtime="00:06:32.38" resultid="1558" heatid="2392" lane="7" entrytime="00:06:55.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.64" />
                    <SPLIT distance="200" swimtime="00:03:12.55" />
                    <SPLIT distance="300" swimtime="00:04:55.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Fonseca Ribeiro" birthdate="2016-02-25" gender="F" nation="BRA" license="412016" swrid="5740011" athleteid="1820" externalid="412016">
              <RESULTS>
                <RESULT eventid="1060" status="DNS" swimtime="00:00:00.00" resultid="1821" heatid="2326" lane="3" />
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="1822" heatid="2343" lane="2" entrytime="00:01:06.47" entrycourse="LCM" />
                <RESULT eventid="1120" status="DNS" swimtime="00:00:00.00" resultid="1823" heatid="2399" lane="3" entrytime="00:00:53.85" entrycourse="LCM" />
                <RESULT eventid="1104" status="DNS" swimtime="00:00:00.00" resultid="1824" heatid="2380" lane="2" entrytime="00:01:08.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Gonçalves Sperandio" birthdate="2013-05-22" gender="M" nation="BRA" license="376980" swrid="5588851" athleteid="1435" externalid="376980">
              <RESULTS>
                <RESULT eventid="1101" points="153" swimtime="00:00:41.58" resultid="1436" heatid="2375" lane="3" />
                <RESULT eventid="1073" points="243" swimtime="00:03:02.64" resultid="1437" heatid="2341" lane="7" entrytime="00:03:08.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="278" swimtime="00:05:37.02" resultid="1438" heatid="2397" lane="8" entrytime="00:05:49.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.58" />
                    <SPLIT distance="200" swimtime="00:02:46.75" />
                    <SPLIT distance="300" swimtime="00:04:14.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="182" swimtime="00:00:45.76" resultid="1439" heatid="2437" lane="3" entrytime="00:00:49.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Betina" lastname="Vieira Pellanda" birthdate="2014-02-16" gender="F" nation="BRA" license="391041" swrid="5602589" athleteid="1609" externalid="391041">
              <RESULTS>
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="1610" heatid="2347" lane="5" entrytime="00:00:57.62" entrycourse="LCM" />
                <RESULT eventid="1064" status="DNS" swimtime="00:00:00.00" resultid="1611" heatid="2330" lane="3" entrytime="00:03:19.95" entrycourse="LCM" />
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="1612" heatid="2405" lane="1" entrytime="00:00:47.06" entrycourse="LCM" />
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="1613" heatid="2385" lane="6" entrytime="00:03:51.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Spadari Soso" birthdate="2012-12-28" gender="F" nation="BRA" license="377313" swrid="5588921" athleteid="1748" externalid="377313">
              <RESULTS>
                <RESULT eventid="1086" points="414" swimtime="00:01:09.37" resultid="1749" heatid="2357" lane="6" entrytime="00:01:20.12" entrycourse="LCM" />
                <RESULT eventid="1070" points="346" swimtime="00:02:59.58" resultid="1750" heatid="2335" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="412" swimtime="00:05:16.11" resultid="1751" heatid="2391" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.24" />
                    <SPLIT distance="200" swimtime="00:02:40.82" />
                    <SPLIT distance="300" swimtime="00:04:01.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="294" swimtime="00:00:43.82" resultid="1752" heatid="2433" lane="7" entrytime="00:00:44.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Wolf Macedo" birthdate="2012-01-27" gender="F" nation="BRA" license="369277" swrid="5602592" athleteid="1343" externalid="369277">
              <RESULTS>
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="1344" heatid="2374" lane="4" entrytime="00:00:33.76" entrycourse="LCM" />
                <RESULT eventid="1070" points="332" swimtime="00:03:02.10" resultid="1345" heatid="2338" lane="5" entrytime="00:02:56.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" status="DNS" swimtime="00:00:00.00" resultid="1346" heatid="2393" lane="7" entrytime="00:05:29.09" entrycourse="LCM" />
                <RESULT eventid="1142" status="DNS" swimtime="00:00:00.00" resultid="1347" heatid="2433" lane="3" entrytime="00:00:43.41" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia" lastname="Ziliotto Mehl" birthdate="2015-10-09" gender="F" nation="BRA" license="400122" swrid="5652905" athleteid="1703" externalid="400122">
              <RESULTS>
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="1704" heatid="2347" lane="3" entrytime="00:00:58.04" entrycourse="LCM" />
                <RESULT eventid="1064" status="DNS" swimtime="00:00:00.00" resultid="1705" heatid="2329" lane="6" entrytime="00:03:48.96" entrycourse="LCM" />
                <RESULT eventid="1136" status="DNS" swimtime="00:00:00.00" resultid="1706" heatid="2423" lane="3" entrytime="00:00:40.85" entrycourse="LCM" />
                <RESULT eventid="1108" status="DNS" swimtime="00:00:00.00" resultid="1707" heatid="2384" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Carcereri Navarro" birthdate="2013-12-19" gender="M" nation="BRA" license="376962" swrid="5588576" athleteid="1398" externalid="376962">
              <RESULTS>
                <RESULT eventid="1101" points="182" swimtime="00:00:39.28" resultid="1399" heatid="2377" lane="3" entrytime="00:00:40.67" entrycourse="LCM" />
                <RESULT eventid="1073" points="171" swimtime="00:03:25.35" resultid="1400" heatid="2339" lane="4" entrytime="00:03:25.77" entrycourse="LCM" />
                <RESULT eventid="1117" points="171" swimtime="00:06:36.34" resultid="1401" heatid="2395" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.16" />
                    <SPLIT distance="200" swimtime="00:03:14.96" />
                    <SPLIT distance="300" swimtime="00:04:56.97" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.4 - Movimentos das pernas não simultâneos.  (Horário: 19:26)" eventid="1145" status="DSQ" swimtime="00:00:44.23" resultid="1402" heatid="2438" lane="7" entrytime="00:00:45.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Calvo Ribas" birthdate="2016-01-09" gender="M" nation="BRA" license="415014" swrid="5755331" athleteid="1856" externalid="415014">
              <RESULTS>
                <RESULT eventid="1078" points="67" swimtime="00:00:57.81" resultid="1857" heatid="2344" lane="4" entrytime="00:00:55.21" entrycourse="LCM" />
                <RESULT eventid="1122" points="35" swimtime="00:01:03.34" resultid="1858" heatid="2401" lane="6" entrytime="00:01:05.06" entrycourse="LCM" />
                <RESULT eventid="1106" status="DNS" swimtime="00:00:00.00" resultid="1859" heatid="2381" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Corte Flor" birthdate="2016-12-03" gender="M" nation="BRA" license="412013" swrid="5740007" athleteid="1809" externalid="412013">
              <RESULTS>
                <RESULT eventid="1078" status="DNS" swimtime="00:00:00.00" resultid="1810" heatid="2344" lane="2" entrytime="00:01:09.91" entrycourse="LCM" />
                <RESULT eventid="1122" points="54" swimtime="00:00:55.25" resultid="1811" heatid="2400" lane="3" />
                <RESULT eventid="1106" points="52" swimtime="00:01:09.40" resultid="1812" heatid="2381" lane="5" entrytime="00:01:10.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Poletto Abrahao" birthdate="2014-10-20" gender="M" nation="BRA" license="382128" swrid="5602571" athleteid="1534" externalid="382128">
              <RESULTS>
                <RESULT eventid="1083" points="192" swimtime="00:00:44.97" resultid="1535" heatid="2352" lane="4" entrytime="00:00:44.75" entrycourse="LCM" />
                <RESULT eventid="1067" points="196" swimtime="00:02:55.44" resultid="1536" heatid="2334" lane="7" entrytime="00:03:05.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="150" swimtime="00:00:44.27" resultid="1537" heatid="2410" lane="2" entrytime="00:00:44.51" entrycourse="LCM" />
                <RESULT eventid="1111" points="220" swimtime="00:03:08.70" resultid="1538" heatid="2389" lane="4" entrytime="00:03:23.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Prosdocimo" birthdate="2012-11-30" gender="M" nation="BRA" license="369272" swrid="5602575" athleteid="1328" externalid="369272">
              <RESULTS>
                <RESULT eventid="1101" points="190" swimtime="00:00:38.68" resultid="1329" heatid="2375" lane="6" />
                <RESULT eventid="1089" points="324" swimtime="00:01:08.19" resultid="1330" heatid="2363" lane="5" entrytime="00:01:15.98" entrycourse="LCM" />
                <RESULT eventid="1133" points="232" swimtime="00:01:23.86" resultid="1331" heatid="2420" lane="1" entrytime="00:01:27.62" entrycourse="LCM" />
                <RESULT eventid="1117" points="324" swimtime="00:05:20.38" resultid="1332" heatid="2397" lane="4" entrytime="00:05:28.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.89" />
                    <SPLIT distance="200" swimtime="00:02:39.18" />
                    <SPLIT distance="300" swimtime="00:04:02.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="De Almeida Dias" birthdate="2012-02-18" gender="F" nation="BRA" license="369262" swrid="5588638" athleteid="1298" externalid="369262">
              <RESULTS>
                <RESULT eventid="1098" points="294" swimtime="00:00:36.74" resultid="1299" heatid="2371" lane="5" />
                <RESULT eventid="1086" points="452" swimtime="00:01:07.37" resultid="1300" heatid="2358" lane="4" entrytime="00:01:07.35" entrycourse="LCM" />
                <RESULT eventid="1130" points="351" swimtime="00:01:21.24" resultid="1301" heatid="2415" lane="6" entrytime="00:01:21.59" entrycourse="LCM" />
                <RESULT eventid="1114" points="434" swimtime="00:05:10.71" resultid="1302" heatid="2393" lane="6" entrytime="00:05:14.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.91" />
                    <SPLIT distance="200" swimtime="00:02:32.34" />
                    <SPLIT distance="300" swimtime="00:03:52.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Lauand Lorenci" birthdate="2013-03-06" gender="M" nation="BRA" license="376982" swrid="5588764" athleteid="1445" externalid="376982">
              <RESULTS>
                <RESULT eventid="1101" points="155" swimtime="00:00:41.38" resultid="1446" heatid="2377" lane="5" entrytime="00:00:39.74" entrycourse="LCM" />
                <RESULT eventid="1073" points="224" swimtime="00:03:07.51" resultid="1447" heatid="2340" lane="5" entrytime="00:03:10.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="236" swimtime="00:05:55.86" resultid="1448" heatid="2394" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.35" />
                    <SPLIT distance="200" swimtime="00:02:57.31" />
                    <SPLIT distance="300" swimtime="00:04:28.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="201" swimtime="00:00:44.28" resultid="1449" heatid="2438" lane="2" entrytime="00:00:43.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Lazzarotti Matias" birthdate="2012-03-19" gender="F" nation="BRA" license="391026" swrid="5602552" athleteid="1599" externalid="391026">
              <RESULTS>
                <RESULT eventid="1086" points="379" swimtime="00:01:11.44" resultid="1600" heatid="2354" lane="4" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 10:21), Na volta dos 150m (Medley Individual, Peito)." eventid="1070" status="DSQ" swimtime="00:03:02.35" resultid="1601" heatid="2338" lane="8" entrytime="00:03:04.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="386" swimtime="00:01:18.73" resultid="1602" heatid="2415" lane="3" entrytime="00:01:19.89" entrycourse="LCM" />
                <RESULT eventid="1142" points="249" swimtime="00:00:46.29" resultid="1603" heatid="2432" lane="5" entrytime="00:00:47.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Liam" lastname="Batista Grise" birthdate="2014-03-27" gender="M" nation="BRA" license="391008" swrid="5602514" athleteid="1544" externalid="391008">
              <RESULTS>
                <RESULT eventid="1095" points="65" swimtime="00:00:55.26" resultid="1545" heatid="2368" lane="1" />
                <RESULT eventid="1083" points="96" swimtime="00:00:56.64" resultid="1546" heatid="2351" lane="7" entrytime="00:00:54.92" entrycourse="LCM" />
                <RESULT eventid="1127" points="92" swimtime="00:00:52.09" resultid="1547" heatid="2408" lane="5" entrytime="00:00:56.44" entrycourse="LCM" />
                <RESULT eventid="1139" points="124" swimtime="00:00:41.90" resultid="1548" heatid="2427" lane="7" entrytime="00:00:43.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Weber Boguszewski" birthdate="2016-10-07" gender="M" nation="BRA" license="415255" swrid="5755346" athleteid="1860" externalid="415255">
              <RESULTS>
                <RESULT eventid="1078" points="29" swimtime="00:01:16.28" resultid="1861" heatid="2344" lane="3" entrytime="00:01:03.08" entrycourse="LCM" />
                <RESULT eventid="1122" points="53" swimtime="00:00:55.40" resultid="1862" heatid="2401" lane="7" entrytime="00:01:10.83" entrycourse="LCM" />
                <RESULT eventid="1106" points="30" swimtime="00:01:22.96" resultid="1863" heatid="2381" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivia" lastname="Mayer Paludetto" birthdate="2016-04-01" gender="F" nation="BRA" license="412014" swrid="5740014" athleteid="1813" externalid="412014">
              <RESULTS>
                <RESULT eventid="1060" points="25" swimtime="00:01:22.83" resultid="1814" heatid="2326" lane="4" entrytime="00:01:15.73" entrycourse="LCM" />
                <RESULT eventid="1076" points="83" swimtime="00:01:01.42" resultid="1815" heatid="2343" lane="4" entrytime="00:00:56.13" entrycourse="LCM" />
                <RESULT eventid="1120" points="72" swimtime="00:00:56.69" resultid="1816" heatid="2399" lane="4" entrytime="00:00:50.17" entrycourse="LCM" />
                <RESULT eventid="1104" points="107" swimtime="00:01:01.35" resultid="1817" heatid="2380" lane="5" entrytime="00:01:02.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Karam Barbosa Lima" birthdate="2012-12-11" gender="F" nation="BRA" license="376956" swrid="5588758" athleteid="1383" externalid="376956">
              <RESULTS>
                <RESULT eventid="1086" points="356" swimtime="00:01:12.91" resultid="1384" heatid="2358" lane="7" entrytime="00:01:14.88" entrycourse="LCM" />
                <RESULT eventid="1070" points="319" swimtime="00:03:04.43" resultid="1385" heatid="2337" lane="2" entrytime="00:03:11.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="283" swimtime="00:01:27.29" resultid="1386" heatid="2415" lane="2" entrytime="00:01:25.05" entrycourse="LCM" />
                <RESULT eventid="1114" points="378" swimtime="00:05:25.28" resultid="1387" heatid="2392" lane="5" entrytime="00:05:46.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.43" />
                    <SPLIT distance="200" swimtime="00:02:40.95" />
                    <SPLIT distance="300" swimtime="00:04:05.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Fernandes Tramujas" birthdate="2015-01-15" gender="F" nation="BRA" license="406750" swrid="5717263" athleteid="1743" externalid="406750">
              <RESULTS>
                <RESULT eventid="1080" points="76" swimtime="00:01:08.82" resultid="1744" heatid="2346" lane="1" entrytime="00:01:10.52" entrycourse="LCM" />
                <RESULT eventid="1064" points="122" swimtime="00:03:47.12" resultid="1745" heatid="2329" lane="8" entrytime="00:04:11.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="117" swimtime="00:00:48.20" resultid="1746" heatid="2422" lane="8" entrytime="00:00:47.76" entrycourse="LCM" />
                <RESULT eventid="1108" points="88" swimtime="00:04:43.47" resultid="1747" heatid="2383" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:26.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Dolberth Alcantara" birthdate="2014-09-26" gender="F" nation="BRA" license="382124" swrid="5602532" athleteid="1519" externalid="382124">
              <RESULTS>
                <RESULT eventid="1092" points="140" swimtime="00:00:47.01" resultid="1520" heatid="2367" lane="1" entrytime="00:00:46.74" entrycourse="LCM" />
                <RESULT eventid="1064" points="172" swimtime="00:03:22.78" resultid="1521" heatid="2328" lane="3" entrytime="00:04:19.57" entrycourse="LCM" />
                <RESULT eventid="1124" points="159" swimtime="00:00:49.51" resultid="1522" heatid="2404" lane="4" entrytime="00:00:48.62" entrycourse="LCM" />
                <RESULT eventid="1108" points="185" swimtime="00:03:41.06" resultid="1523" heatid="2385" lane="8" entrytime="00:03:57.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Emilia Abrahao" birthdate="2016-06-14" gender="F" nation="BRA" license="412012" swrid="5740010" athleteid="1806" externalid="412012">
              <RESULTS>
                <RESULT eventid="1120" status="DNS" swimtime="00:00:00.00" resultid="1807" heatid="2399" lane="2" entrytime="00:01:01.96" entrycourse="LCM" />
                <RESULT eventid="1104" status="DNS" swimtime="00:00:00.00" resultid="1808" heatid="2380" lane="6" entrytime="00:01:07.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Massimo" lastname="Puppi Cardoso" birthdate="2015-03-30" gender="M" nation="BRA" license="406742" swrid="5717290" athleteid="1723" externalid="406742">
              <RESULTS>
                <RESULT eventid="1083" status="DNS" swimtime="00:00:00.00" resultid="1724" heatid="2350" lane="4" entrytime="00:00:57.41" entrycourse="LCM" />
                <RESULT eventid="1067" status="DNS" swimtime="00:00:00.00" resultid="1725" heatid="2332" lane="6" />
                <RESULT eventid="1111" status="DNS" swimtime="00:00:00.00" resultid="1726" heatid="2388" lane="8" entrytime="00:04:46.93" entrycourse="LCM" />
                <RESULT eventid="1139" status="DNS" swimtime="00:00:00.00" resultid="1727" heatid="2426" lane="3" entrytime="00:00:48.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ravi" lastname="Osternack Erbe" birthdate="2013-08-10" gender="M" nation="BRA" license="372681" swrid="5588841" athleteid="1368" externalid="372681">
              <RESULTS>
                <RESULT eventid="1101" points="215" swimtime="00:00:37.15" resultid="1369" heatid="2377" lane="6" entrytime="00:00:40.83" entrycourse="LCM" />
                <RESULT eventid="1089" points="251" swimtime="00:01:14.27" resultid="1370" heatid="2362" lane="4" entrytime="00:01:21.15" entrycourse="LCM" />
                <RESULT eventid="1133" points="186" swimtime="00:01:30.33" resultid="1371" heatid="2420" lane="7" entrytime="00:01:27.59" entrycourse="LCM" />
                <RESULT eventid="1117" points="244" swimtime="00:05:52.09" resultid="1372" heatid="2394" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.14" />
                    <SPLIT distance="200" swimtime="00:02:55.97" />
                    <SPLIT distance="300" swimtime="00:04:27.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Trevisan De Paula" birthdate="2014-01-27" gender="M" nation="BRA" license="377152" swrid="5602568" athleteid="1504" externalid="377152">
              <RESULTS>
                <RESULT eventid="1095" points="192" swimtime="00:00:38.57" resultid="1505" heatid="2370" lane="4" entrytime="00:00:37.55" entrycourse="LCM" />
                <RESULT eventid="1067" points="220" swimtime="00:02:48.94" resultid="1506" heatid="2334" lane="4" entrytime="00:02:53.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="194" swimtime="00:03:16.59" resultid="1507" heatid="2389" lane="5" entrytime="00:03:25.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="223" swimtime="00:00:34.46" resultid="1508" heatid="2429" lane="4" entrytime="00:00:33.59" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13068" nation="BRA" region="PR" clubid="1934" swrid="93787" name="Sociedade Morgenau" shortname="Morgenau">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Cecilia Carstens" birthdate="2014-02-22" gender="F" nation="BRA" license="406721" swrid="5717251" athleteid="1970" externalid="406721">
              <RESULTS>
                <RESULT eventid="1136" points="188" swimtime="00:00:41.20" resultid="1971" heatid="2422" lane="5" entrytime="00:00:42.96" entrycourse="LCM" />
                <RESULT eventid="1108" points="159" swimtime="00:03:52.79" resultid="1972" heatid="2383" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:51.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Lara" birthdate="2014-09-02" gender="F" nation="BRA" license="406686" swrid="5717259" athleteid="1957" externalid="406686">
              <RESULTS>
                <RESULT eventid="1092" points="98" swimtime="00:00:52.89" resultid="1958" heatid="2366" lane="8" entrytime="00:00:53.72" entrycourse="LCM" />
                <RESULT eventid="1080" points="121" swimtime="00:00:58.81" resultid="1959" heatid="2346" lane="3" entrytime="00:01:03.13" entrycourse="LCM" />
                <RESULT eventid="1136" points="207" swimtime="00:00:39.86" resultid="1960" heatid="2423" lane="4" entrytime="00:00:40.41" entrycourse="LCM" />
                <RESULT eventid="1108" points="151" swimtime="00:03:56.47" resultid="1961" heatid="2384" lane="5" entrytime="00:04:34.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:52.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Seiffert Mafra" birthdate="2013-01-11" gender="F" nation="BRA" license="406729" swrid="5717296" athleteid="1978" externalid="406729">
              <RESULTS>
                <RESULT eventid="1098" points="87" swimtime="00:00:55.13" resultid="1979" heatid="2371" lane="3" />
                <RESULT eventid="1086" points="140" swimtime="00:01:39.58" resultid="1980" heatid="2355" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Fernanda De Lima" birthdate="2013-09-26" gender="F" nation="BRA" license="378290" swrid="5588693" athleteid="1940" externalid="378290">
              <RESULTS>
                <RESULT eventid="1098" points="113" swimtime="00:00:50.53" resultid="1941" heatid="2371" lane="4" />
                <RESULT eventid="1086" points="220" swimtime="00:01:25.65" resultid="1942" heatid="2356" lane="8" entrytime="00:01:33.38" entrycourse="LCM" />
                <RESULT eventid="1142" points="137" swimtime="00:00:56.45" resultid="1943" heatid="2431" lane="3" entrytime="00:01:01.33" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Paes Pereira" birthdate="2013-03-11" gender="M" nation="BRA" license="391137" swrid="5602567" athleteid="1944" externalid="391137">
              <RESULTS>
                <RESULT eventid="1101" points="102" swimtime="00:00:47.54" resultid="1945" heatid="2376" lane="6" entrytime="00:01:05.21" entrycourse="LCM" />
                <RESULT eventid="1089" points="141" swimtime="00:01:30.00" resultid="1946" heatid="2360" lane="3" entrytime="00:01:44.10" entrycourse="LCM" />
                <RESULT eventid="1133" points="109" swimtime="00:01:47.80" resultid="1947" heatid="2417" lane="1" />
                <RESULT eventid="1117" points="140" swimtime="00:07:03.56" resultid="1948" heatid="2394" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.86" />
                    <SPLIT distance="200" swimtime="00:03:25.98" />
                    <SPLIT distance="300" swimtime="00:05:17.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Gavinski Alves" birthdate="2012-10-12" gender="M" nation="BRA" license="369324" swrid="5588674" athleteid="1935" externalid="369324">
              <RESULTS>
                <RESULT eventid="1089" points="279" swimtime="00:01:11.69" resultid="1936" heatid="2363" lane="2" entrytime="00:01:18.86" entrycourse="LCM" />
                <RESULT eventid="1073" points="254" swimtime="00:02:59.98" resultid="1937" heatid="2341" lane="2" entrytime="00:03:05.09" entrycourse="LCM" />
                <RESULT eventid="1133" points="314" swimtime="00:01:15.85" resultid="1938" heatid="2420" lane="5" entrytime="00:01:19.94" entrycourse="LCM" />
                <RESULT eventid="1145" points="148" swimtime="00:00:48.99" resultid="1939" heatid="2434" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Tomaz Zmievski" birthdate="2012-09-20" gender="F" nation="BRA" license="406725" swrid="5717300" athleteid="1973" externalid="406725">
              <RESULTS>
                <RESULT eventid="1086" points="249" swimtime="00:01:22.16" resultid="1974" heatid="2356" lane="3" entrytime="00:01:26.76" entrycourse="LCM" />
                <RESULT eventid="1070" points="217" swimtime="00:03:29.75" resultid="1975" heatid="2336" lane="3" entrytime="00:03:35.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="214" swimtime="00:01:35.84" resultid="1976" heatid="2413" lane="1" />
                <RESULT eventid="1142" points="163" swimtime="00:00:53.35" resultid="1977" heatid="2431" lane="4" entrytime="00:00:57.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Melo" birthdate="2015-02-07" gender="F" nation="BRA" license="406717" swrid="5717280" athleteid="1962" externalid="406717">
              <RESULTS>
                <RESULT eventid="1092" points="103" swimtime="00:00:52.09" resultid="1963" heatid="2366" lane="3" entrytime="00:00:50.43" entrycourse="LCM" />
                <RESULT eventid="1080" points="93" swimtime="00:01:04.34" resultid="1964" heatid="2345" lane="3" />
                <RESULT eventid="1124" points="192" swimtime="00:00:46.48" resultid="1965" heatid="2405" lane="5" entrytime="00:00:43.99" entrycourse="LCM" />
                <RESULT eventid="1108" points="148" swimtime="00:03:58.05" resultid="1966" heatid="2383" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maryana" lastname="Lemos Carvalho" birthdate="2014-02-10" gender="F" nation="BRA" license="406718" swrid="5717278" athleteid="1967" externalid="406718">
              <RESULTS>
                <RESULT eventid="1064" points="127" swimtime="00:03:44.14" resultid="1968" heatid="2329" lane="1" entrytime="00:04:10.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="138" swimtime="00:00:51.93" resultid="1969" heatid="2403" lane="4" entrytime="00:00:56.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Nitz Costa" birthdate="2015-02-09" gender="F" nation="BRA" license="397328" swrid="5641773" athleteid="1952" externalid="397328">
              <RESULTS>
                <RESULT eventid="1092" points="159" swimtime="00:00:45.08" resultid="1953" heatid="2367" lane="2" entrytime="00:00:43.07" entrycourse="LCM" />
                <RESULT eventid="1064" points="239" swimtime="00:03:01.67" resultid="1954" heatid="2330" lane="6" entrytime="00:03:20.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="251" swimtime="00:00:37.42" resultid="1955" heatid="2424" lane="6" entrytime="00:00:37.75" entrycourse="LCM" />
                <RESULT eventid="1108" points="201" swimtime="00:03:35.30" resultid="1956" heatid="2383" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Felipe Kuhn" birthdate="2014-03-22" gender="M" nation="BRA" license="392121" swrid="5602536" athleteid="1949" externalid="392121">
              <RESULTS>
                <RESULT eventid="1095" points="112" swimtime="00:00:46.11" resultid="1950" heatid="2368" lane="2" />
                <RESULT eventid="1083" points="142" swimtime="00:00:49.69" resultid="1951" heatid="2352" lane="6" entrytime="00:00:50.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11303" nation="BRA" region="PR" clubid="1242" swrid="93760" name="Associação De Talentos Da Natação" shortname="Atn/Curitiba">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Eduarda Guedes Braga" birthdate="2013-04-09" gender="F" nation="BRA" license="385009" swrid="5602534" athleteid="1243" externalid="385009">
              <RESULTS>
                <RESULT eventid="1098" points="160" swimtime="00:00:45.00" resultid="1244" heatid="2372" lane="5" entrytime="00:00:50.46" entrycourse="LCM" />
                <RESULT eventid="1086" points="286" swimtime="00:01:18.46" resultid="1245" heatid="2358" lane="1" entrytime="00:01:14.94" entrycourse="LCM" />
                <RESULT eventid="1130" points="238" swimtime="00:01:32.40" resultid="1246" heatid="2414" lane="6" entrytime="00:01:33.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maximilian" lastname="Hock" birthdate="2016-11-20" gender="M" nation="DEU" license="408352" athleteid="1270" externalid="408352">
              <RESULTS>
                <RESULT eventid="1078" points="70" swimtime="00:00:57.00" resultid="1271" heatid="2344" lane="5" entrytime="00:01:00.03" entrycourse="LCM" />
                <RESULT eventid="1122" points="91" swimtime="00:00:46.44" resultid="1272" heatid="2401" lane="4" entrytime="00:00:47.58" entrycourse="LCM" />
                <RESULT eventid="1106" points="69" swimtime="00:01:03.07" resultid="1273" heatid="2381" lane="4" entrytime="00:01:02.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Manuela Souza" birthdate="2016-07-07" gender="F" nation="BRA" license="406759" swrid="5717282" athleteid="1261" externalid="406759">
              <RESULTS>
                <RESULT eventid="1076" points="85" swimtime="00:01:00.94" resultid="1262" heatid="2343" lane="3" entrytime="00:01:02.34" entrycourse="LCM" />
                <RESULT eventid="1120" points="98" swimtime="00:00:51.10" resultid="1263" heatid="2399" lane="6" entrytime="00:00:53.99" entrycourse="LCM" />
                <RESULT eventid="1104" points="129" swimtime="00:00:57.69" resultid="1264" heatid="2380" lane="4" entrytime="00:00:58.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Lemes Luis" birthdate="2013-10-14" gender="M" nation="BRA" license="410105" swrid="5740012" athleteid="1274" externalid="410105">
              <RESULTS>
                <RESULT eventid="1101" points="64" swimtime="00:00:55.51" resultid="1275" heatid="2375" lane="5" />
                <RESULT eventid="1089" points="121" swimtime="00:01:34.60" resultid="1276" heatid="2361" lane="8" entrytime="00:01:31.33" entrycourse="LCM" />
                <RESULT eventid="1133" points="129" swimtime="00:01:41.86" resultid="1277" heatid="2418" lane="5" />
                <RESULT eventid="1145" points="130" swimtime="00:00:51.12" resultid="1278" heatid="2435" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Goncalves Ghion" birthdate="2014-10-15" gender="F" nation="BRA" license="406912" swrid="5717269" athleteid="1265" externalid="406912">
              <RESULTS>
                <RESULT eventid="1092" points="79" swimtime="00:00:56.90" resultid="1266" heatid="2365" lane="8" />
                <RESULT eventid="1080" points="123" swimtime="00:00:58.62" resultid="1267" heatid="2347" lane="2" entrytime="00:00:58.47" entrycourse="LCM" />
                <RESULT eventid="1136" points="151" swimtime="00:00:44.24" resultid="1268" heatid="2423" lane="2" entrytime="00:00:41.59" entrycourse="LCM" />
                <RESULT eventid="1124" points="109" swimtime="00:00:56.12" resultid="1269" heatid="2403" lane="7" entrytime="00:00:57.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Duarte De Almeida" birthdate="2013-12-09" gender="M" nation="BRA" license="385711" swrid="5588666" athleteid="1250" externalid="385711">
              <RESULTS>
                <RESULT eventid="1089" points="277" swimtime="00:01:11.83" resultid="1251" heatid="2363" lane="7" entrytime="00:01:20.03" entrycourse="LCM" />
                <RESULT eventid="1073" points="219" swimtime="00:03:09.09" resultid="1252" heatid="2339" lane="5" entrytime="00:03:26.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="197" swimtime="00:00:44.59" resultid="1253" heatid="2437" lane="4" entrytime="00:00:45.96" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isis" lastname="De Miranda" birthdate="2012-01-10" gender="F" nation="BRA" license="397278" swrid="5652886" athleteid="1254" externalid="397278">
              <RESULTS>
                <RESULT eventid="1098" points="206" swimtime="00:00:41.31" resultid="1255" heatid="2373" lane="6" entrytime="00:00:44.36" entrycourse="LCM" />
                <RESULT eventid="1086" points="301" swimtime="00:01:17.11" resultid="1256" heatid="2357" lane="8" entrytime="00:01:21.23" entrycourse="LCM" />
                <RESULT eventid="1114" points="304" swimtime="00:05:49.86" resultid="1257" heatid="2392" lane="3" entrytime="00:06:03.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.55" />
                    <SPLIT distance="200" swimtime="00:02:50.90" />
                    <SPLIT distance="300" swimtime="00:04:20.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Leal Kuss" birthdate="2012-10-20" gender="M" nation="BRA" license="385085" swrid="5588768" athleteid="1247" externalid="385085">
              <RESULTS>
                <RESULT eventid="1101" points="210" swimtime="00:00:37.43" resultid="1248" heatid="2378" lane="6" entrytime="00:00:36.21" entrycourse="LCM" />
                <RESULT eventid="1089" points="244" swimtime="00:01:14.92" resultid="1249" heatid="2362" lane="1" entrytime="00:01:24.89" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isaac" lastname="Zonta" birthdate="2012-11-14" gender="M" nation="BRA" license="414857" swrid="5755348" athleteid="1279" externalid="414857">
              <RESULTS>
                <RESULT eventid="1089" points="199" swimtime="00:01:20.26" resultid="1280" heatid="2359" lane="6" />
                <RESULT eventid="1145" points="111" swimtime="00:00:53.95" resultid="1281" heatid="2435" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yohanna" lastname="Vitoria Sena" birthdate="2012-01-20" gender="F" nation="BRA" license="406710" swrid="5717302" athleteid="1258" externalid="406710">
              <RESULTS>
                <RESULT eventid="1086" points="200" swimtime="00:01:28.29" resultid="1259" heatid="2355" lane="3" entrytime="00:01:42.36" entrycourse="LCM" />
                <RESULT eventid="1130" points="121" swimtime="00:01:55.87" resultid="1260" heatid="2413" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2864" nation="BRA" region="PR" clubid="1148" swrid="93756" name="Associacao De Pais E Amigos Da Natacao De Ponta Gr" shortname="Apan Ponta Grossa">
          <ATHLETES>
            <ATHLETE firstname="Theo" lastname="Campagnoli" birthdate="2013-03-13" gender="M" nation="BRA" license="370651" swrid="5602519" athleteid="1151" externalid="370651">
              <RESULTS>
                <RESULT eventid="1101" points="246" swimtime="00:00:35.53" resultid="1152" heatid="2378" lane="3" entrytime="00:00:35.66" entrycourse="LCM" />
                <RESULT eventid="1089" points="281" swimtime="00:01:11.50" resultid="1153" heatid="2364" lane="6" entrytime="00:01:10.40" entrycourse="LCM" />
                <RESULT eventid="1133" points="261" swimtime="00:01:20.70" resultid="1154" heatid="2420" lane="3" entrytime="00:01:22.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Clara Domingues" birthdate="2012-01-19" gender="F" nation="BRA" license="377291" swrid="5588599" athleteid="1149" externalid="377291">
              <RESULTS>
                <RESULT eventid="1086" points="282" swimtime="00:01:18.79" resultid="1150" heatid="2356" lane="6" entrytime="00:01:27.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Clara Rigailo" birthdate="2013-04-06" gender="F" nation="BRA" license="396828" swrid="5641758" athleteid="1168" externalid="396828">
              <RESULTS>
                <RESULT eventid="1086" points="259" swimtime="00:01:21.08" resultid="1169" heatid="2354" lane="6" />
                <RESULT eventid="1142" points="300" swimtime="00:00:43.54" resultid="1170" heatid="2433" lane="2" entrytime="00:00:44.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Bischof Rogoski" birthdate="2014-10-03" gender="M" nation="BRA" license="401860" swrid="5661341" athleteid="1174" externalid="401860">
              <RESULTS>
                <RESULT eventid="1095" points="123" swimtime="00:00:44.70" resultid="1175" heatid="2370" lane="1" entrytime="00:00:42.79" entrycourse="LCM" />
                <RESULT eventid="1083" points="153" swimtime="00:00:48.45" resultid="1176" heatid="2352" lane="2" entrytime="00:00:50.23" entrycourse="LCM" />
                <RESULT eventid="1139" points="199" swimtime="00:00:35.76" resultid="1177" heatid="2429" lane="1" entrytime="00:00:36.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Victoria Borges" birthdate="2014-01-16" gender="F" nation="BRA" license="376737" swrid="5602587" athleteid="1155" externalid="376737">
              <RESULTS>
                <RESULT eventid="1092" points="99" swimtime="00:00:52.66" resultid="1156" heatid="2366" lane="7" entrytime="00:00:52.55" entrycourse="LCM" />
                <RESULT eventid="1064" points="179" swimtime="00:03:20.04" resultid="1157" heatid="2330" lane="1" entrytime="00:03:35.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="230" swimtime="00:00:38.53" resultid="1158" heatid="2424" lane="3" entrytime="00:00:37.71" entrycourse="LCM" />
                <RESULT eventid="1124" points="175" swimtime="00:00:47.95" resultid="1159" heatid="2405" lane="7" entrytime="00:00:46.32" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Hilgenberg Lievore" birthdate="2014-04-23" gender="M" nation="BRA" license="391167" swrid="5602546" athleteid="1165" externalid="391167">
              <RESULTS>
                <RESULT eventid="1127" points="167" swimtime="00:00:42.68" resultid="1166" heatid="2410" lane="6" entrytime="00:00:43.29" entrycourse="LCM" />
                <RESULT eventid="1139" points="166" swimtime="00:00:38.00" resultid="1167" heatid="2428" lane="4" entrytime="00:00:36.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Miretzki" birthdate="2014-09-17" gender="F" nation="BRA" license="414996" swrid="5755341" athleteid="1178" externalid="414996">
              <RESULTS>
                <RESULT eventid="1080" points="112" swimtime="00:01:00.32" resultid="1179" heatid="2347" lane="7" entrytime="00:00:59.88" entrycourse="LCM" />
                <RESULT eventid="1136" points="206" swimtime="00:00:39.96" resultid="1180" heatid="2421" lane="2" />
                <RESULT eventid="1124" points="144" swimtime="00:00:51.13" resultid="1181" heatid="2402" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emanuel" lastname="Lucas Ribeiro" birthdate="2014-03-28" gender="M" nation="BRA" license="414997" swrid="5755338" athleteid="1182" externalid="414997">
              <RESULTS>
                <RESULT eventid="1083" points="97" swimtime="00:00:56.34" resultid="1183" heatid="2351" lane="8" entrytime="00:00:56.03" entrycourse="LCM" />
                <RESULT eventid="1127" points="81" swimtime="00:00:54.42" resultid="1184" heatid="2409" lane="1" entrytime="00:00:55.42" entrycourse="LCM" />
                <RESULT eventid="1139" points="95" swimtime="00:00:45.74" resultid="1185" heatid="2427" lane="8" entrytime="00:00:45.56" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolly" lastname="Victoria Souza" birthdate="2015-11-15" gender="F" nation="BRA" license="400091" swrid="5652902" athleteid="1171" externalid="400091">
              <RESULTS>
                <RESULT eventid="1080" points="160" swimtime="00:00:53.65" resultid="1172" heatid="2348" lane="8" entrytime="00:00:54.46" entrycourse="LCM" />
                <RESULT eventid="1136" points="156" swimtime="00:00:43.78" resultid="1173" heatid="2423" lane="8" entrytime="00:00:42.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariana" lastname="Brunetti Silva" birthdate="2014-03-24" gender="F" nation="BRA" license="390878" swrid="5602517" athleteid="1160" externalid="390878">
              <RESULTS>
                <RESULT eventid="1092" points="66" swimtime="00:01:00.35" resultid="1161" heatid="2366" lane="1" entrytime="00:00:53.21" entrycourse="LCM" />
                <RESULT eventid="1080" points="152" swimtime="00:00:54.55" resultid="1162" heatid="2347" lane="4" entrytime="00:00:54.91" entrycourse="LCM" />
                <RESULT eventid="1136" points="215" swimtime="00:00:39.40" resultid="1163" heatid="2423" lane="5" entrytime="00:00:40.65" entrycourse="LCM" />
                <RESULT eventid="1124" points="147" swimtime="00:00:50.78" resultid="1164" heatid="2404" lane="3" entrytime="00:00:50.19" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1007" nation="BRA" region="PR" clubid="1981" swrid="93785" name="Santa Mônica Clube De Campo" shortname="Santa Mônica">
          <ATHLETES>
            <ATHLETE firstname="Pedro" lastname="Marini" birthdate="2014-04-09" gender="M" nation="BRA" license="382247" swrid="5684582" athleteid="2017" externalid="382247">
              <RESULTS>
                <RESULT eventid="1095" points="128" swimtime="00:00:44.12" resultid="2018" heatid="2370" lane="8" entrytime="00:00:43.78" entrycourse="LCM" />
                <RESULT eventid="1083" points="95" swimtime="00:00:56.74" resultid="2019" heatid="2350" lane="2" entrytime="00:01:01.99" entrycourse="LCM" />
                <RESULT eventid="1111" points="134" swimtime="00:03:42.55" resultid="2020" heatid="2386" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="144" swimtime="00:00:39.87" resultid="2021" heatid="2428" lane="8" entrytime="00:00:40.41" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Szpak Costa" birthdate="2015-05-19" gender="M" nation="BRA" license="416974" athleteid="2151" externalid="416974">
              <RESULTS>
                <RESULT eventid="1127" points="45" swimtime="00:01:05.88" resultid="2152" heatid="2406" lane="4" />
                <RESULT eventid="1139" points="54" swimtime="00:00:55.02" resultid="2153" heatid="2425" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Hugo Dos Santos" birthdate="2014-07-25" gender="M" nation="BRA" license="397420" swrid="5641766" athleteid="2085" externalid="397420">
              <RESULTS>
                <RESULT eventid="1095" points="55" swimtime="00:00:58.31" resultid="2086" heatid="2369" lane="7" entrytime="00:00:56.06" entrycourse="LCM" />
                <RESULT eventid="1083" points="91" swimtime="00:00:57.60" resultid="2087" heatid="2351" lane="1" entrytime="00:00:55.67" entrycourse="LCM" />
                <RESULT eventid="1111" points="99" swimtime="00:04:05.79" resultid="2088" heatid="2388" lane="5" entrytime="00:04:13.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:04.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="153" swimtime="00:00:39.06" resultid="2089" heatid="2427" lane="3" entrytime="00:00:40.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helloisa" lastname="De Bassani" birthdate="2012-09-23" gender="F" nation="BRA" license="403403" swrid="5676296" athleteid="2118" externalid="403403">
              <RESULTS>
                <RESULT eventid="1086" points="153" swimtime="00:01:36.60" resultid="2119" heatid="2355" lane="7" entrytime="00:02:17.31" entrycourse="LCM" />
                <RESULT comment="SW 6.4 - A virada não foi iniciada após a conclusão do movimento de braço, após sair da posição de costas.  (Horário: 18:16), Na volta dos 50 m " eventid="1130" status="DSQ" swimtime="00:01:56.89" resultid="2120" heatid="2412" lane="4" />
                <RESULT eventid="1142" points="105" swimtime="00:01:01.75" resultid="2121" heatid="2431" lane="5" entrytime="00:00:58.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Luiza Rocha Batista" birthdate="2013-11-24" gender="F" nation="BRA" license="387379" swrid="5588784" athleteid="2046" externalid="387379">
              <RESULTS>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 12:10)" eventid="1098" status="DSQ" swimtime="00:00:47.48" resultid="2047" heatid="2373" lane="1" entrytime="00:00:49.00" entrycourse="LCM" />
                <RESULT eventid="1086" points="267" swimtime="00:01:20.21" resultid="2048" heatid="2356" lane="5" entrytime="00:01:25.62" entrycourse="LCM" />
                <RESULT eventid="1130" points="204" swimtime="00:01:37.32" resultid="2049" heatid="2411" lane="5" />
                <RESULT eventid="1114" points="215" swimtime="00:06:32.60" resultid="2050" heatid="2391" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.28" />
                    <SPLIT distance="300" swimtime="00:04:56.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cleverson" lastname="Cardoso" birthdate="2013-07-20" gender="M" nation="BRA" license="387382" swrid="5588577" athleteid="2051" externalid="387382">
              <RESULTS>
                <RESULT eventid="1101" points="80" swimtime="00:00:51.52" resultid="2052" heatid="2376" lane="2" />
                <RESULT eventid="1089" points="194" swimtime="00:01:20.85" resultid="2053" heatid="2361" lane="5" entrytime="00:01:27.27" entrycourse="LCM" />
                <RESULT eventid="1133" points="143" swimtime="00:01:38.53" resultid="2054" heatid="2417" lane="6" />
                <RESULT eventid="1145" points="152" swimtime="00:00:48.62" resultid="2055" heatid="2437" lane="6" entrytime="00:00:50.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mathias" lastname="Bernardo" birthdate="2014-05-17" gender="M" nation="BRA" license="387376" swrid="5652880" athleteid="2036" externalid="387376">
              <RESULTS>
                <RESULT eventid="1095" points="65" swimtime="00:00:55.11" resultid="2037" heatid="2369" lane="6" entrytime="00:00:50.94" entrycourse="LCM" />
                <RESULT eventid="1083" points="102" swimtime="00:00:55.43" resultid="2038" heatid="2350" lane="6" entrytime="00:01:01.30" entrycourse="LCM" />
                <RESULT eventid="1127" points="112" swimtime="00:00:48.72" resultid="2039" heatid="2409" lane="7" entrytime="00:00:51.01" entrycourse="LCM" />
                <RESULT eventid="1111" points="146" swimtime="00:03:36.18" resultid="2040" heatid="2387" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="Cirilo Da Cunha" birthdate="2013-05-26" gender="F" nation="BRA" license="377316" swrid="5588595" athleteid="1997" externalid="377316">
              <RESULTS>
                <RESULT eventid="1086" points="274" swimtime="00:01:19.58" resultid="1998" heatid="2357" lane="2" entrytime="00:01:20.49" entrycourse="LCM" />
                <RESULT eventid="1070" points="271" swimtime="00:03:14.75" resultid="1999" heatid="2336" lane="4" entrytime="00:03:29.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="247" swimtime="00:01:31.31" resultid="2000" heatid="2412" lane="5" />
                <RESULT eventid="1114" points="275" swimtime="00:06:01.59" resultid="2001" heatid="2390" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.36" />
                    <SPLIT distance="200" swimtime="00:03:02.70" />
                    <SPLIT distance="300" swimtime="00:04:35.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Luiz Cruz" birthdate="2012-10-13" gender="M" nation="BRA" license="393209" swrid="5616447" athleteid="2066" externalid="393209">
              <RESULTS>
                <RESULT eventid="1101" points="185" swimtime="00:00:39.07" resultid="2067" heatid="2377" lane="2" entrytime="00:00:42.41" entrycourse="LCM" />
                <RESULT eventid="1073" points="175" swimtime="00:03:23.50" resultid="2068" heatid="2339" lane="6" entrytime="00:03:42.84" entrycourse="LCM" />
                <RESULT eventid="1117" points="221" swimtime="00:06:03.72" resultid="2069" heatid="2396" lane="2" entrytime="00:06:39.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.25" />
                    <SPLIT distance="200" swimtime="00:02:58.10" />
                    <SPLIT distance="300" swimtime="00:04:30.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="140" swimtime="00:00:49.91" resultid="2070" heatid="2437" lane="7" entrytime="00:00:51.13" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Strapasson" birthdate="2012-03-01" gender="M" nation="BRA" license="371377" swrid="5602585" athleteid="1982" externalid="371377">
              <RESULTS>
                <RESULT eventid="1101" points="209" swimtime="00:00:37.51" resultid="1983" heatid="2377" lane="7" entrytime="00:00:43.06" entrycourse="LCM" />
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 11:49)" eventid="1089" status="DSQ" swimtime="00:01:06.12" resultid="1984" heatid="2364" lane="5" entrytime="00:01:07.75" entrycourse="LCM" />
                <RESULT eventid="1117" points="292" swimtime="00:05:31.60" resultid="1985" heatid="2397" lane="7" entrytime="00:05:41.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.57" />
                    <SPLIT distance="200" swimtime="00:02:40.86" />
                    <SPLIT distance="300" swimtime="00:04:06.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="295" swimtime="00:00:38.95" resultid="1986" heatid="2438" lane="5" entrytime="00:00:40.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Prestes" birthdate="2014-01-16" gender="M" nation="BRA" license="382249" swrid="5602574" athleteid="2022" externalid="382249">
              <RESULTS>
                <RESULT eventid="1083" points="159" swimtime="00:00:47.83" resultid="2023" heatid="2352" lane="5" entrytime="00:00:47.63" entrycourse="LCM" />
                <RESULT eventid="1067" points="178" swimtime="00:03:01.23" resultid="2024" heatid="2334" lane="1" entrytime="00:03:14.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="140" swimtime="00:00:45.35" resultid="2025" heatid="2410" lane="7" entrytime="00:00:44.77" entrycourse="LCM" />
                <RESULT eventid="1139" points="205" swimtime="00:00:35.44" resultid="2026" heatid="2429" lane="7" entrytime="00:00:36.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Camily Moraes" birthdate="2014-07-13" gender="F" nation="BRA" license="397159" swrid="5641755" athleteid="2080" externalid="397159">
              <RESULTS>
                <RESULT eventid="1092" points="89" swimtime="00:00:54.52" resultid="2081" heatid="2365" lane="4" entrytime="00:00:54.48" entrycourse="LCM" />
                <RESULT eventid="1080" points="134" swimtime="00:00:56.92" resultid="2082" heatid="2345" lane="4" entrytime="00:01:33.18" entrycourse="LCM" />
                <RESULT eventid="1136" points="199" swimtime="00:00:40.38" resultid="2083" heatid="2424" lane="7" entrytime="00:00:38.59" entrycourse="LCM" />
                <RESULT eventid="1124" points="197" swimtime="00:00:46.16" resultid="2084" heatid="2405" lane="2" entrytime="00:00:46.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Zanotto Souza" birthdate="2015-07-01" gender="M" nation="BRA" license="415249" swrid="5755347" athleteid="2143" externalid="415249">
              <RESULTS>
                <RESULT eventid="1127" points="64" swimtime="00:00:58.66" resultid="2144" heatid="2407" lane="3" />
                <RESULT eventid="1139" points="98" swimtime="00:00:45.29" resultid="2145" heatid="2426" lane="4" entrytime="00:00:46.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lais" lastname="Manika Broto" birthdate="2013-03-27" gender="F" nation="BRA" license="378054" swrid="5588795" athleteid="2012" externalid="378054">
              <RESULTS>
                <RESULT eventid="1086" points="339" swimtime="00:01:14.15" resultid="2013" heatid="2358" lane="5" entrytime="00:01:11.50" entrycourse="LCM" />
                <RESULT eventid="1070" points="338" swimtime="00:03:00.90" resultid="2014" heatid="2338" lane="7" entrytime="00:03:04.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1114" points="379" swimtime="00:05:25.21" resultid="2015" heatid="2393" lane="1" entrytime="00:05:34.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.28" />
                    <SPLIT distance="200" swimtime="00:02:39.99" />
                    <SPLIT distance="300" swimtime="00:04:06.06" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.4 - A cabeça não rompeu a superfície durante cada ciclo do nado.  (Horário: 19:05)" eventid="1142" status="DSQ" swimtime="00:00:46.69" resultid="2016" heatid="2430" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Gabriel Broto" birthdate="2014-09-14" gender="M" nation="BRA" license="402171" swrid="5661345" athleteid="2109" externalid="402171">
              <RESULTS>
                <RESULT eventid="1083" points="32" swimtime="00:01:21.68" resultid="2110" heatid="2349" lane="6" />
                <RESULT eventid="1067" points="77" swimtime="00:03:59.74" resultid="2111" heatid="2331" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="54" swimtime="00:01:02.30" resultid="2112" heatid="2407" lane="5" entrytime="00:01:09.72" entrycourse="LCM" />
                <RESULT eventid="1139" points="69" swimtime="00:00:50.93" resultid="2113" heatid="2426" lane="8" entrytime="00:00:57.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Zattar" birthdate="2012-04-19" gender="F" nation="BRA" license="401736" swrid="5661351" athleteid="2104" externalid="401736">
              <RESULTS>
                <RESULT eventid="1098" points="330" swimtime="00:00:35.32" resultid="2105" heatid="2372" lane="1" />
                <RESULT eventid="1070" points="334" swimtime="00:03:01.70" resultid="2106" heatid="2337" lane="8" entrytime="00:03:18.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="244" swimtime="00:01:31.67" resultid="2107" heatid="2414" lane="3" entrytime="00:01:32.30" entrycourse="LCM" />
                <RESULT eventid="1142" points="328" swimtime="00:00:42.26" resultid="2108" heatid="2432" lane="4" entrytime="00:00:46.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Victoria De Medeiros" birthdate="2014-08-14" gender="F" nation="BRA" license="403782" swrid="5684611" athleteid="2122" externalid="403782">
              <RESULTS>
                <RESULT eventid="1092" points="76" swimtime="00:00:57.43" resultid="2123" heatid="2365" lane="5" entrytime="00:00:55.20" entrycourse="LCM" />
                <RESULT eventid="1080" points="141" swimtime="00:00:55.90" resultid="2124" heatid="2347" lane="6" entrytime="00:00:58.11" entrycourse="LCM" />
                <RESULT eventid="1136" points="167" swimtime="00:00:42.85" resultid="2125" heatid="2422" lane="2" entrytime="00:00:46.23" entrycourse="LCM" />
                <RESULT eventid="1124" points="113" swimtime="00:00:55.52" resultid="2126" heatid="2403" lane="3" entrytime="00:00:56.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="De Siqueira Machado" birthdate="2012-05-25" gender="F" nation="BRA" license="377312" swrid="5588649" athleteid="1987" externalid="377312">
              <RESULTS>
                <RESULT eventid="1086" points="340" swimtime="00:01:14.07" resultid="1988" heatid="2357" lane="3" entrytime="00:01:18.75" entrycourse="LCM" />
                <RESULT eventid="1070" points="249" swimtime="00:03:20.45" resultid="1989" heatid="2337" lane="7" entrytime="00:03:15.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="274" swimtime="00:01:28.23" resultid="1990" heatid="2414" lane="7" entrytime="00:01:35.94" entrycourse="LCM" />
                <RESULT eventid="1142" points="266" swimtime="00:00:45.33" resultid="1991" heatid="2433" lane="1" entrytime="00:00:44.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Monteiro Reboucas" birthdate="2015-02-23" gender="M" nation="BRA" license="416975" athleteid="2154" externalid="416975">
              <RESULTS>
                <RESULT eventid="1127" points="60" swimtime="00:00:59.90" resultid="2155" heatid="2407" lane="7" />
                <RESULT eventid="1139" points="29" swimtime="00:01:07.35" resultid="2156" heatid="2425" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helenna" lastname="Banzatto Silva" birthdate="2013-07-11" gender="F" nation="BRA" license="393210" swrid="5616439" athleteid="2071" externalid="393210">
              <RESULTS>
                <RESULT eventid="1086" points="86" swimtime="00:01:56.78" resultid="2072" heatid="2355" lane="1" entrytime="00:02:40.28" entrycourse="LCM" />
                <RESULT eventid="1130" points="77" swimtime="00:02:14.39" resultid="2073" heatid="2413" lane="3" />
                <RESULT eventid="1142" points="144" swimtime="00:00:55.51" resultid="2074" heatid="2432" lane="1" entrytime="00:00:55.62" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Borges Piekarzievicz" birthdate="2013-09-10" gender="M" nation="BRA" license="403142" swrid="5676294" athleteid="2114" externalid="403142">
              <RESULTS>
                <RESULT eventid="1101" points="61" swimtime="00:00:56.29" resultid="2115" heatid="2376" lane="8" />
                <RESULT eventid="1089" points="129" swimtime="00:01:32.62" resultid="2116" heatid="2360" lane="4" entrytime="00:01:35.74" entrycourse="LCM" />
                <RESULT eventid="1145" points="105" swimtime="00:00:55.00" resultid="2117" heatid="2436" lane="5" entrytime="00:00:53.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Rodrigues Bortoluzzi" birthdate="2013-10-07" gender="M" nation="BRA" license="387375" swrid="5652897" athleteid="2031" externalid="387375">
              <RESULTS>
                <RESULT eventid="1101" points="89" swimtime="00:00:49.76" resultid="2032" heatid="2375" lane="7" />
                <RESULT eventid="1089" points="190" swimtime="00:01:21.44" resultid="2033" heatid="2361" lane="4" entrytime="00:01:26.64" entrycourse="LCM" />
                <RESULT eventid="1133" points="148" swimtime="00:01:37.39" resultid="2034" heatid="2419" lane="6" entrytime="00:01:36.63" entrycourse="LCM" />
                <RESULT eventid="1117" points="179" swimtime="00:06:30.04" resultid="2035" heatid="2394" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.80" />
                    <SPLIT distance="200" swimtime="00:03:10.12" />
                    <SPLIT distance="300" swimtime="00:04:51.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Julia Rocha" birthdate="2014-02-10" gender="F" nation="BRA" license="397158" swrid="5641767" athleteid="2075" externalid="397158">
              <RESULTS>
                <RESULT eventid="1092" points="224" swimtime="00:00:40.22" resultid="2076" heatid="2367" lane="6" entrytime="00:00:43.01" entrycourse="LCM" />
                <RESULT eventid="1064" points="238" swimtime="00:03:01.99" resultid="2077" heatid="2329" lane="5" entrytime="00:03:43.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="253" swimtime="00:00:42.43" resultid="2078" heatid="2405" lane="4" entrytime="00:00:42.70" entrycourse="LCM" />
                <RESULT eventid="1108" points="251" swimtime="00:03:19.73" resultid="2079" heatid="2384" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Faustino Canjerana" birthdate="2013-09-27" gender="F" nation="BRA" license="416735" athleteid="2146" externalid="416735">
              <RESULTS>
                <RESULT eventid="1098" points="205" swimtime="00:00:41.41" resultid="2147" heatid="2372" lane="7" />
                <RESULT eventid="1086" points="303" swimtime="00:01:16.97" resultid="2148" heatid="2354" lane="1" />
                <RESULT eventid="1130" points="182" swimtime="00:01:41.10" resultid="2149" heatid="2412" lane="7" />
                <RESULT eventid="1142" points="204" swimtime="00:00:49.51" resultid="2150" heatid="2430" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mathias" lastname="Lopes Batista" birthdate="2012-08-22" gender="M" nation="BRA" license="399740" swrid="5652889" athleteid="2090" externalid="399740">
              <RESULTS>
                <RESULT eventid="1089" points="150" swimtime="00:01:28.03" resultid="2091" heatid="2362" lane="6" entrytime="00:01:22.97" entrycourse="LCM" />
                <RESULT eventid="1133" points="172" swimtime="00:01:32.66" resultid="2092" heatid="2419" lane="3" entrytime="00:01:31.14" entrycourse="LCM" />
                <RESULT eventid="1145" points="47" swimtime="00:01:11.73" resultid="2093" heatid="2435" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Wenceslau Bitencourt" birthdate="2012-02-11" gender="M" nation="BRA" license="377318" swrid="5602591" athleteid="2002" externalid="377318">
              <RESULTS>
                <RESULT eventid="1101" points="214" swimtime="00:00:37.22" resultid="2003" heatid="2378" lane="7" entrytime="00:00:37.54" entrycourse="LCM" />
                <RESULT eventid="1073" points="197" swimtime="00:03:15.79" resultid="2004" heatid="2339" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="185" swimtime="00:01:30.49" resultid="2005" heatid="2420" lane="8" entrytime="00:01:29.08" entrycourse="LCM" />
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada.  (Horário: 19:18)" eventid="1145" status="DSQ" swimtime="00:00:51.00" resultid="2006" heatid="2435" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Barbosa Cortes" birthdate="2015-08-04" gender="M" nation="BRA" license="416977" athleteid="2160" externalid="416977">
              <RESULTS>
                <RESULT eventid="1127" points="44" swimtime="00:01:06.45" resultid="2161" heatid="2406" lane="5" />
                <RESULT eventid="1139" points="28" swimtime="00:01:08.44" resultid="2162" heatid="2425" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Ryan Rosa" birthdate="2014-01-14" gender="M" nation="BRA" license="400032" swrid="5652898" athleteid="2099" externalid="400032">
              <RESULTS>
                <RESULT eventid="1095" points="46" swimtime="00:01:01.92" resultid="2100" heatid="2368" lane="3" />
                <RESULT eventid="1083" points="121" swimtime="00:00:52.36" resultid="2101" heatid="2351" lane="3" entrytime="00:00:52.88" entrycourse="LCM" />
                <RESULT eventid="1127" points="114" swimtime="00:00:48.53" resultid="2102" heatid="2409" lane="4" entrytime="00:00:48.27" entrycourse="LCM" />
                <RESULT eventid="1139" points="145" swimtime="00:00:39.75" resultid="2103" heatid="2428" lane="1" entrytime="00:00:40.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Gouvea" birthdate="2013-04-19" gender="M" nation="BRA" license="387378" swrid="5588729" athleteid="2041" externalid="387378">
              <RESULTS>
                <RESULT eventid="1089" points="263" swimtime="00:01:13.05" resultid="2042" heatid="2362" lane="3" entrytime="00:01:22.66" entrycourse="LCM" />
                <RESULT eventid="1073" points="231" swimtime="00:03:05.61" resultid="2043" heatid="2340" lane="6" entrytime="00:03:11.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="233" swimtime="00:05:57.57" resultid="2044" heatid="2394" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.25" />
                    <SPLIT distance="200" swimtime="00:02:58.15" />
                    <SPLIT distance="300" swimtime="00:04:30.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="210" swimtime="00:00:43.59" resultid="2045" heatid="2437" lane="5" entrytime="00:00:49.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Vitor Vicente" birthdate="2012-09-20" gender="M" nation="BRA" license="415246" swrid="5755345" athleteid="2137" externalid="415246">
              <RESULTS>
                <RESULT eventid="1089" points="121" swimtime="00:01:34.58" resultid="2138" heatid="2359" lane="1" />
                <RESULT comment="SW 6.4 - A virada não foi iniciada após a conclusão do movimento de braço, após sair da posição de costas.  (Horário: 18:32), Na volta 50m." eventid="1133" status="DSQ" swimtime="00:02:00.16" resultid="2139" heatid="2417" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Prestes Alves Pinto" birthdate="2012-01-19" gender="F" nation="BRA" license="377324" swrid="5588867" athleteid="2007" externalid="377324">
              <RESULTS>
                <RESULT eventid="1086" points="351" swimtime="00:01:13.28" resultid="2008" heatid="2358" lane="6" entrytime="00:01:12.65" entrycourse="LCM" />
                <RESULT eventid="1070" points="309" swimtime="00:03:06.47" resultid="2009" heatid="2337" lane="6" entrytime="00:03:07.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="275" swimtime="00:01:28.09" resultid="2010" heatid="2415" lane="7" entrytime="00:01:25.74" entrycourse="LCM" />
                <RESULT eventid="1114" points="290" swimtime="00:05:55.48" resultid="2011" heatid="2392" lane="6" entrytime="00:06:05.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.93" />
                    <SPLIT distance="200" swimtime="00:02:52.82" />
                    <SPLIT distance="300" swimtime="00:04:26.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauren" lastname="Kurecki" birthdate="2014-03-06" gender="F" nation="BRA" license="377314" swrid="5602549" athleteid="1992" externalid="377314">
              <RESULTS>
                <RESULT eventid="1092" points="259" swimtime="00:00:38.28" resultid="1993" heatid="2367" lane="4" entrytime="00:00:37.95" entrycourse="LCM" />
                <RESULT eventid="1080" points="311" swimtime="00:00:43.00" resultid="1994" heatid="2348" lane="4" entrytime="00:00:44.66" entrycourse="LCM" />
                <RESULT eventid="1136" points="351" swimtime="00:00:33.45" resultid="1995" heatid="2424" lane="4" entrytime="00:00:33.61" entrycourse="LCM" />
                <RESULT eventid="1108" points="299" swimtime="00:03:08.47" resultid="1996" heatid="2385" lane="5" entrytime="00:03:36.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lis" lastname="Cristini Harmatiuk" birthdate="2014-07-19" gender="F" nation="BRA" license="396830" swrid="5641759" athleteid="2127" externalid="396830">
              <RESULTS>
                <RESULT eventid="1092" points="124" swimtime="00:00:48.91" resultid="2128" heatid="2367" lane="8" entrytime="00:00:47.43" entrycourse="LCM" />
                <RESULT eventid="1080" points="207" swimtime="00:00:49.24" resultid="2129" heatid="2348" lane="3" entrytime="00:00:50.37" entrycourse="LCM" />
                <RESULT eventid="1136" points="216" swimtime="00:00:39.30" resultid="2130" heatid="2424" lane="8" entrytime="00:00:39.67" entrycourse="LCM" />
                <RESULT eventid="1124" points="197" swimtime="00:00:46.15" resultid="2131" heatid="2405" lane="8" entrytime="00:00:47.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Soul Santos" birthdate="2016-05-11" gender="M" nation="BRA" license="415247" swrid="5755343" athleteid="2140" externalid="415247">
              <RESULTS>
                <RESULT eventid="1078" points="45" swimtime="00:01:06.04" resultid="2141" heatid="2344" lane="6" entrytime="00:01:03.93" entrycourse="LCM" />
                <RESULT eventid="1122" points="56" swimtime="00:00:54.44" resultid="2142" heatid="2401" lane="5" entrytime="00:00:58.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Everton" lastname="Rafael Guimaraes" birthdate="2015-08-25" gender="M" nation="BRA" license="416976" athleteid="2157" externalid="416976">
              <RESULTS>
                <RESULT eventid="1127" points="42" swimtime="00:01:07.37" resultid="2158" heatid="2407" lane="6" />
                <RESULT eventid="1139" points="48" swimtime="00:00:57.39" resultid="2159" heatid="2425" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Aparecida Lourenço Alves" birthdate="2013-11-06" gender="F" nation="BRA" license="387374" swrid="5588530" athleteid="2027" externalid="387374">
              <RESULTS>
                <RESULT eventid="1086" points="242" swimtime="00:01:22.87" resultid="2028" heatid="2355" lane="5" entrytime="00:01:39.44" entrycourse="LCM" />
                <RESULT eventid="1130" points="199" swimtime="00:01:38.19" resultid="2029" heatid="2412" lane="3" />
                <RESULT eventid="1142" points="173" swimtime="00:00:52.31" resultid="2030" heatid="2431" lane="6" entrytime="00:01:15.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Hoffmann Zoschke" birthdate="2015-03-22" gender="M" nation="BRA" license="390917" swrid="5602547" athleteid="2061" externalid="390917">
              <RESULTS>
                <RESULT eventid="1083" points="123" swimtime="00:00:52.10" resultid="2062" heatid="2352" lane="8" entrytime="00:00:51.70" entrycourse="LCM" />
                <RESULT eventid="1067" points="186" swimtime="00:02:58.42" resultid="2063" heatid="2334" lane="6" entrytime="00:03:01.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="160" swimtime="00:03:29.90" resultid="2064" heatid="2389" lane="2" entrytime="00:03:35.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="188" swimtime="00:00:36.47" resultid="2065" heatid="2428" lane="5" entrytime="00:00:37.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Zanotto De Souza" birthdate="2013-08-24" gender="M" nation="BRA" license="388361" swrid="5588974" athleteid="2056" externalid="388361">
              <RESULTS>
                <RESULT eventid="1089" points="244" swimtime="00:01:14.98" resultid="2057" heatid="2363" lane="4" entrytime="00:01:15.91" entrycourse="LCM" />
                <RESULT eventid="1073" points="205" swimtime="00:03:13.13" resultid="2058" heatid="2341" lane="1" entrytime="00:03:09.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="159" swimtime="00:01:35.17" resultid="2059" heatid="2418" lane="1" />
                <RESULT eventid="1117" points="245" swimtime="00:05:51.61" resultid="2060" heatid="2397" lane="1" entrytime="00:05:44.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.66" />
                    <SPLIT distance="200" swimtime="00:02:51.82" />
                    <SPLIT distance="300" swimtime="00:04:22.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Andrade Guarido" birthdate="2014-05-17" gender="M" nation="BRA" license="400031" swrid="5652873" athleteid="2094" externalid="400031">
              <RESULTS>
                <RESULT eventid="1095" points="57" swimtime="00:00:57.63" resultid="2095" heatid="2368" lane="4" entrytime="00:00:59.26" entrycourse="LCM" />
                <RESULT eventid="1083" points="125" swimtime="00:00:51.86" resultid="2096" heatid="2351" lane="6" entrytime="00:00:54.04" entrycourse="LCM" />
                <RESULT eventid="1111" points="126" swimtime="00:03:47.34" resultid="2097" heatid="2386" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:57.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="157" swimtime="00:00:38.73" resultid="2098" heatid="2428" lane="7" entrytime="00:00:39.19" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Vieira Coelho" birthdate="2014-09-28" gender="F" nation="BRA" license="406951" swrid="5717301" athleteid="2132" externalid="406951">
              <RESULTS>
                <RESULT eventid="1092" points="87" swimtime="00:00:55.11" resultid="2133" heatid="2366" lane="5" entrytime="00:00:50.21" entrycourse="LCM" />
                <RESULT eventid="1080" points="182" swimtime="00:00:51.39" resultid="2134" heatid="2348" lane="2" entrytime="00:00:52.06" entrycourse="LCM" />
                <RESULT eventid="1136" points="211" swimtime="00:00:39.60" resultid="2135" heatid="2424" lane="1" entrytime="00:00:38.67" entrycourse="LCM" />
                <RESULT eventid="1124" points="180" swimtime="00:00:47.57" resultid="2136" heatid="2402" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16131" nation="BRA" region="PR" clubid="1878" swrid="93766" name="Associação Nadar Colombo" shortname="Equipe Nadar">
          <ATHLETES>
            <ATHLETE firstname="Tayna" lastname="Macedo Gabardo" birthdate="2012-12-01" gender="F" nation="BRA" license="406704" swrid="5717281" athleteid="1879" externalid="406704">
              <RESULTS>
                <RESULT eventid="1098" points="168" swimtime="00:00:44.25" resultid="1880" heatid="2372" lane="3" />
                <RESULT eventid="1086" points="284" swimtime="00:01:18.58" resultid="1881" heatid="2354" lane="5" />
                <RESULT eventid="1130" points="239" swimtime="00:01:32.31" resultid="1882" heatid="2412" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13038" nation="BRA" region="PR" clubid="1186" swrid="93759" name="Associação De Pais E Atletas De Natação Ws/Crb" shortname="Apan/Ws">
          <ATHLETES>
            <ATHLETE firstname="Leon" lastname="Bernardo Bello" birthdate="2014-11-23" gender="M" nation="BRA" license="400324" swrid="5717246" athleteid="1209" externalid="400324">
              <RESULTS>
                <RESULT eventid="1095" points="67" swimtime="00:00:54.60" resultid="1210" heatid="2369" lane="8" entrytime="00:00:58.24" entrycourse="LCM" />
                <RESULT eventid="1083" points="130" swimtime="00:00:51.19" resultid="1211" heatid="2351" lane="5" entrytime="00:00:52.84" entrycourse="LCM" />
                <RESULT eventid="1127" points="144" swimtime="00:00:44.89" resultid="1212" heatid="2409" lane="5" entrytime="00:00:48.42" entrycourse="LCM" />
                <RESULT eventid="1139" points="164" swimtime="00:00:38.14" resultid="1213" heatid="2428" lane="6" entrytime="00:00:37.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Bernardi Iurk" birthdate="2012-04-14" gender="M" nation="BRA" license="408687" swrid="5725984" athleteid="1191" externalid="408687">
              <RESULTS>
                <RESULT eventid="1089" points="207" swimtime="00:01:19.11" resultid="1192" heatid="2361" lane="3" entrytime="00:01:27.74" entrycourse="LCM" />
                <RESULT eventid="1133" points="174" swimtime="00:01:32.31" resultid="1193" heatid="2418" lane="2" />
                <RESULT eventid="1145" points="162" swimtime="00:00:47.55" resultid="1194" heatid="2436" lane="6" entrytime="00:00:54.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Gramms Dallarosa" birthdate="2015-01-14" gender="F" nation="BRA" license="406868" swrid="5717270" athleteid="1219" externalid="406868">
              <RESULTS>
                <RESULT eventid="1080" points="97" swimtime="00:01:03.41" resultid="1220" heatid="2346" lane="4" entrytime="00:01:02.28" entrycourse="LCM" />
                <RESULT eventid="1136" points="132" swimtime="00:00:46.26" resultid="1221" heatid="2421" lane="4" entrytime="00:00:47.79" entrycourse="LCM" />
                <RESULT eventid="1124" points="118" swimtime="00:00:54.70" resultid="1222" heatid="2403" lane="2" entrytime="00:00:57.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Dos Santos" birthdate="2013-06-26" gender="F" nation="BRA" license="387512" swrid="5588662" athleteid="1200" externalid="387512">
              <RESULTS>
                <RESULT eventid="1098" points="154" swimtime="00:00:45.52" resultid="1201" heatid="2373" lane="7" entrytime="00:00:48.13" entrycourse="LCM" />
                <RESULT eventid="1086" points="281" swimtime="00:01:18.89" resultid="1202" heatid="2355" lane="6" entrytime="00:01:42.73" entrycourse="LCM" />
                <RESULT eventid="1130" points="202" swimtime="00:01:37.62" resultid="1203" heatid="2414" lane="1" entrytime="00:01:38.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Da Reginalda" birthdate="2012-11-09" gender="M" nation="BRA" license="400275" swrid="5717253" athleteid="1204" externalid="400275">
              <RESULTS>
                <RESULT eventid="1101" points="189" swimtime="00:00:38.78" resultid="1205" heatid="2375" lane="2" />
                <RESULT eventid="1089" points="247" swimtime="00:01:14.61" resultid="1206" heatid="2363" lane="6" entrytime="00:01:18.12" entrycourse="LCM" />
                <RESULT eventid="1133" points="256" swimtime="00:01:21.20" resultid="1207" heatid="2418" lane="4" />
                <RESULT eventid="1145" points="206" swimtime="00:00:43.87" resultid="1208" heatid="2436" lane="4" entrytime="00:00:52.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Bernardi Iurk" birthdate="2012-04-14" gender="M" nation="BRA" license="406940" swrid="5717245" athleteid="1187" externalid="406940">
              <RESULTS>
                <RESULT eventid="1101" points="172" swimtime="00:00:39.97" resultid="1188" heatid="2376" lane="7" />
                <RESULT eventid="1089" points="270" swimtime="00:01:12.42" resultid="1189" heatid="2361" lane="2" entrytime="00:01:27.99" entrycourse="LCM" />
                <RESULT eventid="1133" points="162" swimtime="00:01:34.47" resultid="1190" heatid="2419" lane="7" entrytime="00:01:43.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Ueda Pritzsche" birthdate="2012-02-07" gender="M" nation="BRA" license="417110" athleteid="1239" externalid="417110">
              <RESULTS>
                <RESULT eventid="1089" points="187" swimtime="00:01:21.86" resultid="1240" heatid="2359" lane="7" />
                <RESULT eventid="1133" points="169" swimtime="00:01:33.29" resultid="1241" heatid="2417" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Cravcenco Marcondes" birthdate="2012-06-23" gender="F" nation="BRA" license="406866" swrid="5725987" athleteid="1214" externalid="406866">
              <RESULTS>
                <RESULT eventid="1098" points="155" swimtime="00:00:45.42" resultid="1215" heatid="2372" lane="6" />
                <RESULT eventid="1086" points="231" swimtime="00:01:24.19" resultid="1216" heatid="2353" lane="3" />
                <RESULT eventid="1130" points="200" swimtime="00:01:38.02" resultid="1217" heatid="2413" lane="7" />
                <RESULT eventid="1142" points="228" swimtime="00:00:47.73" resultid="1218" heatid="2432" lane="6" entrytime="00:00:53.19" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Ferreira" birthdate="2012-12-29" gender="F" nation="BRA" license="382235" swrid="5602538" athleteid="1195" externalid="382235">
              <RESULTS>
                <RESULT eventid="1098" points="254" swimtime="00:00:38.53" resultid="1196" heatid="2374" lane="1" entrytime="00:00:41.41" entrycourse="LCM" />
                <RESULT eventid="1070" points="286" swimtime="00:03:11.32" resultid="1197" heatid="2335" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="269" swimtime="00:01:28.74" resultid="1198" heatid="2413" lane="4" entrytime="00:01:49.36" entrycourse="LCM" />
                <RESULT eventid="1142" points="180" swimtime="00:00:51.56" resultid="1199" heatid="2430" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Leopoldo Goncalves" birthdate="2015-01-10" gender="M" nation="BRA" license="417109" athleteid="1235" externalid="417109">
              <RESULTS>
                <RESULT eventid="1067" points="144" swimtime="00:03:14.16" resultid="1236" heatid="2331" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="157" swimtime="00:00:43.61" resultid="1237" heatid="2407" lane="2" />
                <RESULT eventid="1139" points="177" swimtime="00:00:37.21" resultid="1238" heatid="2425" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Ancai Freire" birthdate="2012-08-11" gender="M" nation="BRA" license="415258" swrid="5754925" athleteid="1226" externalid="415258">
              <RESULTS>
                <RESULT eventid="1089" points="106" swimtime="00:01:38.93" resultid="1227" heatid="2360" lane="1" />
                <RESULT eventid="1133" points="84" swimtime="00:01:57.61" resultid="1228" heatid="2416" lane="3" />
                <RESULT eventid="1145" points="88" swimtime="00:00:58.27" resultid="1229" heatid="2435" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Gabriel Cabral" birthdate="2014-02-11" gender="M" nation="BRA" license="415259" swrid="5755337" athleteid="1230" externalid="415259">
              <RESULTS>
                <RESULT eventid="1083" points="64" swimtime="00:01:04.83" resultid="1231" heatid="2349" lane="2" />
                <RESULT eventid="1067" points="143" swimtime="00:03:14.92" resultid="1232" heatid="2331" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="101" swimtime="00:00:50.42" resultid="1233" heatid="2409" lane="6" entrytime="00:00:49.57" entrycourse="LCM" />
                <RESULT eventid="1139" points="136" swimtime="00:00:40.62" resultid="1234" heatid="2427" lane="6" entrytime="00:00:41.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iasmim" lastname="Ferenczuk" birthdate="2013-06-06" gender="F" nation="BRA" license="414654" swrid="5755335" athleteid="1223" externalid="414654">
              <RESULTS>
                <RESULT eventid="1086" points="133" swimtime="00:01:41.20" resultid="1224" heatid="2354" lane="3" />
                <RESULT eventid="1142" points="123" swimtime="00:00:58.50" resultid="1225" heatid="2431" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
