<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.78979">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Foz do Iguaçu" name="Torneio Regional 3ª Região (Pré-Mirim/Sênior)" course="SCM" deadline="2024-02-21" entrystartdate="2024-02-19" entrytype="INVITATION" hostclub="Prefeitura Municipal de Foz do Iguaçu" hostclub.url="https://www.pmfi.pr.gov.br/" number="38297" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/evento/natacao/38297" startmethod="1" timing="AUTOMATIC" masters="F" withdrawuntil="2024-02-22" state="PR" nation="BRA">
      <AGEDATE value="2024-02-24" type="YEAR" />
      <POOL name="Ginásio de Esportes Costa Cavalcante" lanemin="1" lanemax="6" />
      <FACILITY city="Foz do Iguaçu" name="Ginásio de Esportes Costa Cavalcante" nation="BRA" state="PR" street="Rua Lisboa, 510" street2="Jardim Alice" zip="85858-050" />
      <POINTTABLE pointtableid="3016" name="FINA Point Scoring" version="2023" />
      <QUALIFY from="2023-02-24" until="2024-02-23" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-02-24" daytime="09:10" endtime="12:59" number="1" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1060" daytime="09:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1716" />
                    <RANKING order="2" place="2" resultid="1868" />
                    <RANKING order="3" place="3" resultid="1841" />
                    <RANKING order="4" place="4" resultid="1721" />
                    <RANKING order="5" place="5" resultid="1776" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1782" />
                    <RANKING order="2" place="2" resultid="1663" />
                    <RANKING order="3" place="3" resultid="1558" />
                    <RANKING order="4" place="4" resultid="1371" />
                    <RANKING order="5" place="5" resultid="1874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1669" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1705" />
                    <RANKING order="2" place="2" resultid="1657" />
                    <RANKING order="3" place="3" resultid="1436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1067" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1645" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1904" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1905" daytime="09:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1906" daytime="09:18" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1068" daytime="09:22" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1069" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1709" />
                    <RANKING order="2" place="2" resultid="1692" />
                    <RANKING order="3" place="3" resultid="1814" />
                    <RANKING order="4" place="4" resultid="1728" />
                    <RANKING order="5" place="5" resultid="1852" />
                    <RANKING order="6" place="6" resultid="1607" />
                    <RANKING order="7" place="-1" resultid="1767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1674" />
                    <RANKING order="2" place="2" resultid="1569" />
                    <RANKING order="3" place="3" resultid="1681" />
                    <RANKING order="4" place="-1" resultid="1788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1734" />
                    <RANKING order="2" place="2" resultid="1651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1639" />
                    <RANKING order="2" place="2" resultid="1491" />
                    <RANKING order="3" place="3" resultid="1795" />
                    <RANKING order="4" place="4" resultid="1747" />
                    <RANKING order="5" place="5" resultid="1456" />
                    <RANKING order="6" place="6" resultid="1522" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1687" />
                    <RANKING order="2" place="2" resultid="1516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1633" />
                    <RANKING order="2" place="2" resultid="1485" />
                    <RANKING order="3" place="3" resultid="1740" />
                    <RANKING order="4" place="-1" resultid="1474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1480" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1907" daytime="09:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1908" daytime="09:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1909" daytime="09:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="1910" daytime="09:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="1911" daytime="09:38" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1076" daytime="09:42" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1077" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1374" />
                    <RANKING order="2" place="-1" resultid="1628" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1534" />
                    <RANKING order="2" place="2" resultid="1836" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1912" daytime="09:42" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1079" daytime="09:46" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1080" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1805" />
                    <RANKING order="2" place="2" resultid="1564" />
                    <RANKING order="3" place="3" resultid="1752" />
                    <RANKING order="4" place="4" resultid="1575" />
                    <RANKING order="5" place="-1" resultid="1620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1699" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1913" daytime="09:46" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1082" daytime="09:50" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1083" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1402" />
                    <RANKING order="2" place="2" resultid="1624" />
                    <RANKING order="3" place="-1" resultid="1821" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1810" />
                    <RANKING order="2" place="2" resultid="1826" />
                    <RANKING order="3" place="3" resultid="1858" />
                    <RANKING order="4" place="4" resultid="1894" />
                    <RANKING order="5" place="5" resultid="1423" />
                    <RANKING order="6" place="6" resultid="1409" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1914" daytime="09:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1915" daytime="09:52" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1085" daytime="09:54" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1086" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1762" />
                    <RANKING order="2" place="2" resultid="1772" />
                    <RANKING order="3" place="3" resultid="1360" />
                    <RANKING order="4" place="4" resultid="1420" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1916" daytime="09:54" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1088" daytime="09:56" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1089" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1353" />
                    <RANKING order="2" place="2" resultid="1334" />
                    <RANKING order="3" place="3" resultid="1596" />
                    <RANKING order="4" place="-1" resultid="1615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1781" />
                    <RANKING order="2" place="2" resultid="1557" />
                    <RANKING order="3" place="3" resultid="1662" />
                    <RANKING order="4" place="4" resultid="1873" />
                    <RANKING order="5" place="5" resultid="1322" />
                    <RANKING order="6" place="6" resultid="1527" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1363" />
                    <RANKING order="2" place="2" resultid="1503" />
                    <RANKING order="3" place="3" resultid="1668" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1092" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1656" />
                    <RANKING order="2" place="2" resultid="1704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1094" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1461" />
                    <RANKING order="2" place="2" resultid="1442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1644" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1917" daytime="09:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1918" daytime="10:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1919" daytime="10:02" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1096" daytime="10:04" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1097" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1606" />
                    <RANKING order="2" place="2" resultid="1590" />
                    <RANKING order="3" place="3" resultid="1851" />
                    <RANKING order="4" place="4" resultid="1406" />
                    <RANKING order="5" place="5" resultid="1602" />
                    <RANKING order="6" place="-1" resultid="1383" />
                    <RANKING order="7" place="-1" resultid="1766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1539" />
                    <RANKING order="2" place="2" resultid="1568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1100" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1638" />
                    <RANKING order="2" place="2" resultid="1794" />
                    <RANKING order="3" place="3" resultid="1746" />
                    <RANKING order="4" place="4" resultid="1340" />
                    <RANKING order="5" place="5" resultid="1455" />
                    <RANKING order="6" place="6" resultid="1521" />
                    <RANKING order="7" place="7" resultid="1509" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1343" />
                    <RANKING order="2" place="2" resultid="1515" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1330" />
                    <RANKING order="2" place="2" resultid="1468" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1920" daytime="10:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1921" daytime="10:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1922" daytime="10:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="1923" daytime="10:12" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1104" daytime="10:14" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1105" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1533" />
                    <RANKING order="2" place="2" resultid="1835" />
                    <RANKING order="3" place="3" resultid="1831" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1924" daytime="10:14" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1107" daytime="10:20" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1108" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1804" />
                    <RANKING order="2" place="2" resultid="1563" />
                    <RANKING order="3" place="3" resultid="1751" />
                    <RANKING order="4" place="4" resultid="1548" />
                    <RANKING order="5" place="5" resultid="1757" />
                    <RANKING order="6" place="6" resultid="1574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1553" />
                    <RANKING order="2" place="2" resultid="1800" />
                    <RANKING order="3" place="3" resultid="1863" />
                    <RANKING order="4" place="4" resultid="1585" />
                    <RANKING order="5" place="5" resultid="1847" />
                    <RANKING order="6" place="-1" resultid="1698" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1925" daytime="10:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1926" daytime="10:26" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1110" daytime="10:30" gender="F" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1111" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="1112" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1545" />
                    <RANKING order="2" place="2" resultid="1857" />
                    <RANKING order="3" place="3" resultid="1580" />
                    <RANKING order="4" place="4" resultid="1893" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1927" daytime="10:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1113" daytime="10:34" gender="M" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1114" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1880" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1771" />
                    <RANKING order="2" place="2" resultid="1393" />
                    <RANKING order="3" place="3" resultid="1884" />
                    <RANKING order="4" place="4" resultid="1761" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1928" daytime="10:34" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1116" daytime="10:36" gender="F" number="13" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1117" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1722" />
                    <RANKING order="2" place="2" resultid="1717" />
                    <RANKING order="3" place="3" resultid="1777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1437" />
                    <RANKING order="2" place="2" resultid="1337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1122" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1929" daytime="10:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1930" daytime="10:58" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1124" daytime="11:22" gender="M" number="14" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1125" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1710" />
                    <RANKING order="2" place="2" resultid="1693" />
                    <RANKING order="3" place="3" resultid="1729" />
                    <RANKING order="4" place="4" resultid="1815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1675" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1492" />
                    <RANKING order="2" place="2" resultid="1510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1498" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1931" daytime="11:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1932" daytime="11:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1132" daytime="12:00" gender="F" number="15" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1133" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1352" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1134" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1136" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1137" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1138" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1441" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1139" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1933" daytime="12:00" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1140" daytime="12:04" gender="M" number="16" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1141" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1396" />
                    <RANKING order="2" place="2" resultid="1601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1143" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1144" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1145" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1146" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1147" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1934" daytime="12:04" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1148" daytime="12:06" gender="F" number="17" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1149" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1378" />
                    <RANKING order="2" place="2" resultid="1356" />
                    <RANKING order="3" place="3" resultid="1888" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1830" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1935" daytime="12:06" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1151" daytime="12:08" gender="M" number="18" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1152" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1547" />
                    <RANKING order="2" place="2" resultid="1756" />
                    <RANKING order="3" place="3" resultid="1389" />
                    <RANKING order="4" place="4" resultid="1619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1552" />
                    <RANKING order="2" place="2" resultid="1799" />
                    <RANKING order="3" place="3" resultid="1862" />
                    <RANKING order="4" place="4" resultid="1584" />
                    <RANKING order="5" place="5" resultid="1846" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1936" daytime="12:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1937" daytime="12:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1154" daytime="12:14" gender="F" number="19" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1155" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1623" />
                    <RANKING order="2" place="-1" resultid="1820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1544" />
                    <RANKING order="2" place="2" resultid="1809" />
                    <RANKING order="3" place="3" resultid="1825" />
                    <RANKING order="4" place="4" resultid="1579" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1938" daytime="12:14" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1157" daytime="12:16" gender="M" number="20" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1158" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1883" />
                    <RANKING order="2" place="2" resultid="1611" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1939" daytime="12:16" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1160" daytime="12:18" gender="F" number="21" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1161" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1715" />
                    <RANKING order="2" place="2" resultid="1867" />
                    <RANKING order="3" place="3" resultid="1840" />
                    <RANKING order="4" place="4" resultid="1775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1162" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1321" />
                    <RANKING order="2" place="2" resultid="1370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1163" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1164" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1703" />
                    <RANKING order="2" place="2" resultid="1435" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1167" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1940" daytime="12:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1941" daytime="12:20" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1168" daytime="12:24" gender="M" number="22" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1169" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1727" />
                    <RANKING order="2" place="2" resultid="1589" />
                    <RANKING order="3" place="-1" resultid="1382" />
                    <RANKING order="4" place="-1" resultid="1765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1538" />
                    <RANKING order="2" place="2" resultid="1787" />
                    <RANKING order="3" place="3" resultid="1680" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1733" />
                    <RANKING order="2" place="2" resultid="1650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1793" />
                    <RANKING order="2" place="2" resultid="1745" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1686" />
                    <RANKING order="2" place="2" resultid="1497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1632" />
                    <RANKING order="2" place="2" resultid="1739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1327" />
                    <RANKING order="2" place="2" resultid="1467" />
                    <RANKING order="3" place="3" resultid="1479" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1942" daytime="12:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1943" daytime="12:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1944" daytime="12:28" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1176" daytime="12:32" gender="F" number="23" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1177" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1333" />
                    <RANKING order="2" place="2" resultid="1595" />
                    <RANKING order="3" place="3" resultid="1614" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1179" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1180" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1181" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1182" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1183" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1945" daytime="12:32" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1184" daytime="12:34" gender="M" number="24" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1185" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1605" />
                    <RANKING order="2" place="2" resultid="1346" />
                    <RANKING order="3" place="3" resultid="1399" />
                    <RANKING order="4" place="4" resultid="1405" />
                    <RANKING order="5" place="5" resultid="1600" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1187" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1188" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1189" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1190" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1946" daytime="12:34" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-02-24" daytime="15:40" endtime="18:51" number="2" officialmeeting="15:00" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1192" daytime="15:40" gender="M" number="25" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1193" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1713" />
                    <RANKING order="2" place="2" resultid="1696" />
                    <RANKING order="3" place="3" resultid="1731" />
                    <RANKING order="4" place="4" resultid="1818" />
                    <RANKING order="5" place="5" resultid="1855" />
                    <RANKING order="6" place="6" resultid="1609" />
                    <RANKING order="7" place="7" resultid="1593" />
                    <RANKING order="8" place="-1" resultid="1769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1678" />
                    <RANKING order="2" place="2" resultid="1542" />
                    <RANKING order="3" place="3" resultid="1791" />
                    <RANKING order="4" place="4" resultid="1684" />
                    <RANKING order="5" place="5" resultid="1572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1654" />
                    <RANKING order="2" place="2" resultid="1737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1196" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1642" />
                    <RANKING order="2" place="2" resultid="1797" />
                    <RANKING order="3" place="3" resultid="1749" />
                    <RANKING order="4" place="4" resultid="1495" />
                    <RANKING order="5" place="5" resultid="1513" />
                    <RANKING order="6" place="6" resultid="1525" />
                    <RANKING order="7" place="7" resultid="1459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1197" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1690" />
                    <RANKING order="2" place="2" resultid="1501" />
                    <RANKING order="3" place="3" resultid="1519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1477" />
                    <RANKING order="2" place="2" resultid="1636" />
                    <RANKING order="3" place="3" resultid="1489" />
                    <RANKING order="4" place="-1" resultid="1743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1199" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1471" />
                    <RANKING order="2" place="2" resultid="1483" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1947" daytime="15:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1948" daytime="15:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1949" daytime="15:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="1950" daytime="16:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="1951" daytime="16:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="1952" daytime="16:16" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1200" daytime="16:22" gender="F" number="26" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1201" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1719" />
                    <RANKING order="2" place="2" resultid="1844" />
                    <RANKING order="3" place="3" resultid="1725" />
                    <RANKING order="4" place="4" resultid="1871" />
                    <RANKING order="5" place="5" resultid="1779" />
                    <RANKING order="6" place="6" resultid="1598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1666" />
                    <RANKING order="2" place="2" resultid="1785" />
                    <RANKING order="3" place="3" resultid="1531" />
                    <RANKING order="4" place="4" resultid="1323" />
                    <RANKING order="5" place="5" resultid="1561" />
                    <RANKING order="6" place="6" resultid="1877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1203" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1507" />
                    <RANKING order="2" place="2" resultid="1672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1204" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1660" />
                    <RANKING order="2" place="2" resultid="1707" />
                    <RANKING order="3" place="3" resultid="1439" />
                    <RANKING order="4" place="4" resultid="1338" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1205" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1206" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1465" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1648" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1953" daytime="16:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1954" daytime="16:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1955" daytime="16:36" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="1956" daytime="16:42" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1208" daytime="16:50" gender="F" number="27" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1209" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1210" daytime="16:50" gender="M" number="28" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1211" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1212" daytime="16:50" gender="F" number="29" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1213" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1823" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1387" />
                    <RANKING order="2" place="2" resultid="1812" />
                    <RANKING order="3" place="3" resultid="1860" />
                    <RANKING order="4" place="4" resultid="1582" />
                    <RANKING order="5" place="5" resultid="1828" />
                    <RANKING order="6" place="6" resultid="1896" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1957" daytime="16:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1958" daytime="16:52" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1215" daytime="16:54" gender="M" number="30" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1216" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="1217" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1773" />
                    <RANKING order="2" place="2" resultid="1886" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1959" daytime="16:54" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1218" daytime="16:56" gender="F" number="31" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1219" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1220" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1838" />
                    <RANKING order="2" place="2" resultid="1833" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1960" daytime="16:56" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1221" daytime="17:00" gender="M" number="32" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1222" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1550" />
                    <RANKING order="2" place="2" resultid="1754" />
                    <RANKING order="3" place="3" resultid="1759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1223" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1555" />
                    <RANKING order="2" place="2" resultid="1865" />
                    <RANKING order="3" place="-1" resultid="1849" />
                    <RANKING order="4" place="-1" resultid="1701" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1961" daytime="17:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1962" daytime="17:04" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1224" daytime="17:08" gender="F" number="33" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1225" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1415" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1963" daytime="17:08" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1226" daytime="17:10" gender="M" number="34" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1227" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1418" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1964" daytime="17:10" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1228" daytime="17:10" gender="F" number="35" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1229" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1778" />
                    <RANKING order="2" place="2" resultid="1870" />
                    <RANKING order="3" place="3" resultid="1843" />
                    <RANKING order="4" place="4" resultid="1335" />
                    <RANKING order="5" place="-1" resultid="1617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1784" />
                    <RANKING order="2" place="2" resultid="1665" />
                    <RANKING order="3" place="3" resultid="1876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1232" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1234" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1235" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1965" daytime="17:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1966" daytime="17:14" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1236" daytime="17:18" gender="M" number="36" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1237" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1712" />
                    <RANKING order="2" place="2" resultid="1730" />
                    <RANKING order="3" place="3" resultid="1854" />
                    <RANKING order="4" place="4" resultid="1817" />
                    <RANKING order="5" place="5" resultid="1407" />
                    <RANKING order="6" place="-1" resultid="1695" />
                    <RANKING order="7" place="-1" resultid="1768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1238" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1677" />
                    <RANKING order="2" place="2" resultid="1790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1239" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1736" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1240" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1494" />
                    <RANKING order="2" place="2" resultid="1748" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1689" />
                    <RANKING order="2" place="2" resultid="1518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1635" />
                    <RANKING order="2" place="2" resultid="1350" />
                    <RANKING order="3" place="3" resultid="1742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1243" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1967" daytime="17:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1968" daytime="17:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1969" daytime="17:22" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1244" daytime="17:26" gender="F" number="37" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1245" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1530" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1248" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1249" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1250" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1251" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1970" daytime="17:26" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1252" daytime="17:28" gender="M" number="38" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1253" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1592" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1254" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1683" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1255" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1653" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1256" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1257" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1344" />
                    <RANKING order="2" place="2" resultid="1500" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1258" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1470" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1971" daytime="17:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1972" daytime="17:30" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1260" daytime="17:32" gender="F" number="39" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1261" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1262" daytime="17:32" gender="M" number="40" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1263" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1264" daytime="17:32" gender="F" number="41" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1265" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1380" />
                    <RANKING order="2" place="2" resultid="1358" />
                    <RANKING order="3" place="3" resultid="1376" />
                    <RANKING order="4" place="4" resultid="1891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1536" />
                    <RANKING order="2" place="2" resultid="1837" />
                    <RANKING order="3" place="3" resultid="1832" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1973" daytime="17:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1974" daytime="17:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1267" daytime="17:38" gender="M" number="42" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1268" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1807" />
                    <RANKING order="2" place="2" resultid="1753" />
                    <RANKING order="3" place="3" resultid="1391" />
                    <RANKING order="4" place="-1" resultid="1566" />
                    <RANKING order="5" place="-1" resultid="1577" />
                    <RANKING order="6" place="-1" resultid="1758" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1269" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1802" />
                    <RANKING order="2" place="2" resultid="1864" />
                    <RANKING order="3" place="-1" resultid="1587" />
                    <RANKING order="4" place="-1" resultid="1700" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1975" daytime="17:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1976" daytime="17:42" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1270" daytime="17:44" gender="F" number="43" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1271" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1718" />
                    <RANKING order="2" place="2" resultid="1842" />
                    <RANKING order="3" place="3" resultid="1869" />
                    <RANKING order="4" place="4" resultid="1723" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1272" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1664" />
                    <RANKING order="2" place="2" resultid="1783" />
                    <RANKING order="3" place="3" resultid="1560" />
                    <RANKING order="4" place="4" resultid="1372" />
                    <RANKING order="5" place="5" resultid="1875" />
                    <RANKING order="6" place="6" resultid="1368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1273" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1670" />
                    <RANKING order="2" place="2" resultid="1506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1274" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1659" />
                    <RANKING order="2" place="2" resultid="1438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1276" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1647" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1977" daytime="17:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1978" daytime="17:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1979" daytime="17:50" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1278" daytime="17:54" gender="M" number="44" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1279" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1694" />
                    <RANKING order="2" place="2" resultid="1711" />
                    <RANKING order="3" place="3" resultid="1816" />
                    <RANKING order="4" place="4" resultid="1853" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1676" />
                    <RANKING order="2" place="2" resultid="1541" />
                    <RANKING order="3" place="3" resultid="1571" />
                    <RANKING order="4" place="4" resultid="1789" />
                    <RANKING order="5" place="5" resultid="1682" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1282" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1493" />
                    <RANKING order="2" place="2" resultid="1640" />
                    <RANKING order="3" place="3" resultid="1458" />
                    <RANKING order="4" place="4" resultid="1524" />
                    <RANKING order="5" place="5" resultid="1512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1283" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1688" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1284" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1476" />
                    <RANKING order="2" place="2" resultid="1488" />
                    <RANKING order="3" place="3" resultid="1634" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1328" />
                    <RANKING order="2" place="2" resultid="1469" />
                    <RANKING order="3" place="3" resultid="1482" />
                    <RANKING order="4" place="4" resultid="1453" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1980" daytime="17:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1981" daytime="17:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1982" daytime="18:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="1983" daytime="18:04" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1286" daytime="18:06" gender="F" number="45" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1287" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1414" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1984" daytime="18:06" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1288" daytime="18:08" gender="M" number="46" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1289" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1417" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1985" daytime="18:08" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1290" daytime="18:10" gender="F" number="47" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1291" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1403" />
                    <RANKING order="2" place="2" resultid="1625" />
                    <RANKING order="3" place="-1" resultid="1822" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1859" />
                    <RANKING order="2" place="2" resultid="1386" />
                    <RANKING order="3" place="3" resultid="1811" />
                    <RANKING order="4" place="4" resultid="1827" />
                    <RANKING order="5" place="5" resultid="1581" />
                    <RANKING order="6" place="6" resultid="1895" />
                    <RANKING order="7" place="7" resultid="1424" />
                    <RANKING order="8" place="8" resultid="1410" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1986" daytime="18:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1987" daytime="18:12" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1293" daytime="18:14" gender="M" number="48" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1294" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="1295" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1394" />
                    <RANKING order="2" place="2" resultid="1885" />
                    <RANKING order="3" place="3" resultid="1763" />
                    <RANKING order="4" place="4" resultid="1361" />
                    <RANKING order="5" place="5" resultid="1421" />
                    <RANKING order="6" place="6" resultid="1612" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1988" daytime="18:14" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1296" daytime="18:16" gender="F" number="49" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1297" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1629" />
                    <RANKING order="2" place="2" resultid="1379" />
                    <RANKING order="3" place="3" resultid="1357" />
                    <RANKING order="4" place="4" resultid="1375" />
                    <RANKING order="5" place="5" resultid="1890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1298" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1535" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1989" daytime="18:16" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1299" daytime="18:18" gender="M" number="50" order="26" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1300" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1549" />
                    <RANKING order="2" place="2" resultid="1806" />
                    <RANKING order="3" place="3" resultid="1565" />
                    <RANKING order="4" place="4" resultid="1576" />
                    <RANKING order="5" place="5" resultid="1621" />
                    <RANKING order="6" place="6" resultid="1390" />
                    <RANKING order="7" place="7" resultid="1412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1301" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1554" />
                    <RANKING order="2" place="2" resultid="1801" />
                    <RANKING order="3" place="3" resultid="1586" />
                    <RANKING order="4" place="4" resultid="1848" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1990" daytime="18:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1991" daytime="18:20" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1302" daytime="18:22" gender="F" number="51" order="27" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1303" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1354" />
                    <RANKING order="2" place="2" resultid="1597" />
                    <RANKING order="3" place="3" resultid="1616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1304" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1559" />
                    <RANKING order="2" place="2" resultid="1529" />
                    <RANKING order="3" place="3" resultid="1367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1305" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1364" />
                    <RANKING order="2" place="2" resultid="1505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1306" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1658" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1307" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1308" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1463" />
                    <RANKING order="2" place="2" resultid="1443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1309" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1646" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1992" daytime="18:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1993" daytime="18:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1994" daytime="18:26" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1310" daytime="18:28" gender="M" number="52" order="28" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1311" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1608" />
                    <RANKING order="2" place="2" resultid="1591" />
                    <RANKING order="3" place="3" resultid="1400" />
                    <RANKING order="4" place="4" resultid="1397" />
                    <RANKING order="5" place="5" resultid="1347" />
                    <RANKING order="6" place="-1" resultid="1384" />
                    <RANKING order="7" place="-1" resultid="1603" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1312" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1570" />
                    <RANKING order="2" place="2" resultid="1540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1313" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1314" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1457" />
                    <RANKING order="2" place="2" resultid="1796" />
                    <RANKING order="3" place="3" resultid="1341" />
                    <RANKING order="4" place="4" resultid="1523" />
                    <RANKING order="5" place="5" resultid="1511" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1315" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1499" />
                    <RANKING order="2" place="2" resultid="1517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1316" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1475" />
                    <RANKING order="2" place="2" resultid="1487" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1317" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1331" />
                    <RANKING order="2" place="2" resultid="1325" />
                    <RANKING order="3" place="3" resultid="1452" />
                    <RANKING order="4" place="4" resultid="1481" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1995" daytime="18:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1996" daytime="18:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1997" daytime="18:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="1998" daytime="18:34" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="3501" nation="BRA" region="PR" clubid="1319" swrid="93752" name="Ortega &amp; De Souza Jesus" shortname="Aquafoz">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Rorato" birthdate="2013-04-18" gender="F" nation="BRA" license="383851" swrid="5596936" athleteid="1377" externalid="383851">
              <RESULTS>
                <RESULT eventid="1148" points="181" swimtime="00:00:44.62" resultid="1378" heatid="1935" lane="3" entrytime="00:00:43.65" entrycourse="SCM" />
                <RESULT eventid="1296" points="206" swimtime="00:00:38.80" resultid="1379" heatid="1989" lane="4" entrytime="00:00:37.27" entrycourse="SCM" />
                <RESULT eventid="1264" points="173" swimtime="00:01:41.25" resultid="1380" heatid="1974" lane="3" entrytime="00:01:41.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Varela" birthdate="2010-05-20" gender="F" nation="BRA" license="365503" swrid="5596942" athleteid="1365" externalid="365503">
              <RESULTS>
                <RESULT eventid="1132" points="229" swimtime="00:00:41.25" resultid="1366" heatid="1933" lane="4" entrytime="00:00:41.38" entrycourse="SCM" />
                <RESULT eventid="1302" points="259" swimtime="00:00:35.94" resultid="1367" heatid="1993" lane="3" entrytime="00:00:34.77" entrycourse="SCM" />
                <RESULT eventid="1270" points="201" swimtime="00:01:33.60" resultid="1368" heatid="1977" lane="4" entrytime="00:01:31.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Wirtti" birthdate="2011-01-14" gender="M" nation="BRA" license="383854" swrid="4917570" athleteid="1381" externalid="383854">
              <RESULTS>
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="1382" heatid="1942" lane="3" />
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="1383" heatid="1921" lane="2" entrytime="00:01:15.61" entrycourse="SCM" />
                <RESULT eventid="1310" status="DNS" swimtime="00:00:00.00" resultid="1384" heatid="1996" lane="5" entrytime="00:00:32.87" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Benicio Martins" birthdate="2013-01-20" gender="M" nation="BRA" license="392831" swrid="5641752" athleteid="1388" externalid="392831">
              <RESULTS>
                <RESULT eventid="1151" points="83" swimtime="00:00:50.53" resultid="1389" heatid="1937" lane="5" entrytime="00:00:51.46" entrycourse="SCM" />
                <RESULT eventid="1299" points="93" swimtime="00:00:44.46" resultid="1390" heatid="1990" lane="4" entrytime="00:00:44.22" entrycourse="SCM" />
                <RESULT eventid="1267" points="74" swimtime="00:01:57.05" resultid="1391" heatid="1976" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Miguel Bogado" birthdate="2013-05-28" gender="M" nation="PRY" license="406649" athleteid="1411" externalid="406649">
              <RESULTS>
                <RESULT eventid="1299" points="45" swimtime="00:00:56.58" resultid="1412" heatid="1990" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="De Albuquerque" birthdate="2014-11-19" gender="F" nation="BRA" license="406648" athleteid="1408" externalid="406648">
              <RESULTS>
                <RESULT eventid="1082" points="32" swimtime="00:01:28.90" resultid="1409" heatid="1914" lane="2" />
                <RESULT eventid="1290" points="49" swimtime="00:01:02.43" resultid="1410" heatid="1986" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Dominguez Olivieski" birthdate="2011-04-27" gender="M" nation="BRA" license="405717" swrid="5664737" athleteid="1404" externalid="405717">
              <RESULTS>
                <RESULT eventid="1184" points="110" swimtime="00:00:52.00" resultid="1405" heatid="1946" lane="1" entrytime="00:00:52.53" entrycourse="SCM" />
                <RESULT eventid="1096" points="156" swimtime="00:01:23.22" resultid="1406" heatid="1920" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="125" swimtime="00:01:50.29" resultid="1407" heatid="1967" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Franco" birthdate="2010-06-09" gender="F" nation="BRA" license="383849" swrid="5596896" athleteid="1320" externalid="383849">
              <RESULTS>
                <RESULT eventid="1160" points="239" swimtime="00:01:27.00" resultid="1321" heatid="1941" lane="1" entrytime="00:01:25.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="328" swimtime="00:01:12.79" resultid="1322" heatid="1918" lane="1" entrytime="00:01:13.24" entrycourse="SCM" />
                <RESULT eventid="1200" points="342" swimtime="00:05:30.74" resultid="1323" heatid="1954" lane="3" entrytime="00:05:35.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="100" swimtime="00:01:17.68" />
                    <SPLIT distance="150" swimtime="00:02:00.03" />
                    <SPLIT distance="200" swimtime="00:02:42.40" />
                    <SPLIT distance="250" swimtime="00:03:25.40" />
                    <SPLIT distance="300" swimtime="00:04:07.49" />
                    <SPLIT distance="350" swimtime="00:04:50.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Voltolini" birthdate="2014-06-29" gender="M" nation="BRA" license="383846" swrid="5596947" athleteid="1359" externalid="383846">
              <RESULTS>
                <RESULT eventid="1085" points="82" swimtime="00:00:57.31" resultid="1360" heatid="1916" lane="2" entrytime="00:00:58.35" entrycourse="SCM" />
                <RESULT eventid="1293" points="87" swimtime="00:00:45.40" resultid="1361" heatid="1988" lane="2" entrytime="00:00:44.07" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julio" lastname="Heck" birthdate="1998-02-15" gender="M" nation="BRA" license="185880" swrid="5596906" athleteid="1329" externalid="185880">
              <RESULTS>
                <RESULT eventid="1096" points="538" swimtime="00:00:55.11" resultid="1330" heatid="1923" lane="3" entrytime="00:00:52.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="515" swimtime="00:00:25.15" resultid="1331" heatid="1998" lane="3" entrytime="00:00:23.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yago" lastname="Simon Pires" birthdate="2008-10-29" gender="M" nation="BRA" license="328942" swrid="5596939" athleteid="1339" externalid="328942">
              <RESULTS>
                <RESULT eventid="1096" points="429" swimtime="00:00:59.45" resultid="1340" heatid="1922" lane="3" entrytime="00:00:59.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="402" swimtime="00:00:27.31" resultid="1341" heatid="1998" lane="6" entrytime="00:00:27.09" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Geórgia" lastname="Adeli Jesus" birthdate="2008-03-27" gender="F" nation="BRA" license="312649" swrid="5596864" athleteid="1336" externalid="312649">
              <RESULTS>
                <RESULT eventid="1116" points="352" swimtime="00:21:25.63" resultid="1337" heatid="1930" lane="4" entrytime="00:21:19.46" entrycourse="SCM" />
                <RESULT eventid="1200" points="393" swimtime="00:05:15.77" resultid="1338" heatid="1955" lane="5" entrytime="00:05:21.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="100" swimtime="00:01:14.41" />
                    <SPLIT distance="150" swimtime="00:01:54.06" />
                    <SPLIT distance="200" swimtime="00:02:34.35" />
                    <SPLIT distance="250" swimtime="00:03:14.28" />
                    <SPLIT distance="300" swimtime="00:03:55.30" />
                    <SPLIT distance="350" swimtime="00:04:35.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Gabriel Serighelli" birthdate="1999-03-12" gender="M" nation="BRA" license="121253" swrid="5596899" athleteid="1324" externalid="121253">
              <RESULTS>
                <RESULT eventid="1310" points="486" swimtime="00:00:25.64" resultid="1325" heatid="1998" lane="4" entrytime="00:00:24.09" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Mussi" birthdate="2006-12-31" gender="M" nation="BRA" license="370567" swrid="5596917" athleteid="1348" externalid="370567">
              <RESULTS>
                <RESULT eventid="1184" points="417" swimtime="00:00:33.37" resultid="1349" heatid="1946" lane="3" entrytime="00:00:32.05" entrycourse="SCM" />
                <RESULT eventid="1236" points="380" swimtime="00:01:16.28" resultid="1350" heatid="1969" lane="4" entrytime="00:01:12.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Marques Lima" birthdate="2010-04-30" gender="F" nation="BRA" license="383051" swrid="5596913" athleteid="1369" externalid="383051">
              <RESULTS>
                <RESULT eventid="1160" points="205" swimtime="00:01:31.54" resultid="1370" heatid="1941" lane="6" entrytime="00:01:28.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="265" swimtime="00:03:09.65" resultid="1371" heatid="1904" lane="4" entrytime="00:03:08.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                    <SPLIT distance="100" swimtime="00:01:26.02" />
                    <SPLIT distance="150" swimtime="00:02:24.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="300" swimtime="00:01:21.99" resultid="1372" heatid="1978" lane="3" entrytime="00:01:20.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Afonso Proteti" birthdate="2002-03-19" gender="M" nation="BRA" license="190464" swrid="5596865" athleteid="1326" externalid="190464">
              <RESULTS>
                <RESULT eventid="1168" points="642" swimtime="00:00:55.37" resultid="1327" heatid="1944" lane="3" entrytime="00:00:55.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="574" swimtime="00:00:58.15" resultid="1328" heatid="1983" lane="3" entrytime="00:00:57.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Garcete" birthdate="2014-01-04" gender="F" nation="BRA" license="383856" swrid="5596904" athleteid="1385" externalid="383856">
              <RESULTS>
                <RESULT eventid="1290" points="175" swimtime="00:00:40.95" resultid="1386" heatid="1987" lane="2" entrytime="00:00:41.24" entrycourse="SCM" />
                <RESULT eventid="1212" points="154" swimtime="00:00:45.48" resultid="1387" heatid="1958" lane="3" entrytime="00:00:45.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Otremba Rouver" birthdate="2007-04-25" gender="M" nation="BRA" license="342152" swrid="5596919" athleteid="1342" externalid="342152">
              <RESULTS>
                <RESULT eventid="1096" points="470" swimtime="00:00:57.67" resultid="1343" heatid="1923" lane="5" entrytime="00:00:56.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="497" swimtime="00:00:27.44" resultid="1344" heatid="1972" lane="2" entrytime="00:00:28.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauan" lastname="Matheus Cunha" birthdate="2011-01-31" gender="M" nation="BRA" license="392834" swrid="5641770" athleteid="1395" externalid="392834">
              <RESULTS>
                <RESULT eventid="1140" points="118" swimtime="00:00:45.04" resultid="1396" heatid="1934" lane="3" entrytime="00:00:45.07" entrycourse="SCM" />
                <RESULT eventid="1310" points="171" swimtime="00:00:36.26" resultid="1397" heatid="1995" lane="3" entrytime="00:00:38.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karim" lastname="Maruan Jaber" birthdate="2014-11-19" gender="M" nation="BRA" license="392833" swrid="5627304" athleteid="1392" externalid="392833">
              <RESULTS>
                <RESULT eventid="1113" points="106" swimtime="00:01:34.58" resultid="1393" heatid="1928" lane="4" entrytime="00:01:38.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1293" points="109" swimtime="00:00:42.08" resultid="1394" heatid="1988" lane="3" entrytime="00:00:41.23" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Blume" birthdate="2013-07-17" gender="F" nation="BRA" license="383850" swrid="5596873" athleteid="1373" externalid="383850">
              <RESULTS>
                <RESULT eventid="1076" points="128" swimtime="00:02:03.73" resultid="1374" heatid="1912" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="139" swimtime="00:00:44.16" resultid="1375" heatid="1989" lane="5" entrytime="00:00:45.81" entrycourse="SCM" />
                <RESULT eventid="1264" points="131" swimtime="00:01:51.24" resultid="1376" heatid="1974" lane="5" entrytime="00:01:57.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Victoria Portela" birthdate="2009-12-04" gender="F" nation="BRA" license="383047" swrid="5596945" athleteid="1362" externalid="383047">
              <RESULTS>
                <RESULT eventid="1088" points="409" swimtime="00:01:07.67" resultid="1363" heatid="1919" lane="1" entrytime="00:01:07.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="432" swimtime="00:00:30.33" resultid="1364" heatid="1994" lane="2" entrytime="00:00:30.06" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emma" lastname="Raquel Nascimento" birthdate="2015-11-06" gender="F" nation="BRA" license="392837" swrid="5641775" athleteid="1401" externalid="392837">
              <RESULTS>
                <RESULT eventid="1082" points="146" swimtime="00:00:53.78" resultid="1402" heatid="1915" lane="3" entrytime="00:00:55.31" entrycourse="SCM" />
                <RESULT eventid="1290" points="138" swimtime="00:00:44.30" resultid="1403" heatid="1987" lane="5" entrytime="00:00:43.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vicente" lastname="Duarte Martins" birthdate="2014-12-23" gender="M" nation="BRA" license="406654" athleteid="1419" externalid="406654">
              <RESULTS>
                <RESULT eventid="1085" points="20" swimtime="00:01:31.16" resultid="1420" heatid="1916" lane="1" />
                <RESULT eventid="1293" points="30" swimtime="00:01:04.88" resultid="1421" heatid="1988" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ian" lastname="Peroni Ottomar" birthdate="2016-07-15" gender="M" nation="BRA" license="406653" athleteid="1416" externalid="406653">
              <RESULTS>
                <RESULT eventid="1288" points="30" swimtime="00:00:29.22" resultid="1417" heatid="1985" lane="3" />
                <RESULT eventid="1226" points="52" swimtime="00:00:27.53" resultid="1418" heatid="1964" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gino" lastname="Benicio Ciallella" birthdate="2012-05-21" gender="M" nation="ARG" license="406735" athleteid="1425" externalid="406735">
              <RESULTS>
                <RESULT eventid="1299" points="34" status="EXH" swimtime="00:01:01.83" resultid="1426" heatid="1990" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daiana" lastname="Safadi Fakih" birthdate="2016-01-16" gender="F" nation="BRA" license="406650" athleteid="1413" externalid="406650">
              <RESULTS>
                <RESULT eventid="1286" points="66" swimtime="00:00:25.84" resultid="1414" heatid="1984" lane="3" />
                <RESULT eventid="1224" points="64" swimtime="00:00:29.63" resultid="1415" heatid="1963" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Maguet" birthdate="2011-07-01" gender="F" nation="BRA" license="370568" swrid="5596911" athleteid="1351" externalid="370568">
              <RESULTS>
                <RESULT eventid="1132" points="200" swimtime="00:00:43.15" resultid="1352" heatid="1933" lane="2" entrytime="00:00:47.52" entrycourse="SCM" />
                <RESULT eventid="1088" points="225" swimtime="00:01:22.59" resultid="1353" heatid="1917" lane="4" entrytime="00:01:25.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="238" swimtime="00:00:37.00" resultid="1354" heatid="1993" lane="4" entrytime="00:00:38.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Gustavo Cunha" birthdate="2011-01-31" gender="M" nation="BRA" license="392836" swrid="5641764" athleteid="1398" externalid="392836">
              <RESULTS>
                <RESULT eventid="1184" points="143" swimtime="00:00:47.71" resultid="1399" heatid="1946" lane="2" entrytime="00:00:45.74" entrycourse="SCM" />
                <RESULT eventid="1310" points="188" swimtime="00:00:35.16" resultid="1400" heatid="1996" lane="6" entrytime="00:00:35.59" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Mendes Portela" birthdate="2014-03-08" gender="F" nation="BRA" license="406656" athleteid="1422" externalid="406656">
              <RESULTS>
                <RESULT eventid="1082" points="42" swimtime="00:01:21.00" resultid="1423" heatid="1915" lane="6" />
                <RESULT eventid="1290" points="51" swimtime="00:01:01.66" resultid="1424" heatid="1986" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Pires" birthdate="2011-04-09" gender="F" nation="BRA" license="383853" swrid="5596927" athleteid="1332" externalid="383853">
              <RESULTS>
                <RESULT eventid="1176" points="193" swimtime="00:00:49.08" resultid="1333" heatid="1945" lane="3" entrytime="00:00:52.06" entrycourse="SCM" />
                <RESULT eventid="1088" points="169" swimtime="00:01:30.75" resultid="1334" heatid="1917" lane="2" entrytime="00:01:32.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="191" swimtime="00:01:48.28" resultid="1335" heatid="1965" lane="3" entrytime="00:01:48.01" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Xavier" birthdate="2011-10-14" gender="M" nation="BRA" license="370564" swrid="5596949" athleteid="1345" externalid="370564">
              <RESULTS>
                <RESULT eventid="1184" points="174" swimtime="00:00:44.69" resultid="1346" heatid="1946" lane="5" entrytime="00:00:46.12" entrycourse="SCM" />
                <RESULT eventid="1310" points="147" swimtime="00:00:38.16" resultid="1347" heatid="1995" lane="4" entrytime="00:00:38.99" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Murakami" birthdate="2013-11-24" gender="F" nation="BRA" license="383844" swrid="5596916" athleteid="1355" externalid="383844">
              <RESULTS>
                <RESULT eventid="1148" points="141" swimtime="00:00:48.47" resultid="1356" heatid="1935" lane="4" entrytime="00:00:48.18" entrycourse="SCM" />
                <RESULT eventid="1296" points="167" swimtime="00:00:41.62" resultid="1357" heatid="1989" lane="2" entrytime="00:00:41.88" entrycourse="SCM" />
                <RESULT eventid="1264" points="169" swimtime="00:01:42.19" resultid="1358" heatid="1974" lane="4" entrytime="00:01:49.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18151" nation="BRA" region="PR" clubid="1626" name="Clube Uniao Recreativo Palmense" shortname="Clube União">
          <ATHLETES>
            <ATHLETE firstname="Luiza" lastname="Langaro Spaniol" birthdate="2013-06-18" gender="F" nation="BRA" license="406600" athleteid="1627" externalid="406600">
              <RESULTS>
                <RESULT eventid="1076" status="DSQ" swimtime="00:01:36.70" resultid="1628" heatid="1912" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="276" swimtime="00:00:35.19" resultid="1629" heatid="1989" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13025" nation="BRA" region="PR" clubid="1433" swrid="93779" name="Instituto Desportos Aquáticos De Foz Do Iguaçu" shortname="Cataratas Natação">
          <ATHLETES>
            <ATHLETE firstname="Vitor" lastname="Marques Petry" birthdate="2008-01-08" gender="M" nation="BRA" license="392352" swrid="4795316" athleteid="1520" externalid="392352" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1096" points="344" swimtime="00:01:03.99" resultid="1521" heatid="1922" lane="1" entrytime="00:01:04.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="292" swimtime="00:02:45.16" resultid="1522" heatid="1908" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:18.55" />
                    <SPLIT distance="150" swimtime="00:02:08.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="331" swimtime="00:00:29.12" resultid="1523" heatid="1997" lane="5" entrytime="00:00:29.13" entrycourse="SCM" />
                <RESULT eventid="1278" points="249" swimtime="00:01:16.77" resultid="1524" heatid="1981" lane="5" entrytime="00:01:16.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="316" swimtime="00:05:11.48" resultid="1525" heatid="1949" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                    <SPLIT distance="100" swimtime="00:01:14.04" />
                    <SPLIT distance="150" swimtime="00:01:53.15" />
                    <SPLIT distance="200" swimtime="00:02:33.09" />
                    <SPLIT distance="250" swimtime="00:03:13.33" />
                    <SPLIT distance="300" swimtime="00:03:52.33" />
                    <SPLIT distance="350" swimtime="00:04:32.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Christopher" lastname="De Araujo" birthdate="2008-08-09" gender="M" nation="BRA" license="366376" swrid="5596884" athleteid="1490" externalid="366376" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1068" points="456" swimtime="00:02:22.43" resultid="1491" heatid="1911" lane="5" entrytime="00:02:23.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                    <SPLIT distance="100" swimtime="00:01:08.93" />
                    <SPLIT distance="150" swimtime="00:01:48.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="473" swimtime="00:18:06.87" resultid="1492" heatid="1931" lane="3" />
                <RESULT eventid="1278" points="366" swimtime="00:01:07.51" resultid="1493" heatid="1983" lane="6" entrytime="00:01:06.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="423" swimtime="00:01:13.62" resultid="1494" heatid="1969" lane="3" entrytime="00:01:12.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="427" swimtime="00:04:41.79" resultid="1495" heatid="1952" lane="2" entrytime="00:04:24.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                    <SPLIT distance="100" swimtime="00:01:04.91" />
                    <SPLIT distance="150" swimtime="00:01:41.29" />
                    <SPLIT distance="200" swimtime="00:02:18.22" />
                    <SPLIT distance="250" swimtime="00:02:54.30" />
                    <SPLIT distance="300" swimtime="00:03:31.22" />
                    <SPLIT distance="350" swimtime="00:04:06.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Marques Petry" birthdate="2008-01-08" gender="M" nation="BRA" license="392351" swrid="4711489" athleteid="1508" externalid="392351" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1096" points="327" swimtime="00:01:05.03" resultid="1509" heatid="1922" lane="6" entrytime="00:01:06.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="299" swimtime="00:21:05.13" resultid="1510" heatid="1931" lane="4" />
                <RESULT eventid="1310" points="304" swimtime="00:00:29.95" resultid="1511" heatid="1996" lane="3" entrytime="00:00:29.77" entrycourse="SCM" />
                <RESULT eventid="1278" points="197" swimtime="00:01:22.94" resultid="1512" heatid="1980" lane="3" entrytime="00:01:23.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="326" swimtime="00:05:08.20" resultid="1513" heatid="1949" lane="3" entrytime="00:05:20.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                    <SPLIT distance="100" swimtime="00:01:14.07" />
                    <SPLIT distance="150" swimtime="00:01:53.12" />
                    <SPLIT distance="200" swimtime="00:02:33.70" />
                    <SPLIT distance="250" swimtime="00:03:13.50" />
                    <SPLIT distance="300" swimtime="00:03:52.30" />
                    <SPLIT distance="350" swimtime="00:04:31.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="De Assis Santos" birthdate="2003-02-21" gender="M" nation="BRA" license="342496" swrid="5596885" athleteid="1478" externalid="342496" level="INTERNE/IT">
              <RESULTS>
                <RESULT eventid="1168" points="359" swimtime="00:01:07.20" resultid="1479" heatid="1942" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="369" swimtime="00:02:32.78" resultid="1480" heatid="1910" lane="5" entrytime="00:02:30.24" entrycourse="SCM" />
                <RESULT eventid="1310" points="433" swimtime="00:00:26.63" resultid="1481" heatid="1997" lane="4" entrytime="00:00:27.37" entrycourse="SCM" />
                <RESULT eventid="1278" points="399" swimtime="00:01:05.62" resultid="1482" heatid="1983" lane="2" entrytime="00:01:02.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="391" swimtime="00:04:50.23" resultid="1483" heatid="1947" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                    <SPLIT distance="100" swimtime="00:01:07.03" />
                    <SPLIT distance="150" swimtime="00:01:43.12" />
                    <SPLIT distance="200" swimtime="00:02:20.29" />
                    <SPLIT distance="250" swimtime="00:02:57.81" />
                    <SPLIT distance="300" swimtime="00:03:35.73" />
                    <SPLIT distance="350" swimtime="00:04:14.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Ferrari Ghellere" birthdate="2014-07-01" gender="F" nation="BRA" license="372038" swrid="5596895" athleteid="1543" externalid="372038" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1154" points="151" swimtime="00:00:47.32" resultid="1544" heatid="1938" lane="4" entrytime="00:00:53.12" entrycourse="SCM" />
                <RESULT eventid="1110" points="196" swimtime="00:01:26.41" resultid="1545" heatid="1927" lane="3" entrytime="00:01:27.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Axel" lastname="Ariel Giménez González" birthdate="2011-06-01" gender="M" nation="BRA" license="365755" swrid="5676299" athleteid="1604" externalid="365755" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1184" points="257" swimtime="00:00:39.21" resultid="1605" heatid="1946" lane="4" entrytime="00:00:43.53" entrycourse="SCM" />
                <RESULT eventid="1096" points="268" swimtime="00:01:09.53" resultid="1606" heatid="1921" lane="4" entrytime="00:01:11.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="222" swimtime="00:03:00.90" resultid="1607" heatid="1907" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="100" swimtime="00:01:27.21" />
                    <SPLIT distance="150" swimtime="00:02:19.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="288" swimtime="00:00:30.52" resultid="1608" heatid="1996" lane="4" entrytime="00:00:30.84" entrycourse="SCM" />
                <RESULT eventid="1192" points="221" swimtime="00:05:50.98" resultid="1609" heatid="1948" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:01:22.82" />
                    <SPLIT distance="150" swimtime="00:02:08.56" />
                    <SPLIT distance="200" swimtime="00:02:55.36" />
                    <SPLIT distance="250" swimtime="00:03:40.66" />
                    <SPLIT distance="300" swimtime="00:04:24.35" />
                    <SPLIT distance="350" swimtime="00:05:08.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Roza" birthdate="2013-06-05" gender="M" nation="BRA" license="374412" swrid="5588949" athleteid="1546" externalid="374412" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1151" points="153" swimtime="00:00:41.28" resultid="1547" heatid="1937" lane="2" entrytime="00:00:49.21" entrycourse="SCM" />
                <RESULT eventid="1107" points="205" swimtime="00:02:48.49" resultid="1548" heatid="1926" lane="2" entrytime="00:02:50.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                    <SPLIT distance="100" swimtime="00:01:21.70" />
                    <SPLIT distance="150" swimtime="00:02:08.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="226" swimtime="00:00:33.05" resultid="1549" heatid="1991" lane="4" entrytime="00:00:33.19" entrycourse="SCM" />
                <RESULT eventid="1221" points="130" swimtime="00:01:34.14" resultid="1550" heatid="1961" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joshua" lastname="Davalos Gimenez" birthdate="2013-10-22" gender="M" nation="PRY" license="380598" athleteid="1562" externalid="380598" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1107" points="206" swimtime="00:02:48.04" resultid="1563" heatid="1926" lane="4" entrytime="00:02:44.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                    <SPLIT distance="100" swimtime="00:01:21.54" />
                    <SPLIT distance="150" swimtime="00:02:06.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="188" swimtime="00:01:36.40" resultid="1564" heatid="1913" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="180" swimtime="00:00:35.69" resultid="1565" heatid="1991" lane="5" entrytime="00:00:35.40" entrycourse="SCM" />
                <RESULT eventid="1267" status="DSQ" swimtime="00:01:35.12" resultid="1566" heatid="1976" lane="2" entrytime="00:01:36.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Sermidi" birthdate="2005-06-15" gender="F" nation="BRA" license="283035" swrid="5596938" athleteid="1440" externalid="283035" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1132" points="393" swimtime="00:00:34.47" resultid="1441" heatid="1933" lane="3" entrytime="00:00:33.22" entrycourse="SCM" />
                <RESULT eventid="1088" points="432" swimtime="00:01:06.43" resultid="1442" heatid="1919" lane="2" entrytime="00:01:06.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="418" swimtime="00:00:30.66" resultid="1443" heatid="1994" lane="4" entrytime="00:00:29.18" entrycourse="SCM" />
                <RESULT eventid="1244" points="367" swimtime="00:00:34.03" resultid="1444" heatid="1970" lane="4" entrytime="00:00:31.38" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ysadora" lastname="Bertoldo" birthdate="2010-04-09" gender="F" nation="BRA" license="376444" swrid="5588553" athleteid="1526" externalid="376444" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1088" points="318" swimtime="00:01:13.58" resultid="1527" heatid="1918" lane="6" entrytime="00:01:14.63" entrycourse="SCM" />
                <RESULT eventid="1116" points="375" swimtime="00:20:58.87" resultid="1528" heatid="1930" lane="2" />
                <RESULT eventid="1302" points="262" swimtime="00:00:35.82" resultid="1529" heatid="1994" lane="6" entrytime="00:00:34.24" entrycourse="SCM" />
                <RESULT eventid="1244" points="256" swimtime="00:00:38.35" resultid="1530" heatid="1970" lane="5" />
                <RESULT eventid="1200" points="359" swimtime="00:05:25.32" resultid="1531" heatid="1955" lane="6" entrytime="00:05:32.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                    <SPLIT distance="100" swimtime="00:01:19.09" />
                    <SPLIT distance="150" swimtime="00:02:00.86" />
                    <SPLIT distance="200" swimtime="00:02:42.35" />
                    <SPLIT distance="250" swimtime="00:03:24.31" />
                    <SPLIT distance="300" swimtime="00:04:05.54" />
                    <SPLIT distance="350" swimtime="00:04:46.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrieli" lastname="Brietzke Sbardelatti" birthdate="2014-07-14" gender="F" nation="BRA" license="400456" swrid="4379861" athleteid="1578" externalid="400456" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1154" points="96" swimtime="00:00:54.99" resultid="1579" heatid="1938" lane="2" entrytime="00:00:53.84" entrycourse="SCM" />
                <RESULT eventid="1110" points="129" swimtime="00:01:39.25" resultid="1580" heatid="1927" lane="2" entrytime="00:01:48.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="132" swimtime="00:00:45.01" resultid="1581" heatid="1986" lane="3" entrytime="00:00:47.82" entrycourse="SCM" />
                <RESULT eventid="1212" points="83" swimtime="00:00:55.83" resultid="1582" heatid="1958" lane="5" entrytime="00:00:58.89" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Leticia Sbardelatti" birthdate="2011-07-28" gender="F" nation="BRA" license="403147" swrid="5676303" athleteid="1594" externalid="403147" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1176" points="182" swimtime="00:00:49.97" resultid="1595" heatid="1945" lane="2" />
                <RESULT eventid="1088" points="167" swimtime="00:01:31.13" resultid="1596" heatid="1917" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="197" swimtime="00:00:39.36" resultid="1597" heatid="1993" lane="2" entrytime="00:00:43.34" entrycourse="SCM" />
                <RESULT eventid="1200" points="127" swimtime="00:07:39.15" resultid="1598" heatid="1953" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.10" />
                    <SPLIT distance="100" swimtime="00:01:43.63" />
                    <SPLIT distance="150" swimtime="00:02:42.64" />
                    <SPLIT distance="200" swimtime="00:03:40.69" />
                    <SPLIT distance="250" swimtime="00:04:40.30" />
                    <SPLIT distance="300" swimtime="00:05:41.39" />
                    <SPLIT distance="350" swimtime="00:06:42.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="De Souza Tulio" birthdate="2006-06-23" gender="F" nation="BRA" license="342344" swrid="5030980" athleteid="1460" externalid="342344" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1088" points="566" swimtime="00:01:00.73" resultid="1461" heatid="1919" lane="3" entrytime="00:00:58.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="501" swimtime="00:19:03.00" resultid="1462" heatid="1929" lane="3" />
                <RESULT eventid="1302" points="493" swimtime="00:00:29.02" resultid="1463" heatid="1994" lane="3" entrytime="00:00:27.92" entrycourse="SCM" />
                <RESULT eventid="1270" points="468" swimtime="00:01:10.68" resultid="1464" heatid="1979" lane="3" entrytime="00:01:05.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="492" swimtime="00:04:52.80" resultid="1465" heatid="1956" lane="4" entrytime="00:04:37.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                    <SPLIT distance="100" swimtime="00:01:09.86" />
                    <SPLIT distance="150" swimtime="00:01:46.94" />
                    <SPLIT distance="200" swimtime="00:02:23.79" />
                    <SPLIT distance="250" swimtime="00:03:00.22" />
                    <SPLIT distance="300" swimtime="00:03:36.85" />
                    <SPLIT distance="350" swimtime="00:04:14.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Resende Ames" birthdate="2010-02-02" gender="M" nation="BRA" license="365505" swrid="5588876" athleteid="1537" externalid="365505" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1168" points="279" swimtime="00:01:13.05" resultid="1538" heatid="1942" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="364" swimtime="00:01:02.80" resultid="1539" heatid="1922" lane="5" entrytime="00:01:04.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="306" swimtime="00:00:29.90" resultid="1540" heatid="1997" lane="1" entrytime="00:00:29.54" entrycourse="SCM" />
                <RESULT eventid="1278" points="355" swimtime="00:01:08.23" resultid="1541" heatid="1982" lane="3" entrytime="00:01:06.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="385" swimtime="00:04:51.55" resultid="1542" heatid="1951" lane="6" entrytime="00:04:47.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                    <SPLIT distance="100" swimtime="00:01:08.43" />
                    <SPLIT distance="150" swimtime="00:01:45.25" />
                    <SPLIT distance="200" swimtime="00:02:21.69" />
                    <SPLIT distance="250" swimtime="00:02:59.56" />
                    <SPLIT distance="300" swimtime="00:03:37.54" />
                    <SPLIT distance="350" swimtime="00:04:14.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jeronimo" lastname="Pujato Flores" birthdate="2013-12-28" gender="M" nation="BRA" license="392839" swrid="5652625" athleteid="1618" externalid="392839" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1151" points="66" swimtime="00:00:54.71" resultid="1619" heatid="1937" lane="1" entrytime="00:00:52.42" entrycourse="SCM" />
                <RESULT eventid="1079" status="DSQ" swimtime="00:02:12.52" resultid="1620" heatid="1913" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="108" swimtime="00:00:42.33" resultid="1621" heatid="1990" lane="2" entrytime="00:00:46.49" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Bailke" birthdate="2007-05-04" gender="M" nation="BRA" license="370566" swrid="5596869" athleteid="1496" externalid="370566" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1168" points="267" swimtime="00:01:14.15" resultid="1497" heatid="1943" lane="4" entrytime="00:01:12.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="333" swimtime="00:20:20.71" resultid="1498" heatid="1931" lane="2" />
                <RESULT eventid="1310" points="314" swimtime="00:00:29.65" resultid="1499" heatid="1997" lane="6" entrytime="00:00:29.62" entrycourse="SCM" />
                <RESULT eventid="1252" points="286" swimtime="00:00:33.00" resultid="1500" heatid="1971" lane="2" />
                <RESULT eventid="1192" points="376" swimtime="00:04:54.06" resultid="1501" heatid="1950" lane="3" entrytime="00:04:50.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                    <SPLIT distance="100" swimtime="00:01:12.87" />
                    <SPLIT distance="150" swimtime="00:01:49.89" />
                    <SPLIT distance="200" swimtime="00:02:28.06" />
                    <SPLIT distance="250" swimtime="00:03:04.89" />
                    <SPLIT distance="300" swimtime="00:03:42.20" />
                    <SPLIT distance="350" swimtime="00:04:18.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mayumi" lastname="Napole" birthdate="2010-02-01" gender="F" nation="BRA" license="376446" swrid="5596918" athleteid="1556" externalid="376446" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1088" points="360" swimtime="00:01:10.60" resultid="1557" heatid="1919" lane="6" entrytime="00:01:08.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="306" swimtime="00:03:00.66" resultid="1558" heatid="1905" lane="5" entrytime="00:02:55.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.20" />
                    <SPLIT distance="100" swimtime="00:01:27.35" />
                    <SPLIT distance="150" swimtime="00:02:19.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="380" swimtime="00:00:31.64" resultid="1559" heatid="1994" lane="5" entrytime="00:00:31.09" entrycourse="SCM" />
                <RESULT eventid="1270" points="311" swimtime="00:01:20.97" resultid="1560" heatid="1979" lane="1" entrytime="00:01:18.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="314" swimtime="00:05:40.18" resultid="1561" heatid="1953" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                    <SPLIT distance="100" swimtime="00:01:21.28" />
                    <SPLIT distance="150" swimtime="00:02:05.52" />
                    <SPLIT distance="200" swimtime="00:02:49.60" />
                    <SPLIT distance="250" swimtime="00:03:33.24" />
                    <SPLIT distance="300" swimtime="00:04:16.59" />
                    <SPLIT distance="350" swimtime="00:04:59.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Luiz Martinazzo" birthdate="2006-05-16" gender="M" nation="BRA" license="345593" swrid="5596910" athleteid="1484" externalid="345593" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1068" points="426" swimtime="00:02:25.62" resultid="1485" heatid="1910" lane="4" entrytime="00:02:25.66" entrycourse="SCM" />
                <RESULT eventid="1124" points="455" swimtime="00:18:20.40" resultid="1486" heatid="1932" lane="4" entrytime="00:17:57.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:18:20.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="448" swimtime="00:00:26.34" resultid="1487" heatid="1995" lane="5" />
                <RESULT eventid="1278" points="399" swimtime="00:01:05.60" resultid="1488" heatid="1983" lane="5" entrytime="00:01:03.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="453" swimtime="00:04:36.21" resultid="1489" heatid="1952" lane="1" entrytime="00:04:25.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                    <SPLIT distance="100" swimtime="00:01:04.05" />
                    <SPLIT distance="150" swimtime="00:01:39.16" />
                    <SPLIT distance="200" swimtime="00:02:13.93" />
                    <SPLIT distance="250" swimtime="00:02:49.21" />
                    <SPLIT distance="300" swimtime="00:03:25.10" />
                    <SPLIT distance="350" swimtime="00:04:00.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Ioris Souza" birthdate="2015-09-10" gender="F" nation="BRA" license="406693" athleteid="1622" externalid="406693" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1154" points="54" swimtime="00:01:06.75" resultid="1623" heatid="1938" lane="6" />
                <RESULT eventid="1082" points="59" swimtime="00:01:12.58" resultid="1624" heatid="1914" lane="4" />
                <RESULT eventid="1290" points="54" swimtime="00:01:00.61" resultid="1625" heatid="1986" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Carvalho Carelli" birthdate="2011-10-15" gender="M" nation="BRA" license="403146" swrid="5676300" athleteid="1588" externalid="403146" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1168" points="150" swimtime="00:01:29.91" resultid="1589" heatid="1943" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="220" swimtime="00:01:14.21" resultid="1590" heatid="1921" lane="6" entrytime="00:01:27.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="215" swimtime="00:00:33.63" resultid="1591" heatid="1996" lane="1" entrytime="00:00:34.88" entrycourse="SCM" />
                <RESULT eventid="1252" points="196" swimtime="00:00:37.38" resultid="1592" heatid="1972" lane="1" entrytime="00:00:41.65" entrycourse="SCM" />
                <RESULT eventid="1192" points="202" swimtime="00:06:01.31" resultid="1593" heatid="1948" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:23.63" />
                    <SPLIT distance="150" swimtime="00:02:10.91" />
                    <SPLIT distance="200" swimtime="00:02:56.87" />
                    <SPLIT distance="250" swimtime="00:03:43.54" />
                    <SPLIT distance="300" swimtime="00:04:27.90" />
                    <SPLIT distance="350" swimtime="00:05:07.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marlon" lastname="Antonio Junior" birthdate="2013-05-12" gender="M" nation="BRA" license="397300" swrid="5641751" athleteid="1573" externalid="397300" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1107" points="139" swimtime="00:03:11.82" resultid="1574" heatid="1925" lane="2" entrytime="00:03:21.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                    <SPLIT distance="100" swimtime="00:01:31.85" />
                    <SPLIT distance="150" swimtime="00:02:24.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="103" swimtime="00:01:57.64" resultid="1575" heatid="1913" lane="1" />
                <RESULT eventid="1299" points="131" swimtime="00:00:39.60" resultid="1576" heatid="1991" lane="6" entrytime="00:00:38.85" entrycourse="SCM" />
                <RESULT eventid="1267" status="DSQ" swimtime="00:01:38.15" resultid="1577" heatid="1975" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Paulo Sales" birthdate="2007-11-07" gender="M" nation="BRA" license="390712" swrid="5596923" athleteid="1514" externalid="390712" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1096" points="283" swimtime="00:01:08.29" resultid="1515" heatid="1921" lane="3" entrytime="00:01:08.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="266" swimtime="00:02:50.31" resultid="1516" heatid="1907" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                    <SPLIT distance="100" swimtime="00:01:19.53" />
                    <SPLIT distance="150" swimtime="00:02:09.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="301" swimtime="00:00:30.08" resultid="1517" heatid="1996" lane="2" entrytime="00:00:31.01" entrycourse="SCM" />
                <RESULT eventid="1236" points="246" swimtime="00:01:28.19" resultid="1518" heatid="1968" lane="6" entrytime="00:01:28.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="282" swimtime="00:05:23.38" resultid="1519" heatid="1947" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                    <SPLIT distance="100" swimtime="00:01:11.67" />
                    <SPLIT distance="150" swimtime="00:01:52.97" />
                    <SPLIT distance="200" swimtime="00:02:35.23" />
                    <SPLIT distance="250" swimtime="00:03:17.84" />
                    <SPLIT distance="300" swimtime="00:04:00.79" />
                    <SPLIT distance="350" swimtime="00:04:43.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edward" lastname="Mikael De Lima" birthdate="2012-03-11" gender="M" nation="BRA" license="376445" swrid="5588816" athleteid="1551" externalid="376445" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1151" points="251" swimtime="00:00:35.03" resultid="1552" heatid="1936" lane="4" />
                <RESULT eventid="1107" points="324" swimtime="00:02:24.63" resultid="1553" heatid="1926" lane="3" entrytime="00:02:25.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:08.86" />
                    <SPLIT distance="150" swimtime="00:01:46.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="309" swimtime="00:00:29.80" resultid="1554" heatid="1991" lane="3" entrytime="00:00:30.23" entrycourse="SCM" />
                <RESULT eventid="1221" points="222" swimtime="00:01:18.84" resultid="1555" heatid="1962" lane="3" entrytime="00:01:22.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katherine" lastname="Kotz" birthdate="2012-05-18" gender="F" nation="BRA" license="390810" swrid="5596907" athleteid="1532" externalid="390810" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1104" points="238" swimtime="00:02:57.84" resultid="1533" heatid="1924" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                    <SPLIT distance="100" swimtime="00:01:29.11" />
                    <SPLIT distance="150" swimtime="00:02:16.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1076" points="222" swimtime="00:01:42.93" resultid="1534" heatid="1912" lane="3" entrytime="00:01:48.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="316" swimtime="00:00:33.66" resultid="1535" heatid="1989" lane="3" entrytime="00:00:33.71" entrycourse="SCM" />
                <RESULT eventid="1264" points="230" swimtime="00:01:32.10" resultid="1536" heatid="1974" lane="2" entrytime="00:01:50.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Mattiello" birthdate="2009-04-11" gender="F" nation="BRA" license="367011" swrid="5596914" athleteid="1502" externalid="367011" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1088" points="392" swimtime="00:01:08.62" resultid="1503" heatid="1918" lane="3" entrytime="00:01:08.32" entrycourse="SCM" />
                <RESULT eventid="1116" points="317" swimtime="00:22:11.43" resultid="1504" heatid="1929" lane="4" />
                <RESULT eventid="1302" points="365" swimtime="00:00:32.06" resultid="1505" heatid="1994" lane="1" entrytime="00:00:31.16" entrycourse="SCM" />
                <RESULT eventid="1270" points="290" swimtime="00:01:22.88" resultid="1506" heatid="1978" lane="2" entrytime="00:01:21.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="373" swimtime="00:05:21.10" resultid="1507" heatid="1955" lane="4" entrytime="00:05:14.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                    <SPLIT distance="100" swimtime="00:01:17.87" />
                    <SPLIT distance="150" swimtime="00:01:24.63" />
                    <SPLIT distance="200" swimtime="00:01:58.36" />
                    <SPLIT distance="250" swimtime="00:02:39.67" />
                    <SPLIT distance="300" swimtime="00:03:21.17" />
                    <SPLIT distance="350" swimtime="00:04:02.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Faisal" lastname="Basem Ghotme" birthdate="2010-12-18" gender="M" nation="BRA" license="390809" swrid="5596871" athleteid="1567" externalid="390809" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1096" points="344" swimtime="00:01:03.96" resultid="1568" heatid="1922" lane="2" entrytime="00:01:03.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="324" swimtime="00:02:39.51" resultid="1569" heatid="1909" lane="5" entrytime="00:02:47.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:14.75" />
                    <SPLIT distance="150" swimtime="00:02:05.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="387" swimtime="00:00:27.65" resultid="1570" heatid="1997" lane="2" entrytime="00:00:27.96" entrycourse="SCM" />
                <RESULT eventid="1278" points="335" swimtime="00:01:09.56" resultid="1571" heatid="1982" lane="1" entrytime="00:01:08.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="282" swimtime="00:05:23.58" resultid="1572" heatid="1948" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="100" swimtime="00:01:15.13" />
                    <SPLIT distance="150" swimtime="00:01:57.30" />
                    <SPLIT distance="200" swimtime="00:02:39.61" />
                    <SPLIT distance="250" swimtime="00:03:23.30" />
                    <SPLIT distance="300" swimtime="00:04:05.13" />
                    <SPLIT distance="350" swimtime="00:04:46.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Omar" lastname="Pinheiro" birthdate="1981-09-04" gender="M" nation="BRA" license="305962" swrid="5596926" athleteid="1451" externalid="305962" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1310" points="472" swimtime="00:00:25.88" resultid="1452" heatid="1998" lane="2" entrytime="00:00:25.15" entrycourse="SCM" />
                <RESULT eventid="1278" points="328" swimtime="00:01:10.04" resultid="1453" heatid="1980" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Abraao" lastname="Felipe Oliveira" birthdate="2012-05-20" gender="M" nation="BRA" license="400457" swrid="5420917" athleteid="1583" externalid="400457" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1151" points="65" swimtime="00:00:54.84" resultid="1584" heatid="1936" lane="3" entrytime="00:00:57.16" entrycourse="SCM" />
                <RESULT eventid="1107" points="115" swimtime="00:03:24.29" resultid="1585" heatid="1925" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.48" />
                    <SPLIT distance="100" swimtime="00:01:36.35" />
                    <SPLIT distance="150" swimtime="00:02:30.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="133" swimtime="00:00:39.46" resultid="1586" heatid="1990" lane="3" entrytime="00:00:39.13" entrycourse="SCM" />
                <RESULT eventid="1267" status="DSQ" swimtime="00:01:45.09" resultid="1587" heatid="1975" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Kasprzak" birthdate="2011-08-09" gender="F" nation="BRA" license="406659" athleteid="1613" externalid="406659" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1176" points="105" swimtime="00:01:00.08" resultid="1614" heatid="1945" lane="4" />
                <RESULT eventid="1088" status="DSQ" swimtime="00:01:54.57" resultid="1615" heatid="1917" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="69" swimtime="00:00:55.65" resultid="1616" heatid="1992" lane="2" />
                <RESULT eventid="1228" status="DSQ" swimtime="00:02:11.53" resultid="1617" heatid="1965" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Carolina Ghellere" birthdate="2007-06-05" gender="F" nation="BRA" license="312662" swrid="5596874" athleteid="1445" externalid="312662" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1160" points="471" swimtime="00:01:09.45" resultid="1446" heatid="1941" lane="3" entrytime="00:01:05.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="486" swimtime="00:02:34.97" resultid="1447" heatid="1906" lane="3" entrytime="00:02:32.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                    <SPLIT distance="100" swimtime="00:01:13.23" />
                    <SPLIT distance="150" swimtime="00:01:59.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="451" swimtime="00:00:29.89" resultid="1448" heatid="1992" lane="4" />
                <RESULT eventid="1244" points="429" swimtime="00:00:32.32" resultid="1449" heatid="1970" lane="3" entrytime="00:00:30.19" entrycourse="SCM" />
                <RESULT eventid="1200" points="501" swimtime="00:04:51.19" resultid="1450" heatid="1956" lane="3" entrytime="00:04:27.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                    <SPLIT distance="100" swimtime="00:01:09.73" />
                    <SPLIT distance="150" swimtime="00:01:46.77" />
                    <SPLIT distance="200" swimtime="00:02:23.73" />
                    <SPLIT distance="250" swimtime="00:02:59.63" />
                    <SPLIT distance="300" swimtime="00:03:36.66" />
                    <SPLIT distance="350" swimtime="00:04:14.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Targat Pinheiro" birthdate="2008-09-04" gender="F" nation="BRA" license="331610" swrid="5596894" athleteid="1434" externalid="331610" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1160" points="422" swimtime="00:01:12.03" resultid="1435" heatid="1941" lane="2" entrytime="00:01:12.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="411" swimtime="00:02:43.78" resultid="1436" heatid="1906" lane="5" entrytime="00:02:38.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:14.45" />
                    <SPLIT distance="150" swimtime="00:02:04.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="431" swimtime="00:20:01.76" resultid="1437" heatid="1930" lane="3" entrytime="00:19:51.15" entrycourse="SCM" />
                <RESULT eventid="1270" points="349" swimtime="00:01:17.94" resultid="1438" heatid="1979" lane="2" entrytime="00:01:15.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="424" swimtime="00:05:07.70" resultid="1439" heatid="1956" lane="5" entrytime="00:04:57.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:11.99" />
                    <SPLIT distance="150" swimtime="00:01:51.12" />
                    <SPLIT distance="200" swimtime="00:02:30.32" />
                    <SPLIT distance="250" swimtime="00:03:09.72" />
                    <SPLIT distance="300" swimtime="00:03:50.09" />
                    <SPLIT distance="350" swimtime="00:04:29.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Gabriel Dreher" birthdate="2011-12-05" gender="M" nation="BRA" license="403148" swrid="5676302" athleteid="1599" externalid="403148" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1184" points="84" swimtime="00:00:56.95" resultid="1600" heatid="1946" lane="6" />
                <RESULT eventid="1140" points="98" swimtime="00:00:47.84" resultid="1601" heatid="1934" lane="4" />
                <RESULT eventid="1096" points="101" swimtime="00:01:35.97" resultid="1602" heatid="1920" lane="3" entrytime="00:01:47.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" status="DNS" swimtime="00:00:00.00" resultid="1603" heatid="1995" lane="2" entrytime="00:00:43.48" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Resende Ames" birthdate="2006-02-10" gender="M" nation="BRA" license="365657" swrid="5596931" athleteid="1472" externalid="365657" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1096" points="538" swimtime="00:00:55.10" resultid="1473" heatid="1923" lane="4" entrytime="00:00:54.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" status="DSQ" swimtime="00:00:00.00" resultid="1474" heatid="1908" lane="1" />
                <RESULT eventid="1310" points="494" swimtime="00:00:25.49" resultid="1475" heatid="1998" lane="5" entrytime="00:00:25.94" entrycourse="SCM" />
                <RESULT eventid="1278" points="400" swimtime="00:01:05.59" resultid="1476" heatid="1982" lane="4" entrytime="00:01:07.09" entrycourse="SCM" />
                <RESULT eventid="1192" points="564" swimtime="00:04:16.79" resultid="1477" heatid="1952" lane="4" entrytime="00:04:16.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.90" />
                    <SPLIT distance="100" swimtime="00:01:01.16" />
                    <SPLIT distance="150" swimtime="00:01:33.57" />
                    <SPLIT distance="200" swimtime="00:02:05.77" />
                    <SPLIT distance="250" swimtime="00:02:37.85" />
                    <SPLIT distance="300" swimtime="00:03:10.50" />
                    <SPLIT distance="350" swimtime="00:03:43.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaleo" lastname="Bruno Da Luz" birthdate="2014-03-11" gender="M" nation="BRA" license="406658" athleteid="1610" externalid="406658" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1157" points="22" swimtime="00:01:18.70" resultid="1611" heatid="1939" lane="2" />
                <RESULT eventid="1293" points="26" swimtime="00:01:07.30" resultid="1612" heatid="1988" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Oliveira" birthdate="2003-07-16" gender="M" nation="BRA" license="295723" swrid="5596944" athleteid="1466" externalid="295723" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1168" points="469" swimtime="00:01:01.49" resultid="1467" heatid="1944" lane="4" entrytime="00:00:59.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="470" swimtime="00:00:57.65" resultid="1468" heatid="1920" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="415" swimtime="00:01:04.77" resultid="1469" heatid="1983" lane="4" entrytime="00:01:00.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="506" swimtime="00:00:27.29" resultid="1470" heatid="1972" lane="3" entrytime="00:00:26.34" entrycourse="SCM" />
                <RESULT eventid="1192" points="460" swimtime="00:04:34.79" resultid="1471" heatid="1947" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.49" />
                    <SPLIT distance="100" swimtime="00:01:06.51" />
                    <SPLIT distance="150" swimtime="00:01:41.40" />
                    <SPLIT distance="200" swimtime="00:02:16.11" />
                    <SPLIT distance="250" swimtime="00:02:51.05" />
                    <SPLIT distance="300" swimtime="00:03:26.00" />
                    <SPLIT distance="350" swimtime="00:04:00.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Rogge" birthdate="2008-09-02" gender="M" nation="BRA" license="383387" swrid="4883279" athleteid="1454" externalid="383387" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1096" points="428" swimtime="00:00:59.50" resultid="1455" heatid="1923" lane="1" entrytime="00:00:58.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="307" swimtime="00:02:42.36" resultid="1456" heatid="1908" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:10.98" />
                    <SPLIT distance="150" swimtime="00:02:02.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="450" swimtime="00:00:26.29" resultid="1457" heatid="1998" lane="1" entrytime="00:00:26.54" entrycourse="SCM" />
                <RESULT eventid="1278" points="331" swimtime="00:01:09.80" resultid="1458" heatid="1982" lane="2" entrytime="00:01:07.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="259" swimtime="00:05:32.59" resultid="1459" heatid="1948" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:15.37" />
                    <SPLIT distance="150" swimtime="00:01:56.83" />
                    <SPLIT distance="200" swimtime="00:02:39.69" />
                    <SPLIT distance="250" swimtime="00:03:23.09" />
                    <SPLIT distance="300" swimtime="00:04:06.42" />
                    <SPLIT distance="350" swimtime="00:04:48.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="NATION" code="729" nation="PAR" clubid="1897" name="Seleção do Paraguai" shortname="Paraguai">
          <ATHLETES>
            <ATHLETE firstname="Cristhiane" lastname="Añasco Kliemann" birthdate="2009-02-03" gender="F" nation="PAR" license="V381201" swrid="5654088" athleteid="1898" externalid="V381201">
              <RESULTS>
                <RESULT eventid="1160" points="362" status="EXH" swimtime="00:01:15.82" resultid="1899" heatid="1940" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="550" status="EXH" swimtime="00:00:30.80" resultid="1900" heatid="1933" lane="5" />
                <RESULT eventid="1060" points="453" status="EXH" swimtime="00:02:38.67" resultid="1901" heatid="1904" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:12.09" />
                    <SPLIT distance="150" swimtime="00:02:00.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="504" status="EXH" swimtime="00:01:08.93" resultid="1902" heatid="1977" lane="2" />
                <RESULT eventid="1244" points="483" status="EXH" swimtime="00:00:31.07" resultid="1903" heatid="1970" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="572" nation="BRA" region="RS" clubid="1427" swrid="93767" name="Associação Serrana De Desportos Aquáticos" shortname="Asda">
          <ATHLETES>
            <ATHLETE firstname="Francieli" lastname="Añasco" birthdate="2014-05-27" gender="F" nation="PRY" license="394219" athleteid="1428" externalid="394219">
              <RESULTS>
                <RESULT eventid="1110" points="223" status="EXH" swimtime="00:01:22.83" resultid="1429" heatid="1927" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1082" points="165" status="EXH" swimtime="00:00:51.72" resultid="1430" heatid="1914" lane="5" />
                <RESULT eventid="1290" points="220" status="EXH" swimtime="00:00:37.97" resultid="1431" heatid="1987" lane="3" entrytime="00:00:39.37" entrycourse="SCM" />
                <RESULT eventid="1212" points="180" status="EXH" swimtime="00:00:43.15" resultid="1432" heatid="1957" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="36" nation="BRA" region="PR" clubid="1630" swrid="93753" name="Associação Atlética Comercial" shortname="Comercial Cascavel">
          <ATHLETES>
            <ATHLETE firstname="Helena" lastname="Queiroz Da Costa" birthdate="2014-05-30" gender="F" nation="BRA" license="406698" athleteid="1892" externalid="406698">
              <RESULTS>
                <RESULT eventid="1110" points="90" swimtime="00:01:51.76" resultid="1893" heatid="1927" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1082" points="87" swimtime="00:01:03.99" resultid="1894" heatid="1914" lane="3" />
                <RESULT eventid="1290" points="114" swimtime="00:00:47.22" resultid="1895" heatid="1986" lane="6" />
                <RESULT eventid="1212" points="59" swimtime="00:01:02.51" resultid="1896" heatid="1957" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Emanuel Rech" birthdate="2013-12-02" gender="M" nation="BRA" license="380660" swrid="5588679" athleteid="1750" externalid="380660">
              <RESULTS>
                <RESULT eventid="1107" points="205" swimtime="00:02:48.46" resultid="1751" heatid="1926" lane="6" entrytime="00:02:55.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                    <SPLIT distance="100" swimtime="00:01:21.56" />
                    <SPLIT distance="150" swimtime="00:02:06.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="158" swimtime="00:01:42.19" resultid="1752" heatid="1913" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="172" swimtime="00:01:28.51" resultid="1753" heatid="1976" lane="4" entrytime="00:01:32.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1221" points="100" swimtime="00:01:42.76" resultid="1754" heatid="1961" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Alves Serafini" birthdate="2008-04-15" gender="M" nation="BRA" license="351644" swrid="5596867" athleteid="1792" externalid="351644">
              <RESULTS>
                <RESULT eventid="1168" points="458" swimtime="00:01:01.96" resultid="1793" heatid="1944" lane="5" entrytime="00:01:03.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="463" swimtime="00:00:57.95" resultid="1794" heatid="1923" lane="6" entrytime="00:00:58.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="420" swimtime="00:02:26.34" resultid="1795" heatid="1910" lane="3" entrytime="00:02:25.56" entrycourse="SCM" />
                <RESULT eventid="1310" points="419" swimtime="00:00:26.93" resultid="1796" heatid="1997" lane="3" entrytime="00:00:27.17" entrycourse="SCM" />
                <RESULT eventid="1192" points="478" swimtime="00:04:31.43" resultid="1797" heatid="1951" lane="4" entrytime="00:04:32.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:05.13" />
                    <SPLIT distance="150" swimtime="00:01:39.47" />
                    <SPLIT distance="200" swimtime="00:02:13.66" />
                    <SPLIT distance="250" swimtime="00:02:47.79" />
                    <SPLIT distance="300" swimtime="00:03:22.19" />
                    <SPLIT distance="350" swimtime="00:03:56.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Vieira Rohnelt" birthdate="2012-05-03" gender="M" nation="BRA" license="365692" swrid="5588952" athleteid="1697" externalid="365692">
              <RESULTS>
                <RESULT eventid="1107" status="WDR" swimtime="00:00:00.00" resultid="1698" heatid="1926" lane="1" entrytime="00:02:51.71" entrycourse="SCM" />
                <RESULT eventid="1079" status="DNS" swimtime="00:00:00.00" resultid="1699" heatid="1913" lane="3" entrytime="00:01:45.30" entrycourse="SCM" />
                <RESULT eventid="1267" status="WDR" swimtime="00:00:00.00" resultid="1700" heatid="1975" lane="2" />
                <RESULT eventid="1221" status="WDR" swimtime="00:00:00.00" resultid="1701" heatid="1962" lane="4" entrytime="00:01:43.15" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Luiza Bezerra Sedlacek" birthdate="2008-04-18" gender="F" nation="BRA" license="344607" swrid="4496478" athleteid="1655" externalid="344607">
              <RESULTS>
                <RESULT eventid="1088" points="485" swimtime="00:01:03.93" resultid="1656" heatid="1919" lane="4" entrytime="00:01:02.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="458" swimtime="00:02:38.04" resultid="1657" heatid="1906" lane="2" entrytime="00:02:36.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                    <SPLIT distance="100" swimtime="00:01:14.24" />
                    <SPLIT distance="150" swimtime="00:02:01.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="447" swimtime="00:00:29.98" resultid="1658" heatid="1992" lane="3" />
                <RESULT eventid="1270" points="404" swimtime="00:01:14.19" resultid="1659" heatid="1977" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="461" swimtime="00:04:59.27" resultid="1660" heatid="1956" lane="2" entrytime="00:04:47.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:10.69" />
                    <SPLIT distance="150" swimtime="00:01:48.18" />
                    <SPLIT distance="200" swimtime="00:02:26.30" />
                    <SPLIT distance="250" swimtime="00:03:04.59" />
                    <SPLIT distance="300" swimtime="00:03:43.13" />
                    <SPLIT distance="350" swimtime="00:04:21.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luann" lastname="Miguel Mazur" birthdate="2007-01-10" gender="M" nation="BRA" license="365682" swrid="5596915" athleteid="1685" externalid="365682">
              <RESULTS>
                <RESULT eventid="1168" points="327" swimtime="00:01:09.31" resultid="1686" heatid="1942" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="453" swimtime="00:02:22.72" resultid="1687" heatid="1911" lane="2" entrytime="00:02:21.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                    <SPLIT distance="100" swimtime="00:01:08.79" />
                    <SPLIT distance="150" swimtime="00:01:49.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="320" swimtime="00:01:10.60" resultid="1688" heatid="1981" lane="3" entrytime="00:01:11.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="414" swimtime="00:01:14.15" resultid="1689" heatid="1969" lane="5" entrytime="00:01:13.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="453" swimtime="00:04:36.18" resultid="1690" heatid="1951" lane="5" entrytime="00:04:41.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:01:07.03" />
                    <SPLIT distance="150" swimtime="00:01:42.09" />
                    <SPLIT distance="200" swimtime="00:02:17.69" />
                    <SPLIT distance="250" swimtime="00:02:54.12" />
                    <SPLIT distance="300" swimtime="00:03:29.88" />
                    <SPLIT distance="350" swimtime="00:04:02.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Flavia" lastname="De Metz" birthdate="2011-01-07" gender="F" nation="BRA" license="390846" swrid="5596887" athleteid="1839" externalid="390846">
              <RESULTS>
                <RESULT eventid="1160" points="172" swimtime="00:01:37.16" resultid="1840" heatid="1940" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="292" swimtime="00:03:03.54" resultid="1841" heatid="1904" lane="3" entrytime="00:03:04.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.86" />
                    <SPLIT distance="100" swimtime="00:01:29.66" />
                    <SPLIT distance="150" swimtime="00:02:22.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="257" swimtime="00:01:26.30" resultid="1842" heatid="1978" lane="6" entrytime="00:01:23.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="247" swimtime="00:01:39.33" resultid="1843" heatid="1966" lane="6" entrytime="00:01:42.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="361" swimtime="00:05:24.62" resultid="1844" heatid="1955" lane="1" entrytime="00:05:27.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:01:18.76" />
                    <SPLIT distance="150" swimtime="00:01:59.86" />
                    <SPLIT distance="200" swimtime="00:02:41.85" />
                    <SPLIT distance="250" swimtime="00:03:23.07" />
                    <SPLIT distance="300" swimtime="00:04:03.22" />
                    <SPLIT distance="350" swimtime="00:04:44.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marianna" lastname="Galvao Oliveira" birthdate="2014-03-18" gender="F" nation="BRA" license="390835" swrid="5596902" athleteid="1808" externalid="390835">
              <RESULTS>
                <RESULT eventid="1154" points="109" swimtime="00:00:52.74" resultid="1809" heatid="1938" lane="5" entrytime="00:00:54.87" entrycourse="SCM" />
                <RESULT eventid="1082" points="189" swimtime="00:00:49.35" resultid="1810" heatid="1915" lane="4" entrytime="00:00:55.67" entrycourse="SCM" />
                <RESULT eventid="1290" points="145" swimtime="00:00:43.63" resultid="1811" heatid="1987" lane="1" entrytime="00:00:45.28" entrycourse="SCM" />
                <RESULT eventid="1212" points="99" swimtime="00:00:52.68" resultid="1812" heatid="1958" lane="2" entrytime="00:00:54.28" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ramirez Vasconcelos" birthdate="2011-04-06" gender="M" nation="BRA" license="392013" swrid="4863662" athleteid="1850" externalid="392013">
              <RESULTS>
                <RESULT eventid="1096" points="220" swimtime="00:01:14.25" resultid="1851" heatid="1921" lane="1" entrytime="00:01:18.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="223" swimtime="00:03:00.67" resultid="1852" heatid="1908" lane="3" entrytime="00:02:55.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                    <SPLIT distance="100" swimtime="00:01:24.10" />
                    <SPLIT distance="150" swimtime="00:02:18.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="185" swimtime="00:01:24.81" resultid="1853" heatid="1980" lane="2" entrytime="00:02:01.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="237" swimtime="00:01:29.29" resultid="1854" heatid="1967" lane="5" entrytime="00:01:43.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="280" swimtime="00:05:24.10" resultid="1855" heatid="1949" lane="1" entrytime="00:06:42.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:17.30" />
                    <SPLIT distance="150" swimtime="00:01:59.24" />
                    <SPLIT distance="200" swimtime="00:02:41.32" />
                    <SPLIT distance="250" swimtime="00:03:23.42" />
                    <SPLIT distance="300" swimtime="00:04:03.92" />
                    <SPLIT distance="350" swimtime="00:04:45.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jordana" lastname="Rinaldini" birthdate="2004-09-13" gender="F" nation="BRA" license="342426" swrid="5596933" athleteid="1643" externalid="342426">
              <RESULTS>
                <RESULT eventid="1088" points="336" swimtime="00:01:12.26" resultid="1644" heatid="1918" lane="4" entrytime="00:01:09.42" entrycourse="SCM" />
                <RESULT eventid="1060" points="351" swimtime="00:02:52.71" resultid="1645" heatid="1906" lane="6" entrytime="00:02:47.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                    <SPLIT distance="100" swimtime="00:01:20.09" />
                    <SPLIT distance="150" swimtime="00:02:10.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="339" swimtime="00:00:32.86" resultid="1646" heatid="1993" lane="5" />
                <RESULT eventid="1270" points="318" swimtime="00:01:20.41" resultid="1647" heatid="1979" lane="5" entrytime="00:01:17.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="351" swimtime="00:05:27.66" resultid="1648" heatid="1955" lane="2" entrytime="00:05:19.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:17.60" />
                    <SPLIT distance="150" swimtime="00:01:59.23" />
                    <SPLIT distance="200" swimtime="00:02:40.93" />
                    <SPLIT distance="250" swimtime="00:03:22.95" />
                    <SPLIT distance="300" swimtime="00:04:05.19" />
                    <SPLIT distance="350" swimtime="00:04:47.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Claudio" lastname="Rohnelt" birthdate="2010-03-08" gender="M" nation="BRA" license="357954" swrid="5596935" athleteid="1679" externalid="357954">
              <RESULTS>
                <RESULT eventid="1168" points="218" swimtime="00:01:19.28" resultid="1680" heatid="1943" lane="5" entrytime="00:01:17.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="249" swimtime="00:02:54.03" resultid="1681" heatid="1909" lane="6" entrytime="00:02:51.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:22.61" />
                    <SPLIT distance="150" swimtime="00:02:13.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="193" swimtime="00:01:23.50" resultid="1682" heatid="1980" lane="4" entrytime="00:01:23.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="217" swimtime="00:00:36.19" resultid="1683" heatid="1972" lane="5" entrytime="00:00:35.78" entrycourse="SCM" />
                <RESULT eventid="1192" points="303" swimtime="00:05:15.75" resultid="1684" heatid="1949" lane="2" entrytime="00:05:23.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                    <SPLIT distance="100" swimtime="00:01:14.37" />
                    <SPLIT distance="150" swimtime="00:01:53.88" />
                    <SPLIT distance="200" swimtime="00:02:34.28" />
                    <SPLIT distance="250" swimtime="00:03:14.97" />
                    <SPLIT distance="300" swimtime="00:03:55.64" />
                    <SPLIT distance="350" swimtime="00:04:36.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Gaio" birthdate="2014-08-27" gender="F" nation="BRA" license="390841" swrid="5596900" athleteid="1824" externalid="390841">
              <RESULTS>
                <RESULT eventid="1154" points="97" swimtime="00:00:54.79" resultid="1825" heatid="1938" lane="1" entrytime="00:01:02.63" entrycourse="SCM" />
                <RESULT eventid="1082" points="130" swimtime="00:00:56.00" resultid="1826" heatid="1915" lane="1" entrytime="00:01:01.45" entrycourse="SCM" />
                <RESULT eventid="1290" points="136" swimtime="00:00:44.58" resultid="1827" heatid="1986" lane="4" entrytime="00:00:48.27" entrycourse="SCM" />
                <RESULT eventid="1212" points="81" swimtime="00:00:56.30" resultid="1828" heatid="1957" lane="3" entrytime="00:01:25.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Henrique Marca Dos Santos" birthdate="2015-03-28" gender="M" nation="BRA" license="406695" athleteid="1878" externalid="406695">
              <RESULTS>
                <RESULT eventid="1157" points="49" swimtime="00:01:00.14" resultid="1879" heatid="1939" lane="3" />
                <RESULT eventid="1113" points="49" swimtime="00:02:02.34" resultid="1880" heatid="1928" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="51" swimtime="00:01:07.12" resultid="1881" heatid="1916" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Sehn Uren" birthdate="2009-10-15" gender="F" nation="BRA" license="357159" swrid="5596937" athleteid="1667" externalid="357159">
              <RESULTS>
                <RESULT eventid="1088" points="369" swimtime="00:01:10.03" resultid="1668" heatid="1917" lane="3" entrytime="00:01:19.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="388" swimtime="00:02:47.06" resultid="1669" heatid="1905" lane="3" entrytime="00:02:49.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:01:21.66" />
                    <SPLIT distance="150" swimtime="00:02:08.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="304" swimtime="00:01:21.58" resultid="1670" heatid="1978" lane="4" entrytime="00:01:20.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="338" swimtime="00:01:29.50" resultid="1671" heatid="1965" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="326" swimtime="00:05:35.98" resultid="1672" heatid="1954" lane="4" entrytime="00:05:41.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                    <SPLIT distance="100" swimtime="00:01:20.96" />
                    <SPLIT distance="150" swimtime="00:02:03.51" />
                    <SPLIT distance="200" swimtime="00:02:47.23" />
                    <SPLIT distance="250" swimtime="00:03:29.38" />
                    <SPLIT distance="300" swimtime="00:04:12.22" />
                    <SPLIT distance="350" swimtime="00:04:55.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Bertelli Weirich" birthdate="2011-03-18" gender="F" nation="BRA" license="369534" swrid="5588552" athleteid="1714" externalid="369534">
              <RESULTS>
                <RESULT eventid="1160" points="264" swimtime="00:01:24.25" resultid="1715" heatid="1941" lane="5" entrytime="00:01:23.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="341" swimtime="00:02:54.36" resultid="1716" heatid="1905" lane="2" entrytime="00:02:50.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:24.66" />
                    <SPLIT distance="150" swimtime="00:02:14.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="329" swimtime="00:21:54.59" resultid="1717" heatid="1929" lane="2" />
                <RESULT eventid="1270" points="262" swimtime="00:01:25.72" resultid="1718" heatid="1979" lane="6" entrytime="00:01:20.37" entrycourse="SCM" />
                <RESULT eventid="1200" points="365" swimtime="00:05:23.38" resultid="1719" heatid="1955" lane="3" entrytime="00:05:14.63" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Do Prado Martins" birthdate="2008-10-17" gender="F" nation="BRA" license="369419" swrid="5596893" athleteid="1702" externalid="369419">
              <RESULTS>
                <RESULT eventid="1160" points="442" swimtime="00:01:10.93" resultid="1703" heatid="1941" lane="4" entrytime="00:01:11.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="426" swimtime="00:01:06.74" resultid="1704" heatid="1919" lane="5" entrytime="00:01:06.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="465" swimtime="00:02:37.19" resultid="1705" heatid="1906" lane="4" entrytime="00:02:36.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:15.17" />
                    <SPLIT distance="150" swimtime="00:02:00.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="455" swimtime="00:01:21.06" resultid="1706" heatid="1966" lane="3" entrytime="00:01:19.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="432" swimtime="00:05:05.80" resultid="1707" heatid="1956" lane="1" entrytime="00:05:02.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                    <SPLIT distance="100" swimtime="00:01:13.40" />
                    <SPLIT distance="150" swimtime="00:01:52.37" />
                    <SPLIT distance="200" swimtime="00:02:31.64" />
                    <SPLIT distance="250" swimtime="00:03:10.68" />
                    <SPLIT distance="300" swimtime="00:03:49.63" />
                    <SPLIT distance="350" swimtime="00:04:28.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Rinaldini" birthdate="2009-04-09" gender="M" nation="BRA" license="348289" swrid="5596932" athleteid="1649" externalid="348289">
              <RESULTS>
                <RESULT eventid="1168" points="388" swimtime="00:01:05.50" resultid="1650" heatid="1944" lane="6" entrytime="00:01:05.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="411" swimtime="00:02:27.45" resultid="1651" heatid="1911" lane="6" entrytime="00:02:23.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:09.89" />
                    <SPLIT distance="150" swimtime="00:01:54.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="534" swimtime="00:17:23.57" resultid="1652" heatid="1932" lane="3" entrytime="00:17:44.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:17:23.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="378" swimtime="00:00:30.08" resultid="1653" heatid="1971" lane="3" />
                <RESULT eventid="1192" points="505" swimtime="00:04:26.47" resultid="1654" heatid="1952" lane="6" entrytime="00:04:26.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.27" />
                    <SPLIT distance="100" swimtime="00:01:04.49" />
                    <SPLIT distance="150" swimtime="00:01:38.53" />
                    <SPLIT distance="200" swimtime="00:02:12.75" />
                    <SPLIT distance="250" swimtime="00:02:46.52" />
                    <SPLIT distance="300" swimtime="00:03:20.50" />
                    <SPLIT distance="350" swimtime="00:03:54.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Mariotti De Castro" birthdate="2008-06-27" gender="M" nation="BRA" license="329200" swrid="5596912" athleteid="1637" externalid="329200">
              <RESULTS>
                <RESULT eventid="1096" points="481" swimtime="00:00:57.22" resultid="1638" heatid="1923" lane="2" entrytime="00:00:56.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="517" swimtime="00:02:16.54" resultid="1639" heatid="1911" lane="3" entrytime="00:02:12.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                    <SPLIT distance="100" swimtime="00:01:04.48" />
                    <SPLIT distance="150" swimtime="00:01:45.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="332" swimtime="00:01:09.73" resultid="1640" heatid="1983" lane="1" entrytime="00:01:04.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" status="DSQ" swimtime="00:00:29.54" resultid="1641" heatid="1971" lane="4" />
                <RESULT eventid="1192" points="591" swimtime="00:04:12.81" resultid="1642" heatid="1952" lane="3" entrytime="00:04:09.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.50" />
                    <SPLIT distance="100" swimtime="00:01:01.14" />
                    <SPLIT distance="150" swimtime="00:01:33.42" />
                    <SPLIT distance="200" swimtime="00:02:05.89" />
                    <SPLIT distance="250" swimtime="00:02:37.83" />
                    <SPLIT distance="300" swimtime="00:03:10.20" />
                    <SPLIT distance="350" swimtime="00:03:42.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Pedro Signor" birthdate="2005-12-20" gender="M" nation="BRA" license="375814" swrid="5596925" athleteid="1738" externalid="375814">
              <RESULTS>
                <RESULT eventid="1168" points="417" swimtime="00:01:03.95" resultid="1739" heatid="1944" lane="1" entrytime="00:01:04.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="373" swimtime="00:02:32.19" resultid="1740" heatid="1907" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                    <SPLIT distance="100" swimtime="00:01:10.85" />
                    <SPLIT distance="150" swimtime="00:01:58.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="463" swimtime="00:00:28.10" resultid="1741" heatid="1972" lane="4" entrytime="00:00:27.50" entrycourse="SCM" />
                <RESULT eventid="1236" points="360" swimtime="00:01:17.68" resultid="1742" heatid="1969" lane="6" entrytime="00:01:18.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" status="DSQ" swimtime="00:05:02.38" resultid="1743" heatid="1950" lane="5" entrytime="00:05:07.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:12.63" />
                    <SPLIT distance="150" swimtime="00:01:50.34" />
                    <SPLIT distance="200" swimtime="00:02:27.64" />
                    <SPLIT distance="250" swimtime="00:03:05.26" />
                    <SPLIT distance="300" swimtime="00:03:43.32" />
                    <SPLIT distance="350" swimtime="00:04:24.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Pedro Serafini" birthdate="2012-05-15" gender="M" nation="BRA" license="365488" swrid="5596924" athleteid="1798" externalid="365488">
              <RESULTS>
                <RESULT eventid="1151" points="123" swimtime="00:00:44.34" resultid="1799" heatid="1937" lane="4" entrytime="00:00:45.46" entrycourse="SCM" />
                <RESULT eventid="1107" points="168" swimtime="00:02:59.78" resultid="1800" heatid="1925" lane="4" entrytime="00:03:12.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                    <SPLIT distance="100" swimtime="00:01:26.40" />
                    <SPLIT distance="150" swimtime="00:02:24.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="162" swimtime="00:00:36.93" resultid="1801" heatid="1991" lane="1" entrytime="00:00:37.33" entrycourse="SCM" />
                <RESULT eventid="1267" points="138" swimtime="00:01:35.27" resultid="1802" heatid="1976" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Zimmermann" birthdate="2010-01-19" gender="M" nation="BRA" license="357160" swrid="5588977" athleteid="1673" externalid="357160">
              <RESULTS>
                <RESULT eventid="1068" points="444" swimtime="00:02:23.61" resultid="1674" heatid="1911" lane="1" entrytime="00:02:23.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:08.69" />
                    <SPLIT distance="150" swimtime="00:01:50.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="510" swimtime="00:17:39.89" resultid="1675" heatid="1932" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:17:39.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="369" swimtime="00:01:07.37" resultid="1676" heatid="1982" lane="5" entrytime="00:01:08.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="338" swimtime="00:01:19.31" resultid="1677" heatid="1969" lane="1" entrytime="00:01:17.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="494" swimtime="00:04:28.33" resultid="1678" heatid="1951" lane="3" entrytime="00:04:31.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                    <SPLIT distance="100" swimtime="00:01:05.38" />
                    <SPLIT distance="150" swimtime="00:01:39.46" />
                    <SPLIT distance="200" swimtime="00:02:13.73" />
                    <SPLIT distance="250" swimtime="00:02:47.87" />
                    <SPLIT distance="300" swimtime="00:03:22.52" />
                    <SPLIT distance="350" swimtime="00:03:56.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Paiz Ribeiro" birthdate="2006-02-17" gender="M" nation="BRA" license="297583" swrid="5596921" athleteid="1631" externalid="297583">
              <RESULTS>
                <RESULT eventid="1168" points="468" swimtime="00:01:01.50" resultid="1632" heatid="1944" lane="2" entrytime="00:01:00.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="437" swimtime="00:02:24.36" resultid="1633" heatid="1911" lane="4" entrytime="00:02:18.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                    <SPLIT distance="100" swimtime="00:01:08.60" />
                    <SPLIT distance="150" swimtime="00:01:51.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="338" swimtime="00:01:09.37" resultid="1634" heatid="1980" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="388" swimtime="00:01:15.73" resultid="1635" heatid="1969" lane="2" entrytime="00:01:12.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="483" swimtime="00:04:30.38" resultid="1636" heatid="1952" lane="5" entrytime="00:04:25.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                    <SPLIT distance="100" swimtime="00:01:04.93" />
                    <SPLIT distance="150" swimtime="00:01:38.98" />
                    <SPLIT distance="200" swimtime="00:02:13.10" />
                    <SPLIT distance="250" swimtime="00:02:47.46" />
                    <SPLIT distance="300" swimtime="00:03:21.92" />
                    <SPLIT distance="350" swimtime="00:03:56.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Luis Lottermann" birthdate="2014-10-08" gender="M" nation="BRA" license="382237" swrid="5596908" athleteid="1770" externalid="382237">
              <RESULTS>
                <RESULT eventid="1113" points="154" swimtime="00:01:23.55" resultid="1771" heatid="1928" lane="3" entrytime="00:01:20.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="103" swimtime="00:00:53.06" resultid="1772" heatid="1916" lane="4" entrytime="00:00:56.51" entrycourse="SCM" />
                <RESULT eventid="1215" points="99" swimtime="00:00:46.87" resultid="1773" heatid="1959" lane="3" entrytime="00:00:45.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Breno" lastname="Zanella Janke" birthdate="2011-04-26" gender="M" nation="BRA" license="365697" swrid="5588970" athleteid="1708" externalid="365697">
              <RESULTS>
                <RESULT eventid="1068" points="354" swimtime="00:02:34.96" resultid="1709" heatid="1909" lane="3" entrytime="00:02:36.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:12.30" />
                    <SPLIT distance="150" swimtime="00:01:58.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="369" swimtime="00:19:40.58" resultid="1710" heatid="1932" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:19:40.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="235" swimtime="00:01:18.26" resultid="1711" heatid="1981" lane="1" entrytime="00:01:20.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="276" swimtime="00:01:24.81" resultid="1712" heatid="1968" lane="2" entrytime="00:01:25.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="325" swimtime="00:05:08.62" resultid="1713" heatid="1950" lane="2" entrytime="00:05:01.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:14.22" />
                    <SPLIT distance="150" swimtime="00:01:53.96" />
                    <SPLIT distance="200" swimtime="00:02:33.49" />
                    <SPLIT distance="250" swimtime="00:03:12.92" />
                    <SPLIT distance="300" swimtime="00:03:52.20" />
                    <SPLIT distance="350" swimtime="00:04:31.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Colaco Da Conceicao" birthdate="2011-05-25" gender="F" nation="BRA" license="369535" swrid="5588601" athleteid="1720" externalid="369535">
              <RESULTS>
                <RESULT eventid="1060" points="276" swimtime="00:03:06.97" resultid="1721" heatid="1905" lane="1" entrytime="00:03:00.48" entrycourse="SCM" />
                <RESULT eventid="1116" points="337" swimtime="00:21:45.02" resultid="1722" heatid="1930" lane="1" />
                <RESULT eventid="1270" points="245" swimtime="00:01:27.72" resultid="1723" heatid="1977" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1244" points="225" swimtime="00:00:40.06" resultid="1724" heatid="1970" lane="2" entrytime="00:00:42.42" entrycourse="SCM" />
                <RESULT eventid="1200" points="350" swimtime="00:05:28.12" resultid="1725" heatid="1954" lane="5" entrytime="00:05:49.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                    <SPLIT distance="100" swimtime="00:01:16.44" />
                    <SPLIT distance="150" swimtime="00:01:57.44" />
                    <SPLIT distance="200" swimtime="00:02:37.83" />
                    <SPLIT distance="250" swimtime="00:03:20.07" />
                    <SPLIT distance="300" swimtime="00:04:02.42" />
                    <SPLIT distance="350" swimtime="00:04:46.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Bonamigo" birthdate="2013-06-25" gender="M" nation="BRA" license="365484" swrid="5588558" athleteid="1803" externalid="365484">
              <RESULTS>
                <RESULT eventid="1107" points="212" swimtime="00:02:46.47" resultid="1804" heatid="1926" lane="5" entrytime="00:02:51.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                    <SPLIT distance="100" swimtime="00:01:21.30" />
                    <SPLIT distance="150" swimtime="00:02:05.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="202" swimtime="00:01:34.11" resultid="1805" heatid="1913" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="201" swimtime="00:00:34.41" resultid="1806" heatid="1991" lane="2" entrytime="00:00:33.62" entrycourse="SCM" />
                <RESULT eventid="1267" points="192" swimtime="00:01:25.33" resultid="1807" heatid="1976" lane="3" entrytime="00:01:27.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Domingues" birthdate="2013-10-22" gender="M" nation="BRA" license="380661" swrid="5676301" athleteid="1755" externalid="380661">
              <RESULTS>
                <RESULT eventid="1151" points="95" swimtime="00:00:48.41" resultid="1756" heatid="1937" lane="3" entrytime="00:00:44.33" entrycourse="SCM" />
                <RESULT eventid="1107" points="157" swimtime="00:03:03.95" resultid="1757" heatid="1925" lane="5" entrytime="00:03:24.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                    <SPLIT distance="100" swimtime="00:01:28.86" />
                    <SPLIT distance="150" swimtime="00:03:03.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" status="DSQ" swimtime="00:01:51.90" resultid="1758" heatid="1976" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1221" points="57" swimtime="00:02:04.02" resultid="1759" heatid="1961" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Macedo Medeiros" birthdate="2012-05-12" gender="M" nation="BRA" license="392015" swrid="4697574" athleteid="1861" externalid="392015">
              <RESULTS>
                <RESULT eventid="1151" points="76" swimtime="00:00:52.14" resultid="1862" heatid="1937" lane="6" entrytime="00:00:53.38" entrycourse="SCM" />
                <RESULT eventid="1107" points="139" swimtime="00:03:11.42" resultid="1863" heatid="1925" lane="3" entrytime="00:03:11.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                    <SPLIT distance="100" swimtime="00:01:32.06" />
                    <SPLIT distance="150" swimtime="00:02:24.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="123" swimtime="00:01:39.06" resultid="1864" heatid="1975" lane="4" />
                <RESULT eventid="1221" points="82" swimtime="00:01:49.64" resultid="1865" heatid="1962" lane="2" entrytime="00:01:48.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raul" lastname="Bonamigo" birthdate="2010-12-01" gender="M" nation="BRA" license="344397" swrid="5588559" athleteid="1786" externalid="344397">
              <RESULTS>
                <RESULT eventid="1168" points="251" swimtime="00:01:15.67" resultid="1787" heatid="1942" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" status="DSQ" swimtime="00:02:33.41" resultid="1788" heatid="1910" lane="1" entrytime="00:02:34.26" entrycourse="SCM" />
                <RESULT eventid="1278" points="317" swimtime="00:01:10.83" resultid="1789" heatid="1981" lane="4" entrytime="00:01:11.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="245" swimtime="00:01:28.23" resultid="1790" heatid="1968" lane="5" entrytime="00:01:26.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="377" swimtime="00:04:53.77" resultid="1791" heatid="1950" lane="4" entrytime="00:04:57.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:12.37" />
                    <SPLIT distance="150" swimtime="00:01:50.15" />
                    <SPLIT distance="200" swimtime="00:02:27.51" />
                    <SPLIT distance="250" swimtime="00:03:04.95" />
                    <SPLIT distance="300" swimtime="00:03:42.28" />
                    <SPLIT distance="350" swimtime="00:04:18.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Luisa Lottermann" birthdate="2011-08-26" gender="F" nation="BRA" license="382238" swrid="5596909" athleteid="1774" externalid="382238">
              <RESULTS>
                <RESULT eventid="1160" points="154" swimtime="00:01:40.71" resultid="1775" heatid="1940" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="259" swimtime="00:03:10.96" resultid="1776" heatid="1904" lane="2" entrytime="00:03:10.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.49" />
                    <SPLIT distance="100" swimtime="00:01:37.60" />
                    <SPLIT distance="150" swimtime="00:02:27.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="258" swimtime="00:23:46.03" resultid="1777" heatid="1930" lane="5" />
                <RESULT eventid="1228" points="268" swimtime="00:01:36.70" resultid="1778" heatid="1966" lane="1" entrytime="00:01:36.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="280" swimtime="00:05:53.22" resultid="1779" heatid="1953" lane="3" entrytime="00:06:23.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                    <SPLIT distance="100" swimtime="00:01:26.01" />
                    <SPLIT distance="150" swimtime="00:02:11.49" />
                    <SPLIT distance="200" swimtime="00:02:56.80" />
                    <SPLIT distance="250" swimtime="00:03:40.86" />
                    <SPLIT distance="300" swimtime="00:04:25.82" />
                    <SPLIT distance="350" swimtime="00:05:10.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Vitoria Gugel" birthdate="2011-12-08" gender="F" nation="BRA" license="365490" swrid="5588960" athleteid="1866" externalid="365490">
              <RESULTS>
                <RESULT eventid="1160" points="208" swimtime="00:01:31.18" resultid="1867" heatid="1940" lane="3" entrytime="00:01:34.99" entrycourse="SCM" />
                <RESULT eventid="1060" points="304" swimtime="00:03:01.10" resultid="1868" heatid="1905" lane="6" entrytime="00:03:00.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.22" />
                    <SPLIT distance="100" swimtime="00:01:26.98" />
                    <SPLIT distance="150" swimtime="00:02:20.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="248" swimtime="00:01:27.25" resultid="1869" heatid="1978" lane="1" entrytime="00:01:23.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="262" swimtime="00:01:37.41" resultid="1870" heatid="1966" lane="5" entrytime="00:01:36.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="317" swimtime="00:05:38.99" resultid="1871" heatid="1954" lane="2" entrytime="00:05:45.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                    <SPLIT distance="100" swimtime="00:01:19.44" />
                    <SPLIT distance="150" swimtime="00:02:02.43" />
                    <SPLIT distance="200" swimtime="00:02:45.41" />
                    <SPLIT distance="250" swimtime="00:03:29.43" />
                    <SPLIT distance="300" swimtime="00:04:12.94" />
                    <SPLIT distance="350" swimtime="00:04:56.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabelle" lastname="Cordeiro Silva" birthdate="2015-06-14" gender="F" nation="BRA" license="390839" swrid="5596878" athleteid="1819" externalid="390839">
              <RESULTS>
                <RESULT eventid="1154" status="WDR" swimtime="00:00:00.00" resultid="1820" heatid="1938" lane="3" entrytime="00:00:51.43" entrycourse="SCM" />
                <RESULT eventid="1082" status="WDR" swimtime="00:00:00.00" resultid="1821" heatid="1915" lane="5" entrytime="00:00:59.78" entrycourse="SCM" />
                <RESULT eventid="1290" status="WDR" swimtime="00:00:00.00" resultid="1822" heatid="1987" lane="6" entrytime="00:00:45.93" entrycourse="SCM" />
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="1823" heatid="1958" lane="4" entrytime="00:00:54.05" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Tolentino Smarczewski" birthdate="2008-09-01" gender="M" nation="BRA" license="378818" swrid="5596941" athleteid="1744" externalid="378818">
              <RESULTS>
                <RESULT eventid="1168" points="251" swimtime="00:01:15.72" resultid="1745" heatid="1943" lane="2" entrytime="00:01:15.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="434" swimtime="00:00:59.21" resultid="1746" heatid="1922" lane="4" entrytime="00:01:00.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="360" swimtime="00:02:34.08" resultid="1747" heatid="1910" lane="6" entrytime="00:02:35.43" entrycourse="SCM" />
                <RESULT eventid="1236" points="305" swimtime="00:01:22.10" resultid="1748" heatid="1968" lane="4" entrytime="00:01:23.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="429" swimtime="00:04:41.33" resultid="1749" heatid="1951" lane="2" entrytime="00:04:32.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                    <SPLIT distance="100" swimtime="00:01:08.28" />
                    <SPLIT distance="150" swimtime="00:01:44.23" />
                    <SPLIT distance="200" swimtime="00:02:21.22" />
                    <SPLIT distance="250" swimtime="00:02:56.19" />
                    <SPLIT distance="300" swimtime="00:03:30.95" />
                    <SPLIT distance="350" swimtime="00:04:06.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Balduíno" birthdate="2009-06-24" gender="M" nation="BRA" license="370764" swrid="5596870" athleteid="1732" externalid="370764">
              <RESULTS>
                <RESULT eventid="1168" points="405" swimtime="00:01:04.57" resultid="1733" heatid="1943" lane="3" entrytime="00:01:05.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="417" swimtime="00:02:26.70" resultid="1734" heatid="1910" lane="2" entrytime="00:02:27.33" entrycourse="SCM" />
                <RESULT eventid="1278" points="322" swimtime="00:01:10.46" resultid="1735" heatid="1982" lane="6" entrytime="00:01:09.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="311" swimtime="00:01:21.51" resultid="1736" heatid="1968" lane="3" entrytime="00:01:20.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="429" swimtime="00:04:41.33" resultid="1737" heatid="1951" lane="1" entrytime="00:04:43.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                    <SPLIT distance="100" swimtime="00:01:08.02" />
                    <SPLIT distance="150" swimtime="00:01:43.96" />
                    <SPLIT distance="200" swimtime="00:02:20.09" />
                    <SPLIT distance="250" swimtime="00:02:55.92" />
                    <SPLIT distance="300" swimtime="00:03:31.30" />
                    <SPLIT distance="350" swimtime="00:04:06.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose" lastname="Eliziario Filho" birthdate="2014-03-27" gender="M" nation="BRA" license="406696" athleteid="1882" externalid="406696">
              <RESULTS>
                <RESULT eventid="1157" points="59" swimtime="00:00:56.64" resultid="1883" heatid="1939" lane="4" />
                <RESULT eventid="1113" points="105" swimtime="00:01:35.02" resultid="1884" heatid="1928" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1293" points="109" swimtime="00:00:42.17" resultid="1885" heatid="1988" lane="1" />
                <RESULT eventid="1215" points="87" swimtime="00:00:48.90" resultid="1886" heatid="1959" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Bezerra Sedlacek" birthdate="2014-02-26" gender="M" nation="BRA" license="380663" swrid="4300166" athleteid="1760" externalid="380663">
              <RESULTS>
                <RESULT eventid="1113" points="95" swimtime="00:01:37.94" resultid="1761" heatid="1928" lane="2" entrytime="00:01:43.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="106" swimtime="00:00:52.58" resultid="1762" heatid="1916" lane="3" entrytime="00:00:53.70" entrycourse="SCM" />
                <RESULT eventid="1293" points="97" swimtime="00:00:43.79" resultid="1763" heatid="1988" lane="4" entrytime="00:00:42.09" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia" lastname="Oliveira Faria" birthdate="2013-10-04" gender="F" nation="BRA" license="406697" athleteid="1887" externalid="406697">
              <RESULTS>
                <RESULT eventid="1148" points="76" swimtime="00:00:59.39" resultid="1888" heatid="1935" lane="5" />
                <RESULT eventid="1104" points="86" swimtime="00:04:09.43" resultid="1889" heatid="1924" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.43" />
                    <SPLIT distance="100" swimtime="00:01:57.72" />
                    <SPLIT distance="150" swimtime="00:03:03.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="103" swimtime="00:00:48.76" resultid="1890" heatid="1989" lane="6" />
                <RESULT eventid="1264" points="77" swimtime="00:02:12.47" resultid="1891" heatid="1973" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Cordeiro Silva" birthdate="2011-09-04" gender="M" nation="BRA" license="380664" swrid="5596877" athleteid="1764" externalid="380664">
              <RESULTS>
                <RESULT eventid="1168" status="WDR" swimtime="00:00:00.00" resultid="1765" heatid="1942" lane="1" />
                <RESULT eventid="1096" status="WDR" swimtime="00:00:00.00" resultid="1766" heatid="1921" lane="5" entrytime="00:01:15.66" entrycourse="SCM" />
                <RESULT eventid="1068" status="WDR" swimtime="00:00:00.00" resultid="1767" heatid="1908" lane="4" entrytime="00:02:57.90" entrycourse="SCM" />
                <RESULT eventid="1236" status="WDR" swimtime="00:00:00.00" resultid="1768" heatid="1967" lane="2" entrytime="00:01:31.02" entrycourse="SCM" />
                <RESULT eventid="1192" status="WDR" swimtime="00:00:00.00" resultid="1769" heatid="1949" lane="5" entrytime="00:05:40.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Vargas Moreira" birthdate="2014-03-09" gender="F" nation="BRA" license="392014" swrid="4904290" athleteid="1856" externalid="392014">
              <RESULTS>
                <RESULT eventid="1110" points="177" swimtime="00:01:29.46" resultid="1857" heatid="1927" lane="4" entrytime="00:01:32.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1082" points="123" swimtime="00:00:57.04" resultid="1858" heatid="1915" lane="2" entrytime="00:00:57.02" entrycourse="SCM" />
                <RESULT eventid="1290" points="180" swimtime="00:00:40.59" resultid="1859" heatid="1987" lane="4" entrytime="00:00:41.07" entrycourse="SCM" />
                <RESULT eventid="1212" points="98" swimtime="00:00:52.72" resultid="1860" heatid="1958" lane="1" entrytime="00:01:00.81" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Dillenburg Benetti" birthdate="2011-03-10" gender="M" nation="BRA" license="368119" swrid="5588656" athleteid="1691" externalid="368119">
              <RESULTS>
                <RESULT eventid="1068" points="330" swimtime="00:02:38.54" resultid="1692" heatid="1909" lane="4" entrytime="00:02:43.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:01:15.44" />
                    <SPLIT distance="150" swimtime="00:02:01.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="348" swimtime="00:20:03.02" resultid="1693" heatid="1932" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:20:03.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="284" swimtime="00:01:13.52" resultid="1694" heatid="1981" lane="2" entrytime="00:01:14.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" status="DSQ" swimtime="00:01:26.16" resultid="1695" heatid="1968" lane="1" entrytime="00:01:28.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="319" swimtime="00:05:10.37" resultid="1696" heatid="1950" lane="1" entrytime="00:05:16.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:14.15" />
                    <SPLIT distance="150" swimtime="00:01:54.19" />
                    <SPLIT distance="200" swimtime="00:02:33.85" />
                    <SPLIT distance="250" swimtime="00:03:13.24" />
                    <SPLIT distance="300" swimtime="00:03:52.72" />
                    <SPLIT distance="350" swimtime="00:04:31.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Assakura" birthdate="2010-06-29" gender="F" nation="BRA" license="376473" swrid="5596868" athleteid="1780" externalid="376473">
              <RESULTS>
                <RESULT eventid="1088" points="379" swimtime="00:01:09.39" resultid="1781" heatid="1918" lane="2" entrytime="00:01:10.30" entrycourse="SCM" />
                <RESULT eventid="1060" points="388" swimtime="00:02:46.96" resultid="1782" heatid="1905" lane="4" entrytime="00:02:50.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                    <SPLIT distance="100" swimtime="00:01:21.97" />
                    <SPLIT distance="150" swimtime="00:02:08.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="314" swimtime="00:01:20.72" resultid="1783" heatid="1978" lane="5" entrytime="00:01:21.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="374" swimtime="00:01:26.54" resultid="1784" heatid="1966" lane="4" entrytime="00:01:24.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="405" swimtime="00:05:12.46" resultid="1785" heatid="1954" lane="6" entrytime="00:06:02.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                    <SPLIT distance="100" swimtime="00:01:14.27" />
                    <SPLIT distance="150" swimtime="00:01:53.94" />
                    <SPLIT distance="200" swimtime="00:02:33.60" />
                    <SPLIT distance="250" swimtime="00:03:14.62" />
                    <SPLIT distance="300" swimtime="00:03:54.97" />
                    <SPLIT distance="350" swimtime="00:04:36.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Borille Busetti" birthdate="2010-02-17" gender="F" nation="BRA" license="392830" swrid="5622263" athleteid="1872" externalid="392830">
              <RESULTS>
                <RESULT eventid="1088" points="332" swimtime="00:01:12.52" resultid="1873" heatid="1918" lane="5" entrytime="00:01:12.65" entrycourse="SCM" />
                <RESULT eventid="1060" points="201" swimtime="00:03:27.89" resultid="1874" heatid="1904" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.33" />
                    <SPLIT distance="100" swimtime="00:01:36.44" />
                    <SPLIT distance="150" swimtime="00:03:21.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="245" swimtime="00:01:27.64" resultid="1875" heatid="1977" lane="3" entrytime="00:01:31.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="177" swimtime="00:01:50.92" resultid="1876" heatid="1965" lane="4" entrytime="00:01:51.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="262" swimtime="00:06:01.43" resultid="1877" heatid="1954" lane="1" entrytime="00:05:57.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:01:20.02" />
                    <SPLIT distance="150" swimtime="00:02:05.53" />
                    <SPLIT distance="200" swimtime="00:02:52.15" />
                    <SPLIT distance="250" swimtime="00:03:39.61" />
                    <SPLIT distance="300" swimtime="00:04:28.54" />
                    <SPLIT distance="350" swimtime="00:05:16.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emanuel" lastname="Ranieri" birthdate="2011-01-24" gender="M" nation="BRA" license="390838" swrid="5596930" athleteid="1813" externalid="390838">
              <RESULTS>
                <RESULT eventid="1068" points="295" swimtime="00:02:44.62" resultid="1814" heatid="1909" lane="2" entrytime="00:02:44.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                    <SPLIT distance="100" swimtime="00:01:19.53" />
                    <SPLIT distance="150" swimtime="00:02:07.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="282" swimtime="00:21:29.93" resultid="1815" heatid="1931" lane="5" />
                <RESULT eventid="1278" points="201" swimtime="00:01:22.37" resultid="1816" heatid="1981" lane="6" entrytime="00:01:21.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="226" swimtime="00:01:30.63" resultid="1817" heatid="1967" lane="3" entrytime="00:01:29.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="293" swimtime="00:05:19.46" resultid="1818" heatid="1949" lane="4" entrytime="00:05:22.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:01:16.53" />
                    <SPLIT distance="150" swimtime="00:01:57.75" />
                    <SPLIT distance="200" swimtime="00:02:39.61" />
                    <SPLIT distance="250" swimtime="00:03:21.69" />
                    <SPLIT distance="300" swimtime="00:04:03.13" />
                    <SPLIT distance="350" swimtime="00:04:42.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Danilo" lastname="Rodrigues" birthdate="2011-05-23" gender="M" nation="BRA" license="370763" swrid="5596934" athleteid="1726" externalid="370763">
              <RESULTS>
                <RESULT eventid="1168" points="217" swimtime="00:01:19.45" resultid="1727" heatid="1943" lane="1" entrytime="00:01:19.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="281" swimtime="00:02:47.24" resultid="1728" heatid="1909" lane="1" entrytime="00:02:47.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:20.76" />
                    <SPLIT distance="150" swimtime="00:02:09.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="310" swimtime="00:20:51.17" resultid="1729" heatid="1932" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:20:51.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="240" swimtime="00:01:28.93" resultid="1730" heatid="1967" lane="4" entrytime="00:01:30.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="297" swimtime="00:05:17.94" resultid="1731" heatid="1950" lane="6" entrytime="00:05:19.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Gaio" birthdate="2012-11-13" gender="F" nation="BRA" license="390842" swrid="5596901" athleteid="1829" externalid="390842">
              <RESULTS>
                <RESULT eventid="1148" points="60" swimtime="00:01:04.18" resultid="1830" heatid="1935" lane="2" entrytime="00:01:04.13" entrycourse="SCM" />
                <RESULT eventid="1104" points="72" swimtime="00:04:24.23" resultid="1831" heatid="1924" lane="4" entrytime="00:04:26.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.91" />
                    <SPLIT distance="100" swimtime="00:02:05.37" />
                    <SPLIT distance="150" swimtime="00:03:16.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="66" swimtime="00:02:19.35" resultid="1832" heatid="1973" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1218" points="43" swimtime="00:02:34.17" resultid="1833" heatid="1960" lane="4" entrytime="00:02:37.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Stein Duarte" birthdate="2010-10-03" gender="F" nation="BRA" license="351635" swrid="5588923" athleteid="1661" externalid="351635">
              <RESULTS>
                <RESULT eventid="1088" points="360" swimtime="00:01:10.63" resultid="1662" heatid="1917" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="384" swimtime="00:02:47.64" resultid="1663" heatid="1906" lane="1" entrytime="00:02:42.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:01:18.89" />
                    <SPLIT distance="150" swimtime="00:02:07.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="369" swimtime="00:01:16.50" resultid="1664" heatid="1979" lane="4" entrytime="00:01:14.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="313" swimtime="00:01:31.80" resultid="1665" heatid="1966" lane="2" entrytime="00:01:32.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="416" swimtime="00:05:09.84" resultid="1666" heatid="1956" lane="6" entrytime="00:05:09.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:12.86" />
                    <SPLIT distance="150" swimtime="00:01:51.70" />
                    <SPLIT distance="200" swimtime="00:02:31.16" />
                    <SPLIT distance="250" swimtime="00:03:10.51" />
                    <SPLIT distance="300" swimtime="00:03:50.81" />
                    <SPLIT distance="350" swimtime="00:04:30.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gael" lastname="Vicenzo Pereira" birthdate="2012-09-18" gender="M" nation="BRA" license="390847" swrid="5596943" athleteid="1845" externalid="390847">
              <RESULTS>
                <RESULT eventid="1151" points="50" swimtime="00:00:59.67" resultid="1846" heatid="1936" lane="2" />
                <RESULT eventid="1107" points="68" swimtime="00:04:02.77" resultid="1847" heatid="1925" lane="1" entrytime="00:03:57.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.16" />
                    <SPLIT distance="100" swimtime="00:01:50.68" />
                    <SPLIT distance="150" swimtime="00:02:57.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="65" swimtime="00:00:49.97" resultid="1848" heatid="1990" lane="5" entrytime="00:00:48.04" entrycourse="SCM" />
                <RESULT eventid="1221" status="DSQ" swimtime="00:02:40.20" resultid="1849" heatid="1962" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laisa" lastname="Bernardini" birthdate="2012-06-25" gender="F" nation="BRA" license="390843" swrid="5596872" athleteid="1834" externalid="390843">
              <RESULTS>
                <RESULT eventid="1104" points="177" swimtime="00:03:16.10" resultid="1835" heatid="1924" lane="3" entrytime="00:03:06.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.29" />
                    <SPLIT distance="100" swimtime="00:01:34.23" />
                    <SPLIT distance="150" swimtime="00:02:26.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1076" points="194" swimtime="00:01:47.59" resultid="1836" heatid="1912" lane="4" entrytime="00:02:01.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="182" swimtime="00:01:39.56" resultid="1837" heatid="1973" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1218" points="122" swimtime="00:01:48.90" resultid="1838" heatid="1960" lane="3" entrytime="00:01:45.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
