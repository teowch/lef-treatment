<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.79125">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Toledo" name="Torneio Regional da 3ª Região (Pré-Mirim/Sênior)" course="SCM" deadline="2024-03-11" entrystartdate="2024-03-04" entrytype="INVITATION" hostclub="Prefeitura Municipal de Toledo" hostclub.url="https://www.toledo.pr.gov.br/" number="38300" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/evento/natacao/38300" startmethod="1" timing="AUTOMATIC" masters="F" withdrawuntil="2024-03-13" state="PR" nation="BRA">
      <AGEDATE value="2024-03-16" type="YEAR" />
      <POOL name="Piscina Municipal Claus Fuchs" lanemin="1" lanemax="6" />
      <FACILITY city="Toledo" name="Piscina Municipal Claus Fuchs" nation="BRA" state="PR" street="Rua Guanabara, 1040" street2="Jardim Santa Maria" zip="85903-040" />
      <POINTTABLE pointtableid="3016" name="FINA Point Scoring" version="2023" />
      <QUALIFY from="2023-03-16" until="2024-03-15" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99206-4448" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99206-4448" street="Avenida do Batel, 1230" street2="Batel" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-03-16" daytime="09:10" endtime="13:18" number="1" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1060" daytime="09:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1950" />
                    <RANKING order="2" place="2" resultid="1844" />
                    <RANKING order="3" place="3" resultid="1716" />
                    <RANKING order="4" place="4" resultid="1866" />
                    <RANKING order="5" place="5" resultid="1344" />
                    <RANKING order="6" place="6" resultid="1567" />
                    <RANKING order="7" place="7" resultid="1325" />
                    <RANKING order="8" place="8" resultid="1585" />
                    <RANKING order="9" place="-1" resultid="1944" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1932" />
                    <RANKING order="2" place="2" resultid="1312" />
                    <RANKING order="3" place="3" resultid="1506" />
                    <RANKING order="4" place="4" resultid="1361" />
                    <RANKING order="5" place="5" resultid="1937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1352" />
                    <RANKING order="2" place="2" resultid="1476" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1065" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1630" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1436" />
                    <RANKING order="2" place="2" resultid="1920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1625" />
                    <RANKING order="2" place="2" resultid="1914" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1959" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1960" daytime="09:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1961" daytime="09:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="1962" daytime="09:18" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1068" daytime="09:20" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1069" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1688" />
                    <RANKING order="2" place="2" resultid="1576" />
                    <RANKING order="3" place="3" resultid="1850" />
                    <RANKING order="4" place="4" resultid="1367" />
                    <RANKING order="5" place="5" resultid="1771" />
                    <RANKING order="6" place="6" resultid="1393" />
                    <RANKING order="7" place="7" resultid="1378" />
                    <RANKING order="8" place="8" resultid="1571" />
                    <RANKING order="9" place="-1" resultid="1955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1670" />
                    <RANKING order="2" place="2" resultid="1552" />
                    <RANKING order="3" place="3" resultid="1676" />
                    <RANKING order="4" place="-1" resultid="1517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1646" />
                    <RANKING order="2" place="2" resultid="1481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1331" />
                    <RANKING order="2" place="2" resultid="1908" />
                    <RANKING order="3" place="3" resultid="1799" />
                    <RANKING order="4" place="4" resultid="1430" />
                    <RANKING order="5" place="5" resultid="1500" />
                    <RANKING order="6" place="6" resultid="1488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1471" />
                    <RANKING order="2" place="2" resultid="1494" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1449" />
                    <RANKING order="2" place="2" resultid="1459" />
                    <RANKING order="3" place="3" resultid="1926" />
                    <RANKING order="4" place="4" resultid="1741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1321" />
                    <RANKING order="2" place="2" resultid="1443" />
                    <RANKING order="3" place="3" resultid="1316" />
                    <RANKING order="4" place="-1" resultid="1616" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1963" daytime="09:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1964" daytime="09:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1965" daytime="09:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="1966" daytime="09:28" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="1967" daytime="09:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="1968" daytime="09:32" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1076" daytime="09:34" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1077" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1078" daytime="09:34" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1079" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1080" daytime="09:34" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1081" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1855" />
                    <RANKING order="2" place="2" resultid="1522" />
                    <RANKING order="3" place="3" resultid="1752" />
                    <RANKING order="4" place="4" resultid="1558" />
                    <RANKING order="5" place="5" resultid="1815" />
                    <RANKING order="6" place="6" resultid="1542" />
                    <RANKING order="7" place="7" resultid="1897" />
                    <RANKING order="8" place="8" resultid="1829" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1969" daytime="09:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1970" daytime="09:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1083" daytime="09:44" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1084" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="1085" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1776" />
                    <RANKING order="2" place="2" resultid="1547" />
                    <RANKING order="3" place="3" resultid="1765" />
                    <RANKING order="4" place="4" resultid="1887" />
                    <RANKING order="5" place="5" resultid="1877" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1971" daytime="09:44" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1086" daytime="09:50" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1087" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1892" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1511" />
                    <RANKING order="2" place="2" resultid="1838" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1972" daytime="09:50" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1089" daytime="09:54" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1090" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1755" />
                    <RANKING order="2" place="2" resultid="1537" />
                    <RANKING order="3" place="-1" resultid="1760" />
                    <RANKING order="4" place="-1" resultid="1810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1532" />
                    <RANKING order="2" place="2" resultid="1699" />
                    <RANKING order="3" place="3" resultid="1805" />
                    <RANKING order="4" place="-1" resultid="1860" />
                    <RANKING order="5" place="-1" resultid="1563" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1973" daytime="09:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1974" daytime="10:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1092" daytime="10:04" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1093" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1781" />
                    <RANKING order="2" place="2" resultid="1865" />
                    <RANKING order="3" place="3" resultid="1324" />
                    <RANKING order="4" place="-1" resultid="1949" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1788" />
                    <RANKING order="2" place="2" resultid="1658" />
                    <RANKING order="3" place="3" resultid="1936" />
                    <RANKING order="4" place="-1" resultid="1872" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1096" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1652" />
                    <RANKING order="2" place="2" resultid="1704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1427" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1099" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1640" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1975" daytime="10:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1976" daytime="10:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1100" daytime="10:16" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1101" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1711" />
                    <RANKING order="2" place="2" resultid="1693" />
                    <RANKING order="3" place="3" resultid="1728" />
                    <RANKING order="4" place="4" resultid="1819" />
                    <RANKING order="5" place="5" resultid="1770" />
                    <RANKING order="6" place="6" resultid="1849" />
                    <RANKING order="7" place="7" resultid="1575" />
                    <RANKING order="8" place="8" resultid="1337" />
                    <RANKING order="9" place="9" resultid="1381" />
                    <RANKING order="10" place="-1" resultid="1954" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1669" />
                    <RANKING order="2" place="2" resultid="1793" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1104" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1635" />
                    <RANKING order="2" place="2" resultid="1465" />
                    <RANKING order="3" place="3" resultid="1746" />
                    <RANKING order="4" place="4" resultid="1499" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1681" />
                    <RANKING order="2" place="2" resultid="1493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1925" />
                    <RANKING order="2" place="2" resultid="1341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1107" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1977" daytime="10:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1978" daytime="10:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1979" daytime="10:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="1980" daytime="10:28" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1108" daytime="10:32" gender="F" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1109" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1405" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1981" daytime="10:32" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1110" daytime="10:36" gender="M" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1111" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1593" />
                    <RANKING order="2" place="2" resultid="1402" />
                    <RANKING order="3" place="3" resultid="1411" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1982" daytime="10:36" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1112" daytime="10:52" gender="F" number="13" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1113" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1114" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1814" />
                    <RANKING order="2" place="2" resultid="1541" />
                    <RANKING order="3" place="3" resultid="1751" />
                    <RANKING order="4" place="4" resultid="1557" />
                    <RANKING order="5" place="5" resultid="1828" />
                    <RANKING order="6" place="6" resultid="1408" />
                    <RANKING order="7" place="7" resultid="1397" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1983" daytime="10:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1984" daytime="10:54" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1115" daytime="10:58" gender="M" number="14" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1116" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1389" />
                    <RANKING order="2" place="2" resultid="1882" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1117" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1546" />
                    <RANKING order="2" place="2" resultid="1600" />
                    <RANKING order="3" place="3" resultid="1764" />
                    <RANKING order="4" place="4" resultid="1348" />
                    <RANKING order="5" place="5" resultid="1876" />
                    <RANKING order="6" place="6" resultid="1607" />
                    <RANKING order="7" place="7" resultid="1581" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1985" daytime="10:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1986" daytime="11:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1118" daytime="11:02" gender="F" number="15" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1119" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1374" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1510" />
                    <RANKING order="2" place="2" resultid="1834" />
                    <RANKING order="3" place="3" resultid="1597" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1987" daytime="11:02" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1121" daytime="11:06" gender="M" number="16" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1122" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1527" />
                    <RANKING order="2" place="2" resultid="1536" />
                    <RANKING order="3" place="3" resultid="1400" />
                    <RANKING order="4" place="-1" resultid="1809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1531" />
                    <RANKING order="2" place="2" resultid="1804" />
                    <RANKING order="3" place="3" resultid="1562" />
                    <RANKING order="4" place="-1" resultid="1417" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1988" daytime="11:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1989" daytime="11:08" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1124" daytime="11:12" gender="F" number="17" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1125" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1723" />
                    <RANKING order="2" place="2" resultid="1715" />
                    <RANKING order="3" place="3" resultid="1843" />
                    <RANKING order="4" place="4" resultid="1943" />
                    <RANKING order="5" place="5" resultid="1864" />
                    <RANKING order="6" place="6" resultid="1780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1657" />
                    <RANKING order="2" place="2" resultid="1505" />
                    <RANKING order="3" place="3" resultid="1787" />
                    <RANKING order="4" place="4" resultid="1871" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1475" />
                    <RANKING order="2" place="2" resultid="1663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1651" />
                    <RANKING order="2" place="2" resultid="1703" />
                    <RANKING order="3" place="3" resultid="1328" />
                    <RANKING order="4" place="-1" resultid="1422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1131" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1990" daytime="11:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1991" daytime="11:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1992" daytime="11:36" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1132" daytime="11:50" gender="M" number="18" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1133" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1710" />
                    <RANKING order="2" place="2" resultid="1692" />
                    <RANKING order="3" place="3" resultid="1687" />
                    <RANKING order="4" place="4" resultid="1818" />
                    <RANKING order="5" place="5" resultid="1727" />
                    <RANKING order="6" place="6" resultid="1848" />
                    <RANKING order="7" place="7" resultid="1769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1134" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1668" />
                    <RANKING order="2" place="2" resultid="1792" />
                    <RANKING order="3" place="3" resultid="1675" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1645" />
                    <RANKING order="2" place="2" resultid="1734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1634" />
                    <RANKING order="2" place="2" resultid="1464" />
                    <RANKING order="3" place="3" resultid="1798" />
                    <RANKING order="4" place="4" resultid="1745" />
                    <RANKING order="5" place="5" resultid="1487" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1137" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1680" />
                    <RANKING order="2" place="2" resultid="1470" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1621" />
                    <RANKING order="2" place="2" resultid="1740" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1139" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1615" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1993" daytime="11:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1994" daytime="12:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1995" daytime="12:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="1996" daytime="12:26" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1140" daytime="12:38" gender="F" number="19" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1141" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1842" />
                    <RANKING order="2" place="2" resultid="1722" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1656" />
                    <RANKING order="2" place="2" resultid="1931" />
                    <RANKING order="3" place="3" resultid="1786" />
                    <RANKING order="4" place="4" resultid="1360" />
                    <RANKING order="5" place="5" resultid="1870" />
                    <RANKING order="6" place="6" resultid="1355" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1143" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1144" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1145" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1146" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1435" />
                    <RANKING order="2" place="2" resultid="1919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1639" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1997" daytime="12:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1998" daytime="12:44" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1148" daytime="12:48" gender="M" number="20" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1149" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1817" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1516" />
                    <RANKING order="2" place="2" resultid="1551" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1151" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1152" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1907" />
                    <RANKING order="2" place="2" resultid="1429" />
                    <RANKING order="3" place="3" resultid="1498" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1154" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1448" />
                    <RANKING order="2" place="2" resultid="1458" />
                    <RANKING order="3" place="3" resultid="1620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1442" />
                    <RANKING order="2" place="2" resultid="1454" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1999" daytime="12:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2000" daytime="12:52" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1156" daytime="12:58" gender="F" number="21" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1157" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1823" />
                    <RANKING order="2" place="2" resultid="1385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1370" />
                    <RANKING order="2" place="2" resultid="1521" />
                    <RANKING order="3" place="3" resultid="1854" />
                    <RANKING order="4" place="4" resultid="1896" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2001" daytime="12:58" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1159" daytime="13:00" gender="M" number="22" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1160" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1161" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1775" />
                    <RANKING order="2" place="2" resultid="1886" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2002" daytime="13:00" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1162" daytime="13:02" gender="F" number="23" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1163" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1363" />
                    <RANKING order="2" place="2" resultid="1891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1164" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1837" />
                    <RANKING order="2" place="2" resultid="1833" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2003" daytime="13:02" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1165" daytime="13:04" gender="M" number="24" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1166" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1526" />
                    <RANKING order="2" place="2" resultid="1754" />
                    <RANKING order="3" place="3" resultid="1759" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1698" />
                    <RANKING order="2" place="2" resultid="1859" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2004" daytime="13:04" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1168" daytime="13:08" gender="F" number="25" order="26" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1169" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1942" />
                    <RANKING order="2" place="2" resultid="1721" />
                    <RANKING order="3" place="3" resultid="1948" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1930" />
                    <RANKING order="2" place="2" resultid="1504" />
                    <RANKING order="3" place="3" resultid="1311" />
                    <RANKING order="4" place="4" resultid="1359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1662" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1650" />
                    <RANKING order="2" place="-1" resultid="1421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1174" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1175" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1913" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2005" daytime="13:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2006" daytime="13:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1176" daytime="13:14" gender="M" number="26" order="27" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1177" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1686" />
                    <RANKING order="2" place="2" resultid="1709" />
                    <RANKING order="3" place="3" resultid="1366" />
                    <RANKING order="4" place="4" resultid="1377" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1515" />
                    <RANKING order="2" place="2" resultid="1674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1644" />
                    <RANKING order="2" place="2" resultid="1733" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1180" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1463" />
                    <RANKING order="2" place="2" resultid="1906" />
                    <RANKING order="3" place="3" resultid="1486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1181" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1334" />
                    <RANKING order="2" place="2" resultid="1469" />
                    <RANKING order="3" place="3" resultid="1492" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1447" />
                    <RANKING order="2" place="2" resultid="1739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1183" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1318" />
                    <RANKING order="2" place="2" resultid="1315" />
                    <RANKING order="3" place="3" resultid="1441" />
                    <RANKING order="4" place="4" resultid="1453" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2007" daytime="13:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2008" daytime="13:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2009" daytime="13:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2010" daytime="13:20" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-03-16" daytime="15:40" endtime="19:40" number="2" officialmeeting="15:00" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1184" daytime="15:40" gender="F" number="27" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1185" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1719" />
                    <RANKING order="2" place="2" resultid="1868" />
                    <RANKING order="3" place="3" resultid="1725" />
                    <RANKING order="4" place="4" resultid="1846" />
                    <RANKING order="5" place="5" resultid="1784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1660" />
                    <RANKING order="2" place="2" resultid="1790" />
                    <RANKING order="3" place="3" resultid="1874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1666" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1188" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1654" />
                    <RANKING order="2" place="2" resultid="1707" />
                    <RANKING order="3" place="-1" resultid="1425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1189" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1632" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1191" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2011" daytime="15:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2012" daytime="15:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2013" daytime="15:54" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1192" daytime="16:02" gender="M" number="28" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1193" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1713" />
                    <RANKING order="2" place="2" resultid="1696" />
                    <RANKING order="3" place="3" resultid="1731" />
                    <RANKING order="4" place="4" resultid="1821" />
                    <RANKING order="5" place="5" resultid="1852" />
                    <RANKING order="6" place="6" resultid="1773" />
                    <RANKING order="7" place="-1" resultid="1690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1672" />
                    <RANKING order="2" place="2" resultid="1796" />
                    <RANKING order="3" place="3" resultid="1678" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1648" />
                    <RANKING order="2" place="2" resultid="1737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1196" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1637" />
                    <RANKING order="2" place="2" resultid="1467" />
                    <RANKING order="3" place="3" resultid="1802" />
                    <RANKING order="4" place="4" resultid="1749" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1197" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1623" />
                    <RANKING order="2" place="2" resultid="1743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1199" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2014" daytime="16:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2015" daytime="16:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2016" daytime="16:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2017" daytime="16:22" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1200" daytime="16:28" gender="F" number="29" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1201" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1202" daytime="16:28" gender="M" number="30" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1203" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1595" />
                    <RANKING order="2" place="2" resultid="1415" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2018" daytime="16:28" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1204" daytime="16:30" gender="F" number="31" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1205" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1387" />
                    <RANKING order="2" place="2" resultid="1903" />
                    <RANKING order="3" place="3" resultid="1826" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1206" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1524" />
                    <RANKING order="2" place="2" resultid="1857" />
                    <RANKING order="3" place="3" resultid="1544" />
                    <RANKING order="4" place="4" resultid="1560" />
                    <RANKING order="5" place="5" resultid="1372" />
                    <RANKING order="6" place="6" resultid="1831" />
                    <RANKING order="7" place="7" resultid="1899" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2019" daytime="16:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2020" daytime="16:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1207" daytime="16:38" gender="M" number="32" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1208" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1391" />
                    <RANKING order="2" place="2" resultid="1884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1778" />
                    <RANKING order="2" place="2" resultid="1549" />
                    <RANKING order="3" place="3" resultid="1767" />
                    <RANKING order="4" place="4" resultid="1889" />
                    <RANKING order="5" place="5" resultid="1879" />
                    <RANKING order="6" place="6" resultid="1350" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2021" daytime="16:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2022" daytime="16:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1210" daytime="16:44" gender="F" number="33" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1211" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1894" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1212" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1513" />
                    <RANKING order="2" place="2" resultid="1840" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2023" daytime="16:44" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1213" daytime="16:50" gender="M" number="34" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1214" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1539" />
                    <RANKING order="2" place="2" resultid="1757" />
                    <RANKING order="3" place="3" resultid="1529" />
                    <RANKING order="4" place="-1" resultid="1762" />
                    <RANKING order="5" place="-1" resultid="1812" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1534" />
                    <RANKING order="2" place="2" resultid="1701" />
                    <RANKING order="3" place="3" resultid="1807" />
                    <RANKING order="4" place="4" resultid="1862" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2024" daytime="16:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2025" daytime="16:58" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1216" daytime="17:06" gender="F" number="35" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1217" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1952" />
                    <RANKING order="2" place="2" resultid="1845" />
                    <RANKING order="3" place="3" resultid="1946" />
                    <RANKING order="4" place="4" resultid="1724" />
                    <RANKING order="5" place="5" resultid="1783" />
                    <RANKING order="6" place="6" resultid="1346" />
                    <RANKING order="7" place="7" resultid="1569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1659" />
                    <RANKING order="2" place="2" resultid="1789" />
                    <RANKING order="3" place="3" resultid="1508" />
                    <RANKING order="4" place="4" resultid="1934" />
                    <RANKING order="5" place="5" resultid="1873" />
                    <RANKING order="6" place="6" resultid="1313" />
                    <RANKING order="7" place="7" resultid="1940" />
                    <RANKING order="8" place="8" resultid="1357" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1353" />
                    <RANKING order="2" place="2" resultid="1665" />
                    <RANKING order="3" place="-1" resultid="1478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1220" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1653" />
                    <RANKING order="2" place="2" resultid="1329" />
                    <RANKING order="3" place="-1" resultid="1424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1221" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1631" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1222" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1439" />
                    <RANKING order="2" place="2" resultid="1923" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1223" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1642" />
                    <RANKING order="2" place="2" resultid="1627" />
                    <RANKING order="3" place="3" resultid="1917" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2026" daytime="17:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2027" daytime="17:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2028" daytime="17:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2029" daytime="17:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2030" daytime="17:24" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1224" daytime="17:28" gender="M" number="36" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1225" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1695" />
                    <RANKING order="2" place="2" resultid="1820" />
                    <RANKING order="3" place="3" resultid="1730" />
                    <RANKING order="4" place="4" resultid="1579" />
                    <RANKING order="5" place="5" resultid="1339" />
                    <RANKING order="6" place="6" resultid="1379" />
                    <RANKING order="7" place="7" resultid="1383" />
                    <RANKING order="8" place="8" resultid="1573" />
                    <RANKING order="9" place="-1" resultid="1958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1226" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1671" />
                    <RANKING order="2" place="2" resultid="1795" />
                    <RANKING order="3" place="3" resultid="1519" />
                    <RANKING order="4" place="4" resultid="1555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1227" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1736" />
                    <RANKING order="2" place="2" resultid="1484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1228" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1636" />
                    <RANKING order="2" place="2" resultid="1801" />
                    <RANKING order="3" place="3" resultid="1748" />
                    <RANKING order="4" place="4" resultid="1332" />
                    <RANKING order="5" place="5" resultid="1502" />
                    <RANKING order="6" place="6" resultid="1490" />
                    <RANKING order="7" place="7" resultid="1433" />
                    <RANKING order="8" place="8" resultid="1911" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1229" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1683" />
                    <RANKING order="2" place="2" resultid="1473" />
                    <RANKING order="3" place="3" resultid="1496" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1461" />
                    <RANKING order="2" place="2" resultid="1928" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1445" />
                    <RANKING order="2" place="2" resultid="1618" />
                    <RANKING order="3" place="3" resultid="1322" />
                    <RANKING order="4" place="4" resultid="1456" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2031" daytime="17:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2032" daytime="17:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2033" daytime="17:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2034" daytime="17:42" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2035" daytime="17:44" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2036" daytime="17:48" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1232" daytime="17:52" gender="F" number="37" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1233" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1406" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2037" daytime="17:52" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1234" daytime="17:54" gender="M" number="38" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1235" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1594" />
                    <RANKING order="2" place="2" resultid="1403" />
                    <RANKING order="3" place="3" resultid="1412" />
                    <RANKING order="4" place="4" resultid="1414" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2038" daytime="17:54" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1236" daytime="18:12" gender="F" number="39" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1237" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1591" />
                    <RANKING order="2" place="2" resultid="1605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1238" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1523" />
                    <RANKING order="2" place="2" resultid="1856" />
                    <RANKING order="3" place="3" resultid="1898" />
                    <RANKING order="4" place="4" resultid="1612" />
                    <RANKING order="5" place="5" resultid="1398" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2039" daytime="18:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2040" daytime="18:14" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1239" daytime="18:16" gender="M" number="40" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1240" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1883" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1878" />
                    <RANKING order="2" place="2" resultid="1888" />
                    <RANKING order="3" place="3" resultid="1602" />
                    <RANKING order="4" place="4" resultid="1609" />
                    <RANKING order="5" place="5" resultid="1583" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2041" daytime="18:16" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1242" daytime="18:20" gender="F" number="41" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1243" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1364" />
                    <RANKING order="2" place="2" resultid="1375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1244" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1839" />
                    <RANKING order="2" place="2" resultid="1598" />
                    <RANKING order="3" place="-1" resultid="1835" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2042" daytime="18:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1245" daytime="18:24" gender="M" number="42" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1246" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1756" />
                    <RANKING order="2" place="-1" resultid="1528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1533" />
                    <RANKING order="2" place="2" resultid="1565" />
                    <RANKING order="3" place="-1" resultid="1418" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2043" daytime="18:24" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1248" daytime="18:26" gender="F" number="43" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1249" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1718" />
                    <RANKING order="2" place="2" resultid="1867" />
                    <RANKING order="3" place="3" resultid="1945" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1250" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1251" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1252" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1706" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1253" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1254" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1255" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2044" daytime="18:26" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1256" daytime="18:30" gender="M" number="44" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1257" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1689" />
                    <RANKING order="2" place="2" resultid="1729" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1258" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1677" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1647" />
                    <RANKING order="2" place="2" resultid="1735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1261" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1472" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1262" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1451" />
                    <RANKING order="2" place="2" resultid="1622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2045" daytime="18:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2046" daytime="18:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1264" daytime="18:40" gender="F" number="45" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1265" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1717" />
                    <RANKING order="2" place="2" resultid="1345" />
                    <RANKING order="3" place="3" resultid="1568" />
                    <RANKING order="4" place="4" resultid="1587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1933" />
                    <RANKING order="2" place="2" resultid="1507" />
                    <RANKING order="3" place="3" resultid="1356" />
                    <RANKING order="4" place="-1" resultid="1939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1267" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1268" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1423" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1269" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1270" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1438" />
                    <RANKING order="2" place="2" resultid="1922" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1271" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1916" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2047" daytime="18:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2048" daytime="18:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2049" daytime="18:46" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1272" daytime="18:48" gender="M" number="46" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1273" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1694" />
                    <RANKING order="2" place="2" resultid="1368" />
                    <RANKING order="3" place="3" resultid="1578" />
                    <RANKING order="4" place="4" resultid="1395" />
                    <RANKING order="5" place="5" resultid="1572" />
                    <RANKING order="6" place="-1" resultid="1957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1274" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1518" />
                    <RANKING order="2" place="2" resultid="1554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1910" />
                    <RANKING order="2" place="2" resultid="1432" />
                    <RANKING order="3" place="3" resultid="1489" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1278" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1460" />
                    <RANKING order="2" place="2" resultid="1742" />
                    <RANKING order="3" place="3" resultid="1450" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1319" />
                    <RANKING order="2" place="2" resultid="1444" />
                    <RANKING order="3" place="3" resultid="1455" />
                    <RANKING order="4" place="4" resultid="1617" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2050" daytime="18:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2051" daytime="18:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2052" daytime="18:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2053" daytime="18:58" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1280" daytime="19:00" gender="F" number="47" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1281" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1386" />
                    <RANKING order="2" place="2" resultid="1825" />
                    <RANKING order="3" place="3" resultid="1902" />
                    <RANKING order="4" place="4" resultid="1590" />
                    <RANKING order="5" place="5" resultid="1604" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1282" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1371" />
                    <RANKING order="2" place="2" resultid="1559" />
                    <RANKING order="3" place="3" resultid="1543" />
                    <RANKING order="4" place="4" resultid="1830" />
                    <RANKING order="5" place="5" resultid="1409" />
                    <RANKING order="6" place="6" resultid="1611" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2054" daytime="19:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2055" daytime="19:02" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1283" daytime="19:04" gender="M" number="48" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1284" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1390" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1777" />
                    <RANKING order="2" place="2" resultid="1548" />
                    <RANKING order="3" place="3" resultid="1766" />
                    <RANKING order="4" place="4" resultid="1601" />
                    <RANKING order="5" place="5" resultid="1349" />
                    <RANKING order="6" place="6" resultid="1582" />
                    <RANKING order="7" place="7" resultid="1608" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2056" daytime="19:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2057" daytime="19:06" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1286" daytime="19:10" gender="F" number="49" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1287" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1893" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1512" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2058" daytime="19:10" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1289" daytime="19:12" gender="M" number="50" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1290" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1538" />
                    <RANKING order="2" place="-1" resultid="1761" />
                    <RANKING order="3" place="-1" resultid="1811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1291" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1861" />
                    <RANKING order="2" place="2" resultid="1700" />
                    <RANKING order="3" place="3" resultid="1564" />
                    <RANKING order="4" place="4" resultid="1806" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2059" daytime="19:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2060" daytime="19:14" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1292" daytime="19:16" gender="F" number="51" order="26" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1293" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1951" />
                    <RANKING order="2" place="2" resultid="1782" />
                    <RANKING order="3" place="3" resultid="1326" />
                    <RANKING order="4" place="4" resultid="1586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1294" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1295" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1296" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1297" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1298" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1437" />
                    <RANKING order="2" place="-1" resultid="1921" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1299" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1641" />
                    <RANKING order="2" place="2" resultid="1915" />
                    <RANKING order="3" place="-1" resultid="1626" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2061" daytime="19:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2062" daytime="19:20" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1300" daytime="19:22" gender="M" number="52" order="27" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1301" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1712" />
                    <RANKING order="2" place="2" resultid="1772" />
                    <RANKING order="3" place="3" resultid="1851" />
                    <RANKING order="4" place="4" resultid="1577" />
                    <RANKING order="5" place="5" resultid="1338" />
                    <RANKING order="6" place="6" resultid="1394" />
                    <RANKING order="7" place="7" resultid="1382" />
                    <RANKING order="8" place="-1" resultid="1956" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1302" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1794" />
                    <RANKING order="2" place="2" resultid="1553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1303" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1304" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1466" />
                    <RANKING order="2" place="2" resultid="1747" />
                    <RANKING order="3" place="3" resultid="1800" />
                    <RANKING order="4" place="4" resultid="1909" />
                    <RANKING order="5" place="5" resultid="1501" />
                    <RANKING order="6" place="6" resultid="1431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1305" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1682" />
                    <RANKING order="2" place="2" resultid="1335" />
                    <RANKING order="3" place="3" resultid="1495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1306" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1927" />
                    <RANKING order="2" place="2" resultid="1342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1307" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2063" daytime="19:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2064" daytime="19:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2065" daytime="19:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2066" daytime="19:30" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="3501" nation="BRA" region="PR" clubid="1309" swrid="93752" name="Ortega &amp; De Souza Jesus" shortname="Aquafoz">
          <ATHLETES>
            <ATHLETE firstname="Emma" lastname="Raquel Nascimento" birthdate="2015-11-06" gender="F" nation="BRA" license="392837" swrid="5641775" athleteid="1384" externalid="392837">
              <RESULTS>
                <RESULT eventid="1156" points="90" swimtime="00:00:54.38" resultid="1385" heatid="2001" lane="4" entrytime="00:00:48.79" entrycourse="SCM" />
                <RESULT eventid="1280" points="144" swimtime="00:00:43.74" resultid="1386" heatid="2055" lane="5" entrytime="00:00:43.96" entrycourse="SCM" />
                <RESULT eventid="1204" points="148" swimtime="00:01:46.77" resultid="1387" heatid="2020" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Wirtti" birthdate="2011-01-14" gender="M" nation="BRA" license="383854" swrid="4917570" athleteid="1365" externalid="383854">
              <RESULTS>
                <RESULT eventid="1176" points="126" swimtime="00:01:35.11" resultid="1366" heatid="2008" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="260" swimtime="00:01:10.23" resultid="1367" heatid="1965" lane="1" entrytime="00:01:15.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="204" swimtime="00:01:22.03" resultid="1368" heatid="2051" lane="2" entrytime="00:01:29.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Varela" birthdate="2010-05-20" gender="F" nation="BRA" license="365503" swrid="5596942" athleteid="1354" externalid="365503">
              <RESULTS>
                <RESULT eventid="1140" points="213" swimtime="00:03:19.08" resultid="1355" heatid="1998" lane="1" entrytime="00:03:22.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.62" />
                    <SPLIT distance="100" swimtime="00:01:37.27" />
                    <SPLIT distance="150" swimtime="00:02:29.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="243" swimtime="00:01:27.96" resultid="1356" heatid="2048" lane="3" entrytime="00:01:31.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="239" swimtime="00:02:57.64" resultid="1357" heatid="2027" lane="2" entrytime="00:03:06.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.34" />
                    <SPLIT distance="100" swimtime="00:01:27.88" />
                    <SPLIT distance="150" swimtime="00:02:15.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="De Zanchet" birthdate="2015-09-16" gender="M" nation="BRA" license="392838" swrid="5641762" athleteid="1388" externalid="392838">
              <RESULTS>
                <RESULT eventid="1115" points="106" swimtime="00:00:52.63" resultid="1389" heatid="1986" lane="2" entrytime="00:00:55.70" entrycourse="SCM" />
                <RESULT eventid="1283" points="89" swimtime="00:00:45.10" resultid="1390" heatid="2056" lane="4" />
                <RESULT eventid="1207" points="75" swimtime="00:01:56.58" resultid="1391" heatid="2021" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Marques Lima" birthdate="2010-04-30" gender="F" nation="BRA" license="383051" swrid="5596913" athleteid="1358" externalid="383051">
              <RESULTS>
                <RESULT eventid="1168" points="200" swimtime="00:01:32.29" resultid="1359" heatid="2006" lane="5" entrytime="00:01:28.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="304" swimtime="00:02:56.70" resultid="1360" heatid="1997" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                    <SPLIT distance="100" swimtime="00:01:25.59" />
                    <SPLIT distance="150" swimtime="00:02:11.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="299" swimtime="00:01:15.10" resultid="1361" heatid="1960" lane="4" entrytime="00:01:20.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isis" lastname="Lukianou Souza" birthdate="2016-09-28" gender="F" nation="BRA" license="406655" athleteid="1404" externalid="406655">
              <RESULTS>
                <RESULT eventid="1108" points="18" swimtime="00:01:34.78" resultid="1405" heatid="1981" lane="3" />
                <RESULT eventid="1232" points="22" swimtime="00:01:21.79" resultid="1406" heatid="2037" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alejandro" lastname="Manuel Melgarejo" birthdate="2016-04-28" gender="M" nation="BRA" license="407315" athleteid="1410" externalid="407315">
              <RESULTS>
                <RESULT eventid="1110" points="42" swimtime="00:01:03.55" resultid="1411" heatid="1982" lane="2" />
                <RESULT eventid="1234" points="36" swimtime="00:01:00.92" resultid="1412" heatid="2038" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Pires" birthdate="2011-04-09" gender="F" nation="BRA" license="383853" swrid="5596927" athleteid="1323" externalid="383853">
              <RESULTS>
                <RESULT eventid="1092" points="193" swimtime="00:03:52.64" resultid="1324" heatid="1975" lane="4" entrytime="00:04:16.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.33" />
                    <SPLIT distance="100" swimtime="00:01:53.41" />
                    <SPLIT distance="150" swimtime="00:02:53.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="192" swimtime="00:01:27.05" resultid="1325" heatid="1960" lane="5" entrytime="00:01:30.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="201" swimtime="00:01:46.33" resultid="1326" heatid="2061" lane="4" entrytime="00:01:48.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julio" lastname="Heck" birthdate="1998-02-15" gender="M" nation="BRA" license="185880" swrid="5596906" athleteid="1320" externalid="185880">
              <RESULTS>
                <RESULT eventid="1068" points="481" swimtime="00:00:57.21" resultid="1321" heatid="1968" lane="3" entrytime="00:00:52.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="386" swimtime="00:02:16.40" resultid="1322" heatid="2035" lane="2" entrytime="00:02:08.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                    <SPLIT distance="100" swimtime="00:01:05.49" />
                    <SPLIT distance="150" swimtime="00:01:42.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Xavier" birthdate="2011-10-14" gender="M" nation="BRA" license="370564" swrid="5596949" athleteid="1336" externalid="370564">
              <RESULTS>
                <RESULT eventid="1100" points="209" swimtime="00:03:22.23" resultid="1337" heatid="1978" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.04" />
                    <SPLIT distance="100" swimtime="00:01:36.84" />
                    <SPLIT distance="150" swimtime="00:02:29.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="202" swimtime="00:01:34.20" resultid="1338" heatid="2064" lane="4" entrytime="00:01:41.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="168" swimtime="00:03:00.03" resultid="1339" heatid="2032" lane="3" entrytime="00:03:10.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.43" />
                    <SPLIT distance="100" swimtime="00:01:28.16" />
                    <SPLIT distance="150" swimtime="00:02:15.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Afonso Proteti" birthdate="2002-03-19" gender="M" nation="BRA" license="190464" swrid="5596865" athleteid="1317" externalid="190464">
              <RESULTS>
                <RESULT eventid="1176" points="593" swimtime="00:00:56.84" resultid="1318" heatid="2010" lane="3" entrytime="00:00:55.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="544" swimtime="00:00:59.17" resultid="1319" heatid="2053" lane="3" entrytime="00:00:57.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Voltolini" birthdate="2014-06-29" gender="M" nation="BRA" license="383846" swrid="5596947" athleteid="1347" externalid="383846">
              <RESULTS>
                <RESULT eventid="1115" points="85" swimtime="00:00:56.71" resultid="1348" heatid="1986" lane="5" entrytime="00:00:57.31" entrycourse="SCM" />
                <RESULT eventid="1283" points="74" swimtime="00:00:47.84" resultid="1349" heatid="2057" lane="5" entrytime="00:00:44.07" entrycourse="SCM" />
                <RESULT eventid="1207" points="73" swimtime="00:01:57.54" resultid="1350" heatid="2021" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Otremba Rouver" birthdate="2007-04-25" gender="M" nation="BRA" license="342152" swrid="5596919" athleteid="1333" externalid="342152">
              <RESULTS>
                <RESULT eventid="1176" points="400" swimtime="00:01:04.80" resultid="1334" heatid="2008" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="401" swimtime="00:01:14.95" resultid="1335" heatid="2064" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Mussi" birthdate="2006-12-31" gender="M" nation="BRA" license="370567" swrid="5596917" athleteid="1340" externalid="370567">
              <RESULTS>
                <RESULT eventid="1100" points="289" swimtime="00:03:01.63" resultid="1341" heatid="1980" lane="1" entrytime="00:02:47.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.28" />
                    <SPLIT distance="100" swimtime="00:01:25.87" />
                    <SPLIT distance="150" swimtime="00:02:13.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="369" swimtime="00:01:17.01" resultid="1342" heatid="2066" lane="2" entrytime="00:01:12.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Franco" birthdate="2010-06-09" gender="F" nation="BRA" license="383849" swrid="5596896" athleteid="1310" externalid="383849">
              <RESULTS>
                <RESULT eventid="1168" points="232" swimtime="00:01:27.91" resultid="1311" heatid="2006" lane="2" entrytime="00:01:25.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="334" swimtime="00:01:12.40" resultid="1312" heatid="1961" lane="1" entrytime="00:01:12.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="294" swimtime="00:02:45.86" resultid="1313" heatid="2028" lane="5" entrytime="00:02:39.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:19.61" />
                    <SPLIT distance="150" swimtime="00:02:03.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Mendes Portela" birthdate="2014-03-08" gender="F" nation="BRA" license="406656" swrid="5117156" athleteid="1407" externalid="406656">
              <RESULTS>
                <RESULT eventid="1112" points="60" swimtime="00:01:12.22" resultid="1408" heatid="1983" lane="4" entrytime="00:01:21.00" entrycourse="SCM" />
                <RESULT eventid="1280" points="78" swimtime="00:00:53.55" resultid="1409" heatid="2054" lane="2" entrytime="00:01:01.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Garcete" birthdate="2014-01-04" gender="F" nation="BRA" license="383856" swrid="5596904" athleteid="1369" externalid="383856">
              <RESULTS>
                <RESULT eventid="1156" points="163" swimtime="00:00:44.62" resultid="1370" heatid="2001" lane="3" entrytime="00:00:45.40" entrycourse="SCM" />
                <RESULT eventid="1280" points="182" swimtime="00:00:40.41" resultid="1371" heatid="2055" lane="3" entrytime="00:00:40.95" entrycourse="SCM" />
                <RESULT eventid="1204" points="137" swimtime="00:01:49.58" resultid="1372" heatid="2020" lane="4" entrytime="00:01:53.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauan" lastname="Matheus Cunha" birthdate="2011-01-31" gender="M" nation="BRA" license="392834" swrid="5641770" athleteid="1376" externalid="392834">
              <RESULTS>
                <RESULT eventid="1176" points="89" swimtime="00:01:46.74" resultid="1377" heatid="2008" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="161" swimtime="00:01:22.39" resultid="1378" heatid="1964" lane="2" entrytime="00:01:28.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="164" swimtime="00:03:01.26" resultid="1379" heatid="2032" lane="2" entrytime="00:03:21.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                    <SPLIT distance="100" swimtime="00:01:28.63" />
                    <SPLIT distance="150" swimtime="00:02:15.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Dominguez Olivieski" birthdate="2011-04-27" gender="M" nation="BRA" license="405717" swrid="5664737" athleteid="1392" externalid="405717">
              <RESULTS>
                <RESULT eventid="1068" points="163" swimtime="00:01:21.97" resultid="1393" heatid="1964" lane="4" entrytime="00:01:23.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="168" swimtime="00:01:40.03" resultid="1394" heatid="2064" lane="2" entrytime="00:01:50.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="154" swimtime="00:01:29.99" resultid="1395" heatid="2051" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Helena Sousa" birthdate="2013-03-20" gender="F" nation="BRA" license="392832" swrid="5641765" athleteid="1373" externalid="392832">
              <RESULTS>
                <RESULT eventid="1118" points="155" swimtime="00:01:33.42" resultid="1374" heatid="1987" lane="4" entrytime="00:01:34.67" entrycourse="SCM" />
                <RESULT eventid="1242" points="128" swimtime="00:01:48.87" resultid="1375" heatid="2042" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Rorato" birthdate="2013-04-18" gender="F" nation="BRA" license="383851" swrid="5596936" athleteid="1362" externalid="383851">
              <RESULTS>
                <RESULT eventid="1162" points="165" swimtime="00:00:44.38" resultid="1363" heatid="2003" lane="3" entrytime="00:00:42.19" entrycourse="SCM" />
                <RESULT eventid="1242" points="190" swimtime="00:01:35.44" resultid="1364" heatid="2042" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Gustavo Cunha" birthdate="2011-01-31" gender="M" nation="BRA" license="392836" swrid="5641764" athleteid="1380" externalid="392836">
              <RESULTS>
                <RESULT eventid="1100" points="164" swimtime="00:03:39.35" resultid="1381" heatid="1978" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.87" />
                    <SPLIT distance="100" swimtime="00:01:46.51" />
                    <SPLIT distance="150" swimtime="00:02:42.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="147" swimtime="00:01:44.54" resultid="1382" heatid="2064" lane="5" entrytime="00:01:52.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="163" swimtime="00:03:01.68" resultid="1383" heatid="2032" lane="4" entrytime="00:03:11.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.12" />
                    <SPLIT distance="100" swimtime="00:01:30.18" />
                    <SPLIT distance="150" swimtime="00:02:17.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ian" lastname="Peroni Ottomar" birthdate="2016-07-15" gender="M" nation="BRA" license="406653" swrid="5258754" athleteid="1401" externalid="406653">
              <RESULTS>
                <RESULT eventid="1110" points="60" swimtime="00:00:56.20" resultid="1402" heatid="1982" lane="3" />
                <RESULT eventid="1234" points="44" swimtime="00:00:56.82" resultid="1403" heatid="2038" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="De Albuquerque" birthdate="2014-11-19" gender="F" nation="BRA" license="406648" swrid="4823632" athleteid="1396" externalid="406648">
              <RESULTS>
                <RESULT eventid="1112" points="39" swimtime="00:01:23.17" resultid="1397" heatid="1983" lane="2" entrytime="00:01:28.90" entrycourse="SCM" />
                <RESULT eventid="1236" points="32" swimtime="00:01:19.41" resultid="1398" heatid="2040" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo" lastname="Antonio Sousa" birthdate="2012-03-17" gender="M" nation="BRA" license="407497" athleteid="1416" externalid="407497">
              <RESULTS>
                <RESULT eventid="1121" status="DSQ" swimtime="00:00:00.00" resultid="1417" heatid="1988" lane="4" />
                <RESULT eventid="1245" status="DSQ" swimtime="00:01:56.72" resultid="1418" heatid="2043" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Geórgia" lastname="Adeli Jesus" birthdate="2008-03-27" gender="F" nation="BRA" license="312649" swrid="5596864" athleteid="1327" externalid="312649">
              <RESULTS>
                <RESULT eventid="1124" points="384" swimtime="00:10:56.73" resultid="1328" heatid="1991" lane="3" entrytime="00:11:16.95" entrycourse="SCM" />
                <RESULT eventid="1216" points="401" swimtime="00:02:29.51" resultid="1329" heatid="2029" lane="4" entrytime="00:02:31.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.21" />
                    <SPLIT distance="150" swimtime="00:01:52.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Marques Voltolini" birthdate="2016-04-25" gender="M" nation="BRA" license="407316" athleteid="1413" externalid="407316">
              <RESULTS>
                <RESULT eventid="1234" points="22" swimtime="00:01:11.56" resultid="1414" heatid="2038" lane="4" />
                <RESULT eventid="1202" points="38" swimtime="00:01:13.69" resultid="1415" heatid="2018" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Maguet" birthdate="2011-07-01" gender="F" nation="BRA" license="370568" swrid="5596911" athleteid="1343" externalid="370568">
              <RESULTS>
                <RESULT eventid="1060" points="242" swimtime="00:01:20.57" resultid="1344" heatid="1960" lane="2" entrytime="00:01:22.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="182" swimtime="00:01:36.83" resultid="1345" heatid="2048" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="236" swimtime="00:02:58.48" resultid="1346" heatid="2027" lane="5" entrytime="00:03:06.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                    <SPLIT distance="100" swimtime="00:01:27.48" />
                    <SPLIT distance="150" swimtime="00:02:14.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Victoria Portela" birthdate="2009-12-04" gender="F" nation="BRA" license="383047" swrid="5596945" athleteid="1351" externalid="383047">
              <RESULTS>
                <RESULT eventid="1060" points="423" swimtime="00:01:06.90" resultid="1352" heatid="1962" lane="2" entrytime="00:01:07.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="398" swimtime="00:02:29.90" resultid="1353" heatid="2029" lane="2" entrytime="00:02:32.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:13.51" />
                    <SPLIT distance="150" swimtime="00:01:52.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Gabriel Serighelli" birthdate="1999-03-12" gender="M" nation="BRA" license="121253" swrid="5596899" athleteid="1314" externalid="121253">
              <RESULTS>
                <RESULT eventid="1176" points="450" swimtime="00:01:02.31" resultid="1315" heatid="2010" lane="4" entrytime="00:00:59.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="467" swimtime="00:00:57.77" resultid="1316" heatid="1968" lane="4" entrytime="00:00:53.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yago" lastname="Simon Pires" birthdate="2008-10-29" gender="M" nation="BRA" license="328942" swrid="5596939" athleteid="1330" externalid="328942">
              <RESULTS>
                <RESULT eventid="1068" points="429" swimtime="00:00:59.41" resultid="1331" heatid="1967" lane="4" entrytime="00:00:59.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="441" swimtime="00:02:10.50" resultid="1332" heatid="2031" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                    <SPLIT distance="100" swimtime="00:01:02.57" />
                    <SPLIT distance="150" swimtime="00:01:36.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Miguel Bogado" birthdate="2013-05-28" gender="M" nation="PRY" license="406649" athleteid="1399" externalid="406649">
              <RESULTS>
                <RESULT eventid="1121" points="40" swimtime="00:02:10.44" resultid="1400" heatid="1988" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3133" nation="BRA" region="PR" clubid="1904" swrid="93768" name="Associação Toledo Natação" shortname="Toledo Natação">
          <ATHLETES>
            <ATHLETE firstname="Isadora" lastname="Marafon" birthdate="2011-03-23" gender="F" nation="BRA" license="380287" swrid="5652623" athleteid="1947" externalid="380287">
              <RESULTS>
                <RESULT eventid="1168" points="164" swimtime="00:01:38.72" resultid="1948" heatid="2005" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" status="DSQ" swimtime="00:03:07.28" resultid="1949" heatid="1975" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                    <SPLIT distance="100" swimtime="00:01:27.18" />
                    <SPLIT distance="150" swimtime="00:02:17.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="406" swimtime="00:01:07.84" resultid="1950" heatid="1961" lane="2" entrytime="00:01:10.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="397" swimtime="00:01:24.84" resultid="1951" heatid="2062" lane="2" entrytime="00:01:27.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="410" swimtime="00:02:28.47" resultid="1952" heatid="2026" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                    <SPLIT distance="100" swimtime="00:01:10.93" />
                    <SPLIT distance="150" swimtime="00:01:49.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Fernando Braga Da Silva" birthdate="2011-01-10" gender="M" nation="BRA" license="380291" swrid="5453344" athleteid="1953" externalid="380291">
              <RESULTS>
                <RESULT eventid="1100" status="DNS" swimtime="00:00:00.00" resultid="1954" heatid="1978" lane="5" />
                <RESULT eventid="1068" status="DNS" swimtime="00:00:00.00" resultid="1955" heatid="1964" lane="3" entrytime="00:01:17.56" entrycourse="SCM" />
                <RESULT eventid="1300" status="DNS" swimtime="00:00:00.00" resultid="1956" heatid="2063" lane="3" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="1957" heatid="2050" lane="4" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="1958" heatid="2033" lane="6" entrytime="00:02:54.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Welter Levandowski" birthdate="2011-05-06" gender="F" nation="BRA" license="380286" swrid="5652626" athleteid="1941" externalid="380286">
              <RESULTS>
                <RESULT eventid="1168" points="241" swimtime="00:01:26.75" resultid="1942" heatid="2006" lane="6" entrytime="00:01:33.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="314" swimtime="00:11:41.77" resultid="1943" heatid="1990" lane="1" />
                <RESULT eventid="1060" status="DSQ" swimtime="00:01:10.77" resultid="1944" heatid="1959" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="236" swimtime="00:03:13.39" resultid="1945" heatid="2044" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                    <SPLIT distance="100" swimtime="00:01:32.19" />
                    <SPLIT distance="150" swimtime="00:02:23.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="373" swimtime="00:02:33.18" resultid="1946" heatid="2028" lane="2" entrytime="00:02:37.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                    <SPLIT distance="150" swimtime="00:01:53.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lavinia" lastname="Martins Paludo" birthdate="2010-09-30" gender="F" nation="BRA" license="347217" swrid="5652624" athleteid="1935" externalid="347217">
              <RESULTS>
                <RESULT eventid="1092" points="264" swimtime="00:03:29.58" resultid="1936" heatid="1975" lane="3" entrytime="00:03:38.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.40" />
                    <SPLIT distance="100" swimtime="00:01:41.35" />
                    <SPLIT distance="150" swimtime="00:02:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="251" swimtime="00:01:19.64" resultid="1937" heatid="1960" lane="3" entrytime="00:01:15.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="246" swimtime="00:01:39.47" resultid="1938" heatid="2061" lane="3" entrytime="00:01:38.23" entrycourse="SCM" />
                <RESULT eventid="1264" status="DNS" swimtime="00:00:00.00" resultid="1939" heatid="2048" lane="4" />
                <RESULT eventid="1216" points="271" swimtime="00:02:50.43" resultid="1940" heatid="2027" lane="3" entrytime="00:02:47.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                    <SPLIT distance="100" swimtime="00:01:20.55" />
                    <SPLIT distance="150" swimtime="00:02:06.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrielly" lastname="Luiza Horn" birthdate="2004-04-03" gender="F" nation="BRA" license="315145" swrid="5622288" athleteid="1912" externalid="315145">
              <RESULTS>
                <RESULT eventid="1168" points="303" swimtime="00:01:20.40" resultid="1913" heatid="2005" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="342" swimtime="00:01:11.79" resultid="1914" heatid="1961" lane="5" entrytime="00:01:12.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="326" swimtime="00:01:30.55" resultid="1915" heatid="2061" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="270" swimtime="00:01:24.90" resultid="1916" heatid="2047" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="289" swimtime="00:02:46.83" resultid="1917" heatid="2027" lane="4" entrytime="00:02:50.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                    <SPLIT distance="100" swimtime="00:01:17.01" />
                    <SPLIT distance="150" swimtime="00:02:02.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Marafon" birthdate="2006-06-17" gender="M" nation="BRA" license="380288" swrid="5622291" athleteid="1924" externalid="380288">
              <RESULTS>
                <RESULT eventid="1100" points="407" swimtime="00:02:42.03" resultid="1925" heatid="1980" lane="5" entrytime="00:02:45.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                    <SPLIT distance="100" swimtime="00:01:18.80" />
                    <SPLIT distance="150" swimtime="00:02:01.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="426" swimtime="00:00:59.58" resultid="1926" heatid="1967" lane="1" entrytime="00:01:00.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="469" swimtime="00:01:11.10" resultid="1927" heatid="2066" lane="3" entrytime="00:01:11.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="316" swimtime="00:02:25.76" resultid="1928" heatid="2031" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:10.27" />
                    <SPLIT distance="150" swimtime="00:01:47.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Feder" birthdate="2008-11-13" gender="M" nation="BRA" license="347224" swrid="5622278" athleteid="1905" externalid="347224">
              <RESULTS>
                <RESULT eventid="1176" points="309" swimtime="00:01:10.64" resultid="1906" heatid="2008" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="363" swimtime="00:02:28.03" resultid="1907" heatid="2000" lane="1" entrytime="00:02:29.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                    <SPLIT distance="100" swimtime="00:01:11.44" />
                    <SPLIT distance="150" swimtime="00:01:50.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="423" swimtime="00:00:59.71" resultid="1908" heatid="1967" lane="5" entrytime="00:00:59.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="273" swimtime="00:01:25.19" resultid="1909" heatid="2063" lane="5" />
                <RESULT eventid="1272" points="381" swimtime="00:01:06.62" resultid="1910" heatid="2053" lane="1" entrytime="00:01:05.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="298" swimtime="00:02:28.75" resultid="1911" heatid="2035" lane="6" entrytime="00:02:16.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:10.46" />
                    <SPLIT distance="150" swimtime="00:01:49.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Torres Romancini" birthdate="2010-05-28" gender="F" nation="BRA" license="347218" swrid="5622309" athleteid="1929" externalid="347218">
              <RESULTS>
                <RESULT eventid="1168" points="241" swimtime="00:01:26.85" resultid="1930" heatid="2005" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="351" swimtime="00:02:48.51" resultid="1931" heatid="1997" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.97" />
                    <SPLIT distance="100" swimtime="00:01:21.09" />
                    <SPLIT distance="150" swimtime="00:02:05.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="336" swimtime="00:01:12.27" resultid="1932" heatid="1959" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="344" swimtime="00:01:18.31" resultid="1933" heatid="2049" lane="5" entrytime="00:01:17.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="336" swimtime="00:02:38.52" resultid="1934" heatid="2026" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:15.08" />
                    <SPLIT distance="150" swimtime="00:01:57.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giullia" lastname="Lagni" birthdate="2006-11-22" gender="F" nation="BRA" license="337671" swrid="5622285" athleteid="1918" externalid="337671">
              <RESULTS>
                <RESULT eventid="1140" points="334" swimtime="00:02:51.27" resultid="1919" heatid="1997" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                    <SPLIT distance="100" swimtime="00:01:21.17" />
                    <SPLIT distance="150" swimtime="00:02:06.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="346" swimtime="00:01:11.56" resultid="1920" heatid="1962" lane="6" entrytime="00:01:09.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" status="DNS" swimtime="00:00:00.00" resultid="1921" heatid="2061" lane="1" />
                <RESULT eventid="1264" points="325" swimtime="00:01:19.83" resultid="1922" heatid="2049" lane="2" entrytime="00:01:16.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="384" swimtime="00:02:31.67" resultid="1923" heatid="2029" lane="6" entrytime="00:02:33.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="100" swimtime="00:01:12.43" />
                    <SPLIT distance="150" swimtime="00:01:52.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="36" nation="BRA" region="PR" clubid="1613" swrid="93753" name="Associação Atlética Comercial" shortname="Comercial Cascavel">
          <ATHLETES>
            <ATHLETE firstname="Isabelle" lastname="Cordeiro Silva" birthdate="2015-06-14" gender="F" nation="BRA" license="390839" swrid="5596878" athleteid="1822" externalid="390839">
              <RESULTS>
                <RESULT eventid="1156" points="96" swimtime="00:00:53.12" resultid="1823" heatid="2001" lane="1" entrytime="00:00:54.05" entrycourse="SCM" />
                <RESULT eventid="1080" points="141" swimtime="00:03:31.57" resultid="1824" heatid="1969" lane="4" />
                <RESULT eventid="1280" points="128" swimtime="00:00:45.44" resultid="1825" heatid="2054" lane="3" entrytime="00:00:45.93" entrycourse="SCM" />
                <RESULT eventid="1204" points="140" swimtime="00:01:48.64" resultid="1826" heatid="2020" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Paese Worm" birthdate="2014-07-23" gender="F" nation="BRA" license="380655" swrid="5596920" athleteid="1750" externalid="380655">
              <RESULTS>
                <RESULT eventid="1112" points="130" swimtime="00:00:55.99" resultid="1751" heatid="1984" lane="2" entrytime="00:00:59.59" entrycourse="SCM" />
                <RESULT eventid="1080" points="167" swimtime="00:03:19.99" resultid="1752" heatid="1969" lane="3" entrytime="00:03:43.28" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Stein Duarte" birthdate="2010-10-03" gender="F" nation="BRA" license="351635" swrid="5588923" athleteid="1655" externalid="351635">
              <RESULTS>
                <RESULT eventid="1140" points="400" swimtime="00:02:41.42" resultid="1656" heatid="1998" lane="4" entrytime="00:02:46.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                    <SPLIT distance="100" swimtime="00:01:18.15" />
                    <SPLIT distance="150" swimtime="00:02:00.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="435" swimtime="00:10:29.97" resultid="1657" heatid="1992" lane="5" entrytime="00:10:35.09" entrycourse="SCM" />
                <RESULT eventid="1092" points="377" swimtime="00:03:06.13" resultid="1658" heatid="1976" lane="5" entrytime="00:03:08.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.69" />
                    <SPLIT distance="100" swimtime="00:01:30.42" />
                    <SPLIT distance="150" swimtime="00:02:18.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="431" swimtime="00:02:26.00" resultid="1659" heatid="2030" lane="6" entrytime="00:02:30.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                    <SPLIT distance="100" swimtime="00:01:11.41" />
                    <SPLIT distance="150" swimtime="00:01:49.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="442" swimtime="00:05:39.75" resultid="1660" heatid="2013" lane="2" entrytime="00:05:44.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:22.29" />
                    <SPLIT distance="150" swimtime="00:02:03.80" />
                    <SPLIT distance="200" swimtime="00:02:43.59" />
                    <SPLIT distance="250" swimtime="00:03:31.94" />
                    <SPLIT distance="300" swimtime="00:04:20.77" />
                    <SPLIT distance="350" swimtime="00:05:00.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Vieira Rohnelt" birthdate="2012-05-03" gender="M" nation="BRA" license="365692" swrid="5588952" athleteid="1697" externalid="365692">
              <RESULTS>
                <RESULT eventid="1165" points="117" swimtime="00:00:44.38" resultid="1698" heatid="2004" lane="2" entrytime="00:00:44.49" entrycourse="SCM" />
                <RESULT eventid="1089" points="185" swimtime="00:03:12.33" resultid="1699" heatid="1974" lane="5" entrytime="00:03:14.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.80" />
                    <SPLIT distance="100" swimtime="00:01:32.28" />
                    <SPLIT distance="150" swimtime="00:02:28.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="131" swimtime="00:00:49.03" resultid="1700" heatid="2060" lane="2" entrytime="00:00:48.53" entrycourse="SCM" />
                <RESULT eventid="1213" points="193" swimtime="00:06:06.80" resultid="1701" heatid="2025" lane="2" entrytime="00:06:30.77" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hendrik" lastname="Alteiro Groenwold" birthdate="2011-03-23" gender="M" nation="BRA" license="365756" swrid="5588520" athleteid="1685" externalid="365756">
              <RESULTS>
                <RESULT eventid="1176" points="304" swimtime="00:01:11.00" resultid="1686" heatid="2009" lane="2" entrytime="00:01:10.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="354" swimtime="00:10:26.41" resultid="1687" heatid="1995" lane="4" />
                <RESULT eventid="1068" points="341" swimtime="00:01:04.15" resultid="1688" heatid="1966" lane="1" entrytime="00:01:04.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="282" swimtime="00:02:42.93" resultid="1689" heatid="2045" lane="4" entrytime="00:02:54.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                    <SPLIT distance="100" swimtime="00:01:18.05" />
                    <SPLIT distance="150" swimtime="00:02:00.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" status="DSQ" swimtime="00:05:38.67" resultid="1690" heatid="2015" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:18.07" />
                    <SPLIT distance="150" swimtime="00:01:59.95" />
                    <SPLIT distance="200" swimtime="00:02:41.07" />
                    <SPLIT distance="250" swimtime="00:03:31.47" />
                    <SPLIT distance="300" swimtime="00:04:22.81" />
                    <SPLIT distance="350" swimtime="00:05:01.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Borille Busetti" birthdate="2010-02-17" gender="F" nation="BRA" license="392830" swrid="5622263" athleteid="1869" externalid="392830">
              <RESULTS>
                <RESULT eventid="1140" points="235" swimtime="00:03:12.73" resultid="1870" heatid="1997" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.65" />
                    <SPLIT distance="100" swimtime="00:01:31.65" />
                    <SPLIT distance="150" swimtime="00:02:22.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="261" swimtime="00:12:26.37" resultid="1871" heatid="1991" lane="5" />
                <RESULT eventid="1092" status="DSQ" swimtime="00:03:42.54" resultid="1872" heatid="1975" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.90" />
                    <SPLIT distance="100" swimtime="00:01:47.42" />
                    <SPLIT distance="150" swimtime="00:02:45.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="304" swimtime="00:02:44.04" resultid="1873" heatid="2028" lane="6" entrytime="00:02:44.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                    <SPLIT distance="100" swimtime="00:01:21.10" />
                    <SPLIT distance="150" swimtime="00:02:04.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="219" swimtime="00:07:09.35" resultid="1874" heatid="2012" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.06" />
                    <SPLIT distance="100" swimtime="00:01:44.82" />
                    <SPLIT distance="150" swimtime="00:02:39.57" />
                    <SPLIT distance="200" swimtime="00:03:34.51" />
                    <SPLIT distance="250" swimtime="00:04:35.56" />
                    <SPLIT distance="300" swimtime="00:05:36.95" />
                    <SPLIT distance="350" swimtime="00:06:25.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Macedo Medeiros" birthdate="2012-05-12" gender="M" nation="BRA" license="392015" swrid="4697574" athleteid="1858" externalid="392015">
              <RESULTS>
                <RESULT eventid="1165" points="95" swimtime="00:00:47.59" resultid="1859" heatid="2004" lane="1" entrytime="00:01:04.81" entrycourse="SCM" />
                <RESULT eventid="1089" status="DSQ" swimtime="00:03:32.23" resultid="1860" heatid="1973" lane="3" entrytime="00:03:46.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.20" />
                    <SPLIT distance="100" swimtime="00:01:43.45" />
                    <SPLIT distance="150" swimtime="00:02:40.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="132" swimtime="00:00:48.99" resultid="1861" heatid="2059" lane="2" entrytime="00:00:55.56" entrycourse="SCM" />
                <RESULT eventid="1213" points="146" swimtime="00:06:42.50" resultid="1862" heatid="2024" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raul" lastname="Bonamigo" birthdate="2010-12-01" gender="M" nation="BRA" license="344397" swrid="5588559" athleteid="1791" externalid="344397">
              <RESULTS>
                <RESULT eventid="1132" points="388" swimtime="00:10:07.60" resultid="1792" heatid="1996" lane="1" entrytime="00:10:01.23" entrycourse="SCM" />
                <RESULT eventid="1100" points="296" swimtime="00:03:00.29" resultid="1793" heatid="1979" lane="1" entrytime="00:03:17.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                    <SPLIT distance="100" swimtime="00:01:25.58" />
                    <SPLIT distance="150" swimtime="00:02:13.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="278" swimtime="00:01:24.60" resultid="1794" heatid="2065" lane="2" entrytime="00:01:26.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="357" swimtime="00:02:19.96" resultid="1795" heatid="2033" lane="5" entrytime="00:02:28.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="100" swimtime="00:01:07.31" />
                    <SPLIT distance="150" swimtime="00:01:43.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="332" swimtime="00:05:38.81" resultid="1796" heatid="2016" lane="4" entrytime="00:05:26.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                    <SPLIT distance="100" swimtime="00:01:20.37" />
                    <SPLIT distance="150" swimtime="00:02:03.18" />
                    <SPLIT distance="200" swimtime="00:02:44.08" />
                    <SPLIT distance="250" swimtime="00:03:33.28" />
                    <SPLIT distance="300" swimtime="00:04:22.38" />
                    <SPLIT distance="350" swimtime="00:05:01.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Bonamigo" birthdate="2013-06-25" gender="M" nation="BRA" license="365484" swrid="5588558" athleteid="1808" externalid="365484">
              <RESULTS>
                <RESULT eventid="1121" status="DNS" swimtime="00:00:00.00" resultid="1809" heatid="1989" lane="3" entrytime="00:01:14.92" entrycourse="SCM" />
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="1810" heatid="1974" lane="4" entrytime="00:03:07.13" entrycourse="SCM" />
                <RESULT eventid="1289" status="DNS" swimtime="00:00:00.00" resultid="1811" heatid="2060" lane="3" entrytime="00:00:41.58" entrycourse="SCM" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="1812" heatid="2025" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Bezerra Sedlacek" birthdate="2014-02-26" gender="M" nation="BRA" license="380663" swrid="4300166" athleteid="1763" externalid="380663">
              <RESULTS>
                <RESULT eventid="1115" points="108" swimtime="00:00:52.39" resultid="1764" heatid="1986" lane="4" entrytime="00:00:52.58" entrycourse="SCM" />
                <RESULT eventid="1083" points="122" swimtime="00:03:19.91" resultid="1765" heatid="1971" lane="5" entrytime="00:03:33.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                    <SPLIT distance="100" swimtime="00:01:34.61" />
                    <SPLIT distance="150" swimtime="00:02:26.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" points="109" swimtime="00:00:42.08" resultid="1766" heatid="2057" lane="2" entrytime="00:00:42.09" entrycourse="SCM" />
                <RESULT eventid="1207" points="106" swimtime="00:01:44.11" resultid="1767" heatid="2022" lane="2" entrytime="00:01:59.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Rinaldini" birthdate="2009-04-09" gender="M" nation="BRA" license="348289" swrid="5596932" athleteid="1643" externalid="348289">
              <RESULTS>
                <RESULT eventid="1176" points="419" swimtime="00:01:03.83" resultid="1644" heatid="2009" lane="3" entrytime="00:01:05.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="550" swimtime="00:09:00.95" resultid="1645" heatid="1995" lane="2" />
                <RESULT eventid="1068" points="437" swimtime="00:00:59.05" resultid="1646" heatid="1963" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="485" swimtime="00:02:15.99" resultid="1647" heatid="2046" lane="2" entrytime="00:02:19.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:04.56" />
                    <SPLIT distance="150" swimtime="00:01:40.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="493" swimtime="00:04:57.20" resultid="1648" heatid="2017" lane="1" entrytime="00:05:03.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                    <SPLIT distance="100" swimtime="00:01:07.37" />
                    <SPLIT distance="150" swimtime="00:01:46.20" />
                    <SPLIT distance="200" swimtime="00:02:24.22" />
                    <SPLIT distance="250" swimtime="00:03:08.55" />
                    <SPLIT distance="300" swimtime="00:03:52.85" />
                    <SPLIT distance="350" swimtime="00:04:26.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose" lastname="Eliziario Filho" birthdate="2014-03-27" gender="M" nation="BRA" license="406696" swrid="4979701" athleteid="1885" externalid="406696">
              <RESULTS>
                <RESULT eventid="1159" points="90" swimtime="00:00:48.42" resultid="1886" heatid="2002" lane="4" entrytime="00:00:48.90" entrycourse="SCM" />
                <RESULT eventid="1083" points="115" swimtime="00:03:23.99" resultid="1887" heatid="1971" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.13" />
                    <SPLIT distance="100" swimtime="00:01:36.66" />
                    <SPLIT distance="150" swimtime="00:02:32.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="75" swimtime="00:00:52.21" resultid="1888" heatid="2041" lane="4" entrytime="00:00:56.64" entrycourse="SCM" />
                <RESULT eventid="1207" points="96" swimtime="00:01:47.33" resultid="1889" heatid="2021" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Gaio" birthdate="2014-08-27" gender="F" nation="BRA" license="390841" swrid="5596900" athleteid="1827" externalid="390841">
              <RESULTS>
                <RESULT eventid="1112" points="113" swimtime="00:00:58.52" resultid="1828" heatid="1984" lane="4" entrytime="00:00:56.00" entrycourse="SCM" />
                <RESULT eventid="1080" points="118" swimtime="00:03:44.69" resultid="1829" heatid="1970" lane="5" entrytime="00:03:35.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.07" />
                    <SPLIT distance="100" swimtime="00:01:49.88" />
                    <SPLIT distance="150" swimtime="00:02:50.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="113" swimtime="00:00:47.35" resultid="1830" heatid="2055" lane="1" entrytime="00:00:44.58" entrycourse="SCM" />
                <RESULT eventid="1204" points="127" swimtime="00:01:52.32" resultid="1831" heatid="2020" lane="2" entrytime="00:02:21.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luann" lastname="Miguel Mazur" birthdate="2007-01-10" gender="M" nation="BRA" license="365682" swrid="5596915" athleteid="1679" externalid="365682">
              <RESULTS>
                <RESULT eventid="1132" points="454" swimtime="00:09:36.70" resultid="1680" heatid="1994" lane="1" />
                <RESULT eventid="1100" points="472" swimtime="00:02:34.28" resultid="1681" heatid="1980" lane="4" entrytime="00:02:37.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                    <SPLIT distance="100" swimtime="00:01:14.69" />
                    <SPLIT distance="150" swimtime="00:01:54.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="460" swimtime="00:01:11.56" resultid="1682" heatid="2066" lane="5" entrytime="00:01:13.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="430" swimtime="00:02:11.61" resultid="1683" heatid="2035" lane="3" entrytime="00:02:08.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:04.86" />
                    <SPLIT distance="150" swimtime="00:01:38.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="488" swimtime="00:04:58.06" resultid="1684" heatid="2017" lane="5" entrytime="00:05:00.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:10.24" />
                    <SPLIT distance="150" swimtime="00:01:49.50" />
                    <SPLIT distance="200" swimtime="00:02:27.75" />
                    <SPLIT distance="250" swimtime="00:03:08.72" />
                    <SPLIT distance="300" swimtime="00:03:50.27" />
                    <SPLIT distance="350" swimtime="00:04:24.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Vitoria Gugel" birthdate="2011-12-08" gender="F" nation="BRA" license="365490" swrid="5588960" athleteid="1863" externalid="365490">
              <RESULTS>
                <RESULT eventid="1124" points="306" swimtime="00:11:48.42" resultid="1864" heatid="1991" lane="1" />
                <RESULT eventid="1092" points="305" swimtime="00:03:19.81" resultid="1865" heatid="1975" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.49" />
                    <SPLIT distance="100" swimtime="00:01:37.73" />
                    <SPLIT distance="150" swimtime="00:02:28.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="297" swimtime="00:01:15.25" resultid="1866" heatid="1959" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="250" swimtime="00:03:09.62" resultid="1867" heatid="2044" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.23" />
                    <SPLIT distance="100" swimtime="00:01:31.21" />
                    <SPLIT distance="150" swimtime="00:02:20.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="330" swimtime="00:06:14.51" resultid="1868" heatid="2011" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.91" />
                    <SPLIT distance="100" swimtime="00:01:31.72" />
                    <SPLIT distance="150" swimtime="00:02:20.12" />
                    <SPLIT distance="200" swimtime="00:03:06.54" />
                    <SPLIT distance="250" swimtime="00:03:57.57" />
                    <SPLIT distance="300" swimtime="00:04:49.48" />
                    <SPLIT distance="350" swimtime="00:05:32.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Luisa Lottermann" birthdate="2011-08-26" gender="F" nation="BRA" license="382238" swrid="5596909" athleteid="1779" externalid="382238">
              <RESULTS>
                <RESULT eventid="1124" points="298" swimtime="00:11:54.48" resultid="1780" heatid="1991" lane="6" />
                <RESULT eventid="1092" points="360" swimtime="00:03:09.13" resultid="1781" heatid="1976" lane="6" entrytime="00:03:35.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.56" />
                    <SPLIT distance="100" swimtime="00:01:32.04" />
                    <SPLIT distance="150" swimtime="00:02:20.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="293" swimtime="00:01:33.85" resultid="1782" heatid="2062" lane="6" entrytime="00:01:36.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="283" swimtime="00:02:47.92" resultid="1783" heatid="2027" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.78" />
                    <SPLIT distance="100" swimtime="00:01:22.53" />
                    <SPLIT distance="150" swimtime="00:02:06.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="288" swimtime="00:06:32.06" resultid="1784" heatid="2013" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.15" />
                    <SPLIT distance="100" swimtime="00:01:42.34" />
                    <SPLIT distance="150" swimtime="00:02:35.53" />
                    <SPLIT distance="200" swimtime="00:03:27.16" />
                    <SPLIT distance="250" swimtime="00:04:16.16" />
                    <SPLIT distance="300" swimtime="00:05:06.30" />
                    <SPLIT distance="350" swimtime="00:05:49.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia" lastname="Oliveira Faria" birthdate="2013-10-04" gender="F" nation="BRA" license="406697" swrid="5227019" athleteid="1890" externalid="406697">
              <RESULTS>
                <RESULT eventid="1162" points="68" swimtime="00:00:59.57" resultid="1891" heatid="2003" lane="5" />
                <RESULT eventid="1086" status="DSQ" swimtime="00:04:37.30" resultid="1892" heatid="1972" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.73" />
                    <SPLIT distance="100" swimtime="00:02:07.13" />
                    <SPLIT distance="150" swimtime="00:03:35.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="53" swimtime="00:01:15.20" resultid="1893" heatid="2058" lane="4" />
                <RESULT eventid="1210" points="97" swimtime="00:08:22.03" resultid="1894" heatid="2023" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Cordeiro Silva" birthdate="2011-09-04" gender="M" nation="BRA" license="380664" swrid="5596877" athleteid="1768" externalid="380664">
              <RESULTS>
                <RESULT eventid="1132" points="236" swimtime="00:11:56.74" resultid="1769" heatid="1994" lane="5" />
                <RESULT eventid="1100" points="232" swimtime="00:03:15.33" resultid="1770" heatid="1978" lane="4" entrytime="00:03:28.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.63" />
                    <SPLIT distance="100" swimtime="00:01:34.78" />
                    <SPLIT distance="150" swimtime="00:02:25.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="178" swimtime="00:01:19.69" resultid="1771" heatid="1965" lane="6" entrytime="00:01:15.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="233" swimtime="00:01:29.78" resultid="1772" heatid="2065" lane="6" entrytime="00:01:31.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="219" swimtime="00:06:29.17" resultid="1773" heatid="2015" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.83" />
                    <SPLIT distance="100" swimtime="00:01:33.88" />
                    <SPLIT distance="150" swimtime="00:02:26.30" />
                    <SPLIT distance="200" swimtime="00:03:16.84" />
                    <SPLIT distance="250" swimtime="00:04:10.22" />
                    <SPLIT distance="300" swimtime="00:05:01.83" />
                    <SPLIT distance="350" swimtime="00:05:46.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Zimmermann" birthdate="2010-01-19" gender="M" nation="BRA" license="357160" swrid="5588977" athleteid="1667" externalid="357160">
              <RESULTS>
                <RESULT eventid="1132" points="500" swimtime="00:09:18.40" resultid="1668" heatid="1996" lane="2" entrytime="00:09:14.38" entrycourse="SCM" />
                <RESULT eventid="1100" points="377" swimtime="00:02:46.33" resultid="1669" heatid="1980" lane="6" entrytime="00:02:49.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.95" />
                    <SPLIT distance="100" swimtime="00:01:20.54" />
                    <SPLIT distance="150" swimtime="00:02:03.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="425" swimtime="00:00:59.63" resultid="1670" heatid="1967" lane="6" entrytime="00:01:00.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="467" swimtime="00:02:08.00" resultid="1671" heatid="2035" lane="4" entrytime="00:02:08.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                    <SPLIT distance="100" swimtime="00:01:00.92" />
                    <SPLIT distance="150" swimtime="00:01:27.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="490" swimtime="00:04:57.74" resultid="1672" heatid="2017" lane="6" entrytime="00:05:12.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:10.90" />
                    <SPLIT distance="150" swimtime="00:01:48.17" />
                    <SPLIT distance="200" swimtime="00:02:25.07" />
                    <SPLIT distance="250" swimtime="00:03:07.22" />
                    <SPLIT distance="300" swimtime="00:03:49.56" />
                    <SPLIT distance="350" swimtime="00:04:24.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Emanuel Rech" birthdate="2013-12-02" gender="M" nation="BRA" license="380660" swrid="5588679" athleteid="1753" externalid="380660">
              <RESULTS>
                <RESULT eventid="1165" points="138" swimtime="00:00:41.99" resultid="1754" heatid="2004" lane="4" entrytime="00:00:41.11" entrycourse="SCM" />
                <RESULT eventid="1089" points="198" swimtime="00:03:07.88" resultid="1755" heatid="1974" lane="2" entrytime="00:03:10.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                    <SPLIT distance="100" swimtime="00:01:31.21" />
                    <SPLIT distance="150" swimtime="00:02:26.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1245" points="178" swimtime="00:01:25.79" resultid="1756" heatid="2043" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="192" swimtime="00:06:07.45" resultid="1757" heatid="2024" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Queiroz Da Costa" birthdate="2014-05-30" gender="F" nation="BRA" license="406698" swrid="5335148" athleteid="1895" externalid="406698">
              <RESULTS>
                <RESULT eventid="1156" points="77" swimtime="00:00:57.21" resultid="1896" heatid="2001" lane="6" entrytime="00:01:02.51" entrycourse="SCM" />
                <RESULT eventid="1080" points="132" swimtime="00:03:36.43" resultid="1897" heatid="1969" lane="2" />
                <RESULT eventid="1236" points="88" swimtime="00:00:56.59" resultid="1898" heatid="2039" lane="4" />
                <RESULT eventid="1204" points="103" swimtime="00:02:00.55" resultid="1899" heatid="2020" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Mariotti De Castro" birthdate="2008-06-27" gender="M" nation="BRA" license="329200" swrid="5596912" athleteid="1633" externalid="329200">
              <RESULTS>
                <RESULT eventid="1132" points="625" swimtime="00:08:38.59" resultid="1634" heatid="1996" lane="3" entrytime="00:08:31.20" entrycourse="SCM" />
                <RESULT eventid="1100" points="422" swimtime="00:02:40.13" resultid="1635" heatid="1980" lane="2" entrytime="00:02:43.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:01:18.66" />
                    <SPLIT distance="150" swimtime="00:01:58.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="533" swimtime="00:02:02.54" resultid="1636" heatid="2036" lane="3" entrytime="00:01:58.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                    <SPLIT distance="100" swimtime="00:01:01.25" />
                    <SPLIT distance="150" swimtime="00:01:32.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="554" swimtime="00:04:45.86" resultid="1637" heatid="2017" lane="3" entrytime="00:04:44.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                    <SPLIT distance="100" swimtime="00:01:05.51" />
                    <SPLIT distance="150" swimtime="00:01:42.70" />
                    <SPLIT distance="200" swimtime="00:02:19.14" />
                    <SPLIT distance="250" swimtime="00:03:00.94" />
                    <SPLIT distance="300" swimtime="00:03:42.67" />
                    <SPLIT distance="350" swimtime="00:04:15.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Bertelli Weirich" birthdate="2011-03-18" gender="F" nation="BRA" license="369534" swrid="5588552" athleteid="1714" externalid="369534">
              <RESULTS>
                <RESULT eventid="1124" points="376" swimtime="00:11:01.33" resultid="1715" heatid="1990" lane="4" />
                <RESULT eventid="1060" points="354" swimtime="00:01:10.99" resultid="1716" heatid="1962" lane="5" entrytime="00:01:07.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="287" swimtime="00:01:23.12" resultid="1717" heatid="2049" lane="1" entrytime="00:01:20.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="277" swimtime="00:03:03.30" resultid="1718" heatid="2044" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                    <SPLIT distance="100" swimtime="00:01:26.57" />
                    <SPLIT distance="150" swimtime="00:02:15.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="360" swimtime="00:06:03.70" resultid="1719" heatid="2011" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:01:26.87" />
                    <SPLIT distance="150" swimtime="00:02:14.35" />
                    <SPLIT distance="200" swimtime="00:03:00.02" />
                    <SPLIT distance="250" swimtime="00:03:50.48" />
                    <SPLIT distance="300" swimtime="00:04:42.12" />
                    <SPLIT distance="350" swimtime="00:05:23.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Do Prado Martins" birthdate="2008-10-17" gender="F" nation="BRA" license="369419" swrid="5596893" athleteid="1702" externalid="369419">
              <RESULTS>
                <RESULT eventid="1124" points="397" swimtime="00:10:49.56" resultid="1703" heatid="1990" lane="5" />
                <RESULT eventid="1092" points="407" swimtime="00:03:01.53" resultid="1704" heatid="1976" lane="4" entrytime="00:02:49.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.10" />
                    <SPLIT distance="100" swimtime="00:01:26.82" />
                    <SPLIT distance="150" swimtime="00:02:13.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="411" swimtime="00:01:23.81" resultid="1705" heatid="2062" lane="3" entrytime="00:01:19.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" status="DSQ" swimtime="00:02:49.66" resultid="1706" heatid="2044" lane="3" entrytime="00:02:46.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.13" />
                    <SPLIT distance="100" swimtime="00:01:17.50" />
                    <SPLIT distance="150" swimtime="00:02:02.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="410" swimtime="00:05:48.48" resultid="1707" heatid="2013" lane="3" entrytime="00:05:29.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                    <SPLIT distance="100" swimtime="00:01:17.81" />
                    <SPLIT distance="150" swimtime="00:02:03.22" />
                    <SPLIT distance="200" swimtime="00:02:48.18" />
                    <SPLIT distance="250" swimtime="00:03:36.00" />
                    <SPLIT distance="300" swimtime="00:04:24.56" />
                    <SPLIT distance="350" swimtime="00:05:07.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Luiza Bezerra Sedlacek" birthdate="2008-04-18" gender="F" nation="BRA" license="344607" swrid="4496478" athleteid="1649" externalid="344607">
              <RESULTS>
                <RESULT eventid="1168" points="367" swimtime="00:01:15.47" resultid="1650" heatid="2006" lane="4" entrytime="00:01:12.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="441" swimtime="00:10:26.86" resultid="1651" heatid="1992" lane="2" entrytime="00:10:25.58" entrycourse="SCM" />
                <RESULT eventid="1092" points="411" swimtime="00:03:00.98" resultid="1652" heatid="1975" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.80" />
                    <SPLIT distance="100" swimtime="00:01:25.88" />
                    <SPLIT distance="150" swimtime="00:02:12.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="523" swimtime="00:02:16.83" resultid="1653" heatid="2030" lane="4" entrytime="00:02:13.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:07.02" />
                    <SPLIT distance="150" swimtime="00:01:42.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="465" swimtime="00:05:34.09" resultid="1654" heatid="2013" lane="4" entrytime="00:05:36.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                    <SPLIT distance="100" swimtime="00:01:17.69" />
                    <SPLIT distance="150" swimtime="00:02:00.65" />
                    <SPLIT distance="200" swimtime="00:02:42.59" />
                    <SPLIT distance="250" swimtime="00:03:30.18" />
                    <SPLIT distance="300" swimtime="00:04:18.38" />
                    <SPLIT distance="350" swimtime="00:04:56.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Henrique Marca Dos Santos" birthdate="2015-03-28" gender="M" nation="BRA" license="406695" swrid="4991165" athleteid="1880" externalid="406695">
              <RESULTS>
                <RESULT eventid="1159" points="42" swimtime="00:01:02.22" resultid="1881" heatid="2002" lane="2" />
                <RESULT eventid="1115" points="50" swimtime="00:01:07.42" resultid="1882" heatid="1986" lane="6" entrytime="00:01:07.12" entrycourse="SCM" />
                <RESULT eventid="1239" points="49" swimtime="00:01:00.20" resultid="1883" heatid="2041" lane="2" entrytime="00:01:00.14" entrycourse="SCM" />
                <RESULT eventid="1207" points="57" swimtime="00:02:07.33" resultid="1884" heatid="2022" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Assakura" birthdate="2010-06-29" gender="F" nation="BRA" license="376473" swrid="5596868" athleteid="1785" externalid="376473">
              <RESULTS>
                <RESULT eventid="1140" points="345" swimtime="00:02:49.50" resultid="1786" heatid="1998" lane="5" entrytime="00:02:55.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.01" />
                    <SPLIT distance="100" swimtime="00:01:23.70" />
                    <SPLIT distance="150" swimtime="00:02:07.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="404" swimtime="00:10:45.75" resultid="1787" heatid="1991" lane="2" />
                <RESULT eventid="1092" points="435" swimtime="00:02:57.52" resultid="1788" heatid="1976" lane="1" entrytime="00:03:20.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                    <SPLIT distance="100" swimtime="00:01:25.37" />
                    <SPLIT distance="150" swimtime="00:02:11.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="390" swimtime="00:02:30.90" resultid="1789" heatid="2030" lane="1" entrytime="00:02:30.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:01:12.70" />
                    <SPLIT distance="150" swimtime="00:01:52.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="395" swimtime="00:05:52.69" resultid="1790" heatid="2012" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.67" />
                    <SPLIT distance="100" swimtime="00:01:28.15" />
                    <SPLIT distance="150" swimtime="00:02:12.80" />
                    <SPLIT distance="200" swimtime="00:02:56.56" />
                    <SPLIT distance="250" swimtime="00:03:43.52" />
                    <SPLIT distance="300" swimtime="00:04:30.94" />
                    <SPLIT distance="350" swimtime="00:05:13.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Pedro Signor" birthdate="2005-12-20" gender="M" nation="BRA" license="375814" swrid="5596925" athleteid="1738" externalid="375814">
              <RESULTS>
                <RESULT eventid="1176" points="427" swimtime="00:01:03.44" resultid="1739" heatid="2010" lane="1" entrytime="00:01:03.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="284" swimtime="00:11:14.27" resultid="1740" heatid="1994" lane="4" />
                <RESULT eventid="1068" points="378" swimtime="00:01:01.99" resultid="1741" heatid="1967" lane="2" entrytime="00:00:59.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="366" swimtime="00:01:07.56" resultid="1742" heatid="2052" lane="3" entrytime="00:01:06.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="357" swimtime="00:05:30.70" resultid="1743" heatid="2016" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                    <SPLIT distance="100" swimtime="00:01:17.39" />
                    <SPLIT distance="150" swimtime="00:01:59.98" />
                    <SPLIT distance="200" swimtime="00:02:43.48" />
                    <SPLIT distance="250" swimtime="00:03:29.20" />
                    <SPLIT distance="300" swimtime="00:04:16.20" />
                    <SPLIT distance="350" swimtime="00:04:55.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Claudio" lastname="Rohnelt" birthdate="2010-03-08" gender="M" nation="BRA" license="357954" swrid="5596935" athleteid="1673" externalid="357954">
              <RESULTS>
                <RESULT eventid="1176" points="178" swimtime="00:01:24.85" resultid="1674" heatid="2008" lane="3" entrytime="00:01:17.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="311" swimtime="00:10:53.84" resultid="1675" heatid="1994" lane="6" />
                <RESULT eventid="1068" points="273" swimtime="00:01:09.05" resultid="1676" heatid="1963" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="201" swimtime="00:03:02.40" resultid="1677" heatid="2045" lane="3" entrytime="00:02:52.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:25.52" />
                    <SPLIT distance="150" swimtime="00:02:13.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="262" swimtime="00:06:06.68" resultid="1678" heatid="2014" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.24" />
                    <SPLIT distance="100" swimtime="00:01:27.35" />
                    <SPLIT distance="150" swimtime="00:02:16.49" />
                    <SPLIT distance="200" swimtime="00:03:03.13" />
                    <SPLIT distance="250" swimtime="00:03:55.53" />
                    <SPLIT distance="300" swimtime="00:04:48.54" />
                    <SPLIT distance="350" swimtime="00:05:28.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Vargas Moreira" birthdate="2014-03-09" gender="F" nation="BRA" license="392014" swrid="4904290" athleteid="1853" externalid="392014">
              <RESULTS>
                <RESULT eventid="1156" points="108" swimtime="00:00:51.09" resultid="1854" heatid="2001" lane="5" entrytime="00:00:52.72" entrycourse="SCM" />
                <RESULT eventid="1080" points="223" swimtime="00:03:01.82" resultid="1855" heatid="1970" lane="3" entrytime="00:03:13.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.89" />
                    <SPLIT distance="100" swimtime="00:01:29.32" />
                    <SPLIT distance="150" swimtime="00:02:17.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="117" swimtime="00:00:51.53" resultid="1856" heatid="2040" lane="4" entrytime="00:00:55.15" entrycourse="SCM" />
                <RESULT eventid="1204" points="160" swimtime="00:01:44.05" resultid="1857" heatid="2019" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Colaco Da Conceicao" birthdate="2011-05-25" gender="F" nation="BRA" license="369535" swrid="5588601" athleteid="1720" externalid="369535">
              <RESULTS>
                <RESULT eventid="1168" points="223" swimtime="00:01:29.10" resultid="1721" heatid="2006" lane="1" entrytime="00:01:32.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="265" swimtime="00:03:05.05" resultid="1722" heatid="1997" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.52" />
                    <SPLIT distance="100" swimtime="00:01:30.55" />
                    <SPLIT distance="150" swimtime="00:02:17.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="381" swimtime="00:10:58.38" resultid="1723" heatid="1991" lane="4" />
                <RESULT eventid="1216" points="372" swimtime="00:02:33.35" resultid="1724" heatid="2028" lane="4" entrytime="00:02:35.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                    <SPLIT distance="100" swimtime="00:01:14.58" />
                    <SPLIT distance="150" swimtime="00:01:54.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="314" swimtime="00:06:20.80" resultid="1725" heatid="2012" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.55" />
                    <SPLIT distance="100" swimtime="00:01:32.01" />
                    <SPLIT distance="150" swimtime="00:02:21.09" />
                    <SPLIT distance="200" swimtime="00:03:09.11" />
                    <SPLIT distance="250" swimtime="00:04:00.85" />
                    <SPLIT distance="300" swimtime="00:04:54.30" />
                    <SPLIT distance="350" swimtime="00:05:37.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Paiz Ribeiro" birthdate="2006-02-17" gender="M" nation="BRA" license="297583" swrid="5596921" athleteid="1619" externalid="297583">
              <RESULTS>
                <RESULT eventid="1148" points="359" swimtime="00:02:28.58" resultid="1620" heatid="1999" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:14.77" />
                    <SPLIT distance="150" swimtime="00:01:51.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="506" swimtime="00:09:16.40" resultid="1621" heatid="1993" lane="3" />
                <RESULT eventid="1256" points="481" swimtime="00:02:16.31" resultid="1622" heatid="2046" lane="4" entrytime="00:02:13.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                    <SPLIT distance="100" swimtime="00:01:04.15" />
                    <SPLIT distance="150" swimtime="00:01:39.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="456" swimtime="00:05:05.05" resultid="1623" heatid="2017" lane="4" entrytime="00:04:52.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                    <SPLIT distance="100" swimtime="00:01:06.33" />
                    <SPLIT distance="150" swimtime="00:01:48.01" />
                    <SPLIT distance="200" swimtime="00:02:28.27" />
                    <SPLIT distance="250" swimtime="00:03:11.65" />
                    <SPLIT distance="300" swimtime="00:03:55.91" />
                    <SPLIT distance="350" swimtime="00:04:30.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Domingues" birthdate="2013-10-22" gender="M" nation="BRA" license="380661" swrid="5676301" athleteid="1758" externalid="380661">
              <RESULTS>
                <RESULT eventid="1165" points="99" swimtime="00:00:46.94" resultid="1759" heatid="2004" lane="5" entrytime="00:00:45.02" entrycourse="SCM" />
                <RESULT eventid="1089" status="DSQ" swimtime="00:03:22.55" resultid="1760" heatid="1973" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.26" />
                    <SPLIT distance="100" swimtime="00:01:35.21" />
                    <SPLIT distance="150" swimtime="00:02:39.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" status="DNS" swimtime="00:00:00.00" resultid="1761" heatid="2059" lane="4" entrytime="00:00:54.44" entrycourse="SCM" />
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="1762" heatid="2024" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Breno" lastname="Zanella Janke" birthdate="2011-04-26" gender="M" nation="BRA" license="365697" swrid="5588970" athleteid="1708" externalid="365697">
              <RESULTS>
                <RESULT eventid="1176" points="293" swimtime="00:01:11.86" resultid="1709" heatid="2009" lane="6" entrytime="00:01:16.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="386" swimtime="00:10:08.90" resultid="1710" heatid="1994" lane="2" />
                <RESULT eventid="1100" points="309" swimtime="00:02:57.70" resultid="1711" heatid="1979" lane="2" entrytime="00:03:10.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                    <SPLIT distance="100" swimtime="00:01:25.42" />
                    <SPLIT distance="150" swimtime="00:02:11.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="299" swimtime="00:01:22.66" resultid="1712" heatid="2065" lane="4" entrytime="00:01:24.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="362" swimtime="00:05:29.20" resultid="1713" heatid="2015" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.20" />
                    <SPLIT distance="100" swimtime="00:01:20.08" />
                    <SPLIT distance="150" swimtime="00:02:02.62" />
                    <SPLIT distance="200" swimtime="00:02:43.80" />
                    <SPLIT distance="250" swimtime="00:03:28.98" />
                    <SPLIT distance="300" swimtime="00:04:14.58" />
                    <SPLIT distance="350" swimtime="00:04:52.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Pedro Serafini" birthdate="2012-05-15" gender="M" nation="BRA" license="365488" swrid="5596924" athleteid="1803" externalid="365488">
              <RESULTS>
                <RESULT eventid="1121" points="165" swimtime="00:01:21.73" resultid="1804" heatid="1989" lane="5" entrytime="00:01:23.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1089" points="164" swimtime="00:03:19.98" resultid="1805" heatid="1974" lane="6" entrytime="00:03:24.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.11" />
                    <SPLIT distance="100" swimtime="00:01:36.66" />
                    <SPLIT distance="150" swimtime="00:02:37.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="118" swimtime="00:00:50.73" resultid="1806" heatid="2060" lane="5" entrytime="00:00:52.24" entrycourse="SCM" />
                <RESULT eventid="1213" points="191" swimtime="00:06:08.07" resultid="1807" heatid="2025" lane="4" entrytime="00:06:17.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jordana" lastname="Rinaldini" birthdate="2004-09-13" gender="F" nation="BRA" license="342426" swrid="5596933" athleteid="1638" externalid="342426">
              <RESULTS>
                <RESULT eventid="1140" points="313" swimtime="00:02:55.01" resultid="1639" heatid="1998" lane="2" entrytime="00:02:47.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                    <SPLIT distance="100" swimtime="00:01:23.64" />
                    <SPLIT distance="150" swimtime="00:02:10.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="371" swimtime="00:03:07.12" resultid="1640" heatid="1976" lane="2" entrytime="00:03:01.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                    <SPLIT distance="100" swimtime="00:01:27.10" />
                    <SPLIT distance="150" swimtime="00:02:16.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="345" swimtime="00:01:28.88" resultid="1641" heatid="2062" lane="4" entrytime="00:01:24.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="333" swimtime="00:02:39.09" resultid="1642" heatid="2029" lane="1" entrytime="00:02:33.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                    <SPLIT distance="100" swimtime="00:01:15.25" />
                    <SPLIT distance="150" swimtime="00:01:57.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ramirez Vasconcelos" birthdate="2011-04-06" gender="M" nation="BRA" license="392013" swrid="4863662" athleteid="1847" externalid="392013">
              <RESULTS>
                <RESULT eventid="1132" points="296" swimtime="00:11:05.20" resultid="1848" heatid="1993" lane="2" />
                <RESULT eventid="1100" points="222" swimtime="00:03:18.29" resultid="1849" heatid="1977" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.69" />
                    <SPLIT distance="100" swimtime="00:01:34.22" />
                    <SPLIT distance="150" swimtime="00:02:26.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="275" swimtime="00:01:08.94" resultid="1850" heatid="1965" lane="5" entrytime="00:01:14.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="225" swimtime="00:01:30.85" resultid="1851" heatid="2065" lane="1" entrytime="00:01:29.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="260" swimtime="00:06:07.52" resultid="1852" heatid="2014" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                    <SPLIT distance="100" swimtime="00:01:30.03" />
                    <SPLIT distance="150" swimtime="00:02:17.28" />
                    <SPLIT distance="200" swimtime="00:03:03.26" />
                    <SPLIT distance="250" swimtime="00:03:56.00" />
                    <SPLIT distance="300" swimtime="00:04:49.10" />
                    <SPLIT distance="350" swimtime="00:05:29.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Luis Lottermann" birthdate="2014-10-08" gender="M" nation="BRA" license="382237" swrid="5596908" athleteid="1774" externalid="382237">
              <RESULTS>
                <RESULT eventid="1159" points="111" swimtime="00:00:45.15" resultid="1775" heatid="2002" lane="3" entrytime="00:00:45.02" entrycourse="SCM" />
                <RESULT eventid="1083" points="184" swimtime="00:02:54.46" resultid="1776" heatid="1971" lane="3" entrytime="00:03:03.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.03" />
                    <SPLIT distance="100" swimtime="00:01:25.43" />
                    <SPLIT distance="150" swimtime="00:02:11.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" points="159" swimtime="00:00:37.14" resultid="1777" heatid="2057" lane="3" entrytime="00:00:37.71" entrycourse="SCM" />
                <RESULT eventid="1207" points="149" swimtime="00:01:32.88" resultid="1778" heatid="2022" lane="3" entrytime="00:01:37.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emanuel" lastname="Ranieri" birthdate="2011-01-24" gender="M" nation="BRA" license="390838" swrid="5596930" athleteid="1816" externalid="390838">
              <RESULTS>
                <RESULT eventid="1148" points="263" swimtime="00:02:44.74" resultid="1817" heatid="1999" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:01:21.05" />
                    <SPLIT distance="150" swimtime="00:02:03.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="331" swimtime="00:10:40.77" resultid="1818" heatid="1993" lane="4" />
                <RESULT eventid="1100" points="284" swimtime="00:03:02.65" resultid="1819" heatid="1977" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.22" />
                    <SPLIT distance="100" swimtime="00:01:26.98" />
                    <SPLIT distance="150" swimtime="00:02:14.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="313" swimtime="00:02:26.32" resultid="1820" heatid="2033" lane="2" entrytime="00:02:27.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                    <SPLIT distance="100" swimtime="00:01:12.04" />
                    <SPLIT distance="150" swimtime="00:01:50.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="296" swimtime="00:05:52.20" resultid="1821" heatid="2016" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                    <SPLIT distance="100" swimtime="00:01:27.84" />
                    <SPLIT distance="150" swimtime="00:02:13.29" />
                    <SPLIT distance="200" swimtime="00:02:56.69" />
                    <SPLIT distance="250" swimtime="00:03:44.85" />
                    <SPLIT distance="300" swimtime="00:04:34.33" />
                    <SPLIT distance="350" swimtime="00:05:14.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Tolentino Smarczewski" birthdate="2008-09-01" gender="M" nation="BRA" license="378818" swrid="5596941" athleteid="1744" externalid="378818">
              <RESULTS>
                <RESULT eventid="1132" points="482" swimtime="00:09:25.32" resultid="1745" heatid="1995" lane="6" />
                <RESULT eventid="1100" points="380" swimtime="00:02:45.86" resultid="1746" heatid="1979" lane="3" entrytime="00:02:59.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="100" swimtime="00:01:18.66" />
                    <SPLIT distance="150" swimtime="00:02:01.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="345" swimtime="00:01:18.76" resultid="1747" heatid="2066" lane="6" entrytime="00:01:22.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="453" swimtime="00:02:09.34" resultid="1748" heatid="2036" lane="6" entrytime="00:02:07.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.98" />
                    <SPLIT distance="100" swimtime="00:01:02.63" />
                    <SPLIT distance="150" swimtime="00:01:36.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="358" swimtime="00:05:30.40" resultid="1749" heatid="2016" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                    <SPLIT distance="100" swimtime="00:01:24.99" />
                    <SPLIT distance="150" swimtime="00:02:09.16" />
                    <SPLIT distance="200" swimtime="00:02:52.89" />
                    <SPLIT distance="250" swimtime="00:03:36.98" />
                    <SPLIT distance="300" swimtime="00:04:21.41" />
                    <SPLIT distance="350" swimtime="00:04:56.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Balduíno" birthdate="2009-06-24" gender="M" nation="BRA" license="370764" swrid="5596870" athleteid="1732" externalid="370764">
              <RESULTS>
                <RESULT eventid="1176" points="393" swimtime="00:01:05.20" resultid="1733" heatid="2010" lane="6" entrytime="00:01:04.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="451" swimtime="00:09:37.91" resultid="1734" heatid="1996" lane="5" entrytime="00:09:33.89" entrycourse="SCM" />
                <RESULT eventid="1256" points="380" swimtime="00:02:27.39" resultid="1735" heatid="2046" lane="5" entrytime="00:02:28.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                    <SPLIT distance="150" swimtime="00:01:49.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="428" swimtime="00:02:11.80" resultid="1736" heatid="2034" lane="3" entrytime="00:02:17.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="100" swimtime="00:01:04.12" />
                    <SPLIT distance="150" swimtime="00:01:38.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="430" swimtime="00:05:11.09" resultid="1737" heatid="2016" lane="3" entrytime="00:05:12.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                    <SPLIT distance="100" swimtime="00:01:08.64" />
                    <SPLIT distance="150" swimtime="00:01:49.30" />
                    <SPLIT distance="200" swimtime="00:02:29.22" />
                    <SPLIT distance="250" swimtime="00:03:13.83" />
                    <SPLIT distance="300" swimtime="00:03:59.43" />
                    <SPLIT distance="350" swimtime="00:04:36.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Kupicki" birthdate="2004-03-02" gender="F" nation="BRA" license="311897" swrid="5624094" athleteid="1624" externalid="311897">
              <RESULTS>
                <RESULT eventid="1060" points="355" swimtime="00:01:10.96" resultid="1625" heatid="1962" lane="4" entrytime="00:01:06.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" status="DNS" swimtime="00:00:00.00" resultid="1626" heatid="2062" lane="5" entrytime="00:01:28.08" entrycourse="SCM" />
                <RESULT eventid="1216" points="332" swimtime="00:02:39.25" resultid="1627" heatid="2030" lane="5" entrytime="00:02:27.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.20" />
                    <SPLIT distance="100" swimtime="00:01:13.94" />
                    <SPLIT distance="150" swimtime="00:01:55.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Gaio" birthdate="2012-11-13" gender="F" nation="BRA" license="390842" swrid="5596901" athleteid="1832" externalid="390842">
              <RESULTS>
                <RESULT eventid="1162" points="59" swimtime="00:01:02.36" resultid="1833" heatid="2003" lane="2" entrytime="00:01:04.60" entrycourse="SCM" />
                <RESULT eventid="1118" points="90" swimtime="00:01:51.75" resultid="1834" heatid="1987" lane="2" entrytime="00:02:17.33" entrycourse="SCM" />
                <RESULT eventid="1242" status="DSQ" swimtime="00:02:09.13" resultid="1835" heatid="2042" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Gamero Prado" birthdate="2007-05-16" gender="F" nation="BRA" license="305973" swrid="5596903" athleteid="1628" externalid="305973">
              <RESULTS>
                <RESULT eventid="1124" points="467" swimtime="00:10:15.21" resultid="1629" heatid="1992" lane="3" entrytime="00:10:12.66" entrycourse="SCM" />
                <RESULT eventid="1060" points="435" swimtime="00:01:06.30" resultid="1630" heatid="1961" lane="4" entrytime="00:01:10.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="455" swimtime="00:02:23.37" resultid="1631" heatid="2026" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:09.85" />
                    <SPLIT distance="150" swimtime="00:01:47.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="366" swimtime="00:06:01.78" resultid="1632" heatid="2013" lane="1" entrytime="00:06:06.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                    <SPLIT distance="100" swimtime="00:01:19.54" />
                    <SPLIT distance="150" swimtime="00:02:07.52" />
                    <SPLIT distance="200" swimtime="00:02:54.84" />
                    <SPLIT distance="250" swimtime="00:03:48.57" />
                    <SPLIT distance="300" swimtime="00:04:42.18" />
                    <SPLIT distance="350" swimtime="00:05:22.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laisa" lastname="Bernardini" birthdate="2012-06-25" gender="F" nation="BRA" license="390843" swrid="5596872" athleteid="1836" externalid="390843">
              <RESULTS>
                <RESULT eventid="1162" points="136" swimtime="00:00:47.34" resultid="1837" heatid="2003" lane="4" entrytime="00:00:47.77" entrycourse="SCM" />
                <RESULT eventid="1086" points="200" swimtime="00:03:28.34" resultid="1838" heatid="1972" lane="3" entrytime="00:03:28.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.07" />
                    <SPLIT distance="100" swimtime="00:01:42.54" />
                    <SPLIT distance="150" swimtime="00:02:41.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="178" swimtime="00:01:37.52" resultid="1839" heatid="2042" lane="3" entrytime="00:01:38.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1210" points="200" swimtime="00:06:35.39" resultid="1840" heatid="2023" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Alves Serafini" birthdate="2008-04-15" gender="M" nation="BRA" license="351644" swrid="5596867" athleteid="1797" externalid="351644">
              <RESULTS>
                <RESULT eventid="1132" points="485" swimtime="00:09:24.11" resultid="1798" heatid="1994" lane="3" />
                <RESULT eventid="1068" points="422" swimtime="00:00:59.74" resultid="1799" heatid="1968" lane="1" entrytime="00:00:57.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="307" swimtime="00:01:21.86" resultid="1800" heatid="2066" lane="1" entrytime="00:01:21.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="453" swimtime="00:02:09.32" resultid="1801" heatid="2036" lane="1" entrytime="00:02:07.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                    <SPLIT distance="100" swimtime="00:01:02.67" />
                    <SPLIT distance="150" swimtime="00:01:36.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="402" swimtime="00:05:18.01" resultid="1802" heatid="2016" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:07.29" />
                    <SPLIT distance="150" swimtime="00:01:49.31" />
                    <SPLIT distance="200" swimtime="00:02:30.28" />
                    <SPLIT distance="250" swimtime="00:03:17.05" />
                    <SPLIT distance="300" swimtime="00:04:05.04" />
                    <SPLIT distance="350" swimtime="00:04:41.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Dillenburg Benetti" birthdate="2011-03-10" gender="M" nation="BRA" license="368119" swrid="5588656" athleteid="1691" externalid="368119">
              <RESULTS>
                <RESULT eventid="1132" points="384" swimtime="00:10:09.76" resultid="1692" heatid="1995" lane="5" />
                <RESULT eventid="1100" points="294" swimtime="00:03:00.68" resultid="1693" heatid="1979" lane="6" entrytime="00:03:19.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                    <SPLIT distance="100" swimtime="00:01:25.69" />
                    <SPLIT distance="150" swimtime="00:02:13.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="286" swimtime="00:01:13.29" resultid="1694" heatid="2051" lane="3" entrytime="00:01:13.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="336" swimtime="00:02:22.81" resultid="1695" heatid="2034" lane="5" entrytime="00:02:22.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="100" swimtime="00:01:09.05" />
                    <SPLIT distance="150" swimtime="00:01:46.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="328" swimtime="00:05:40.22" resultid="1696" heatid="2014" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                    <SPLIT distance="100" swimtime="00:01:24.17" />
                    <SPLIT distance="150" swimtime="00:02:07.73" />
                    <SPLIT distance="200" swimtime="00:02:49.18" />
                    <SPLIT distance="250" swimtime="00:03:37.26" />
                    <SPLIT distance="300" swimtime="00:04:25.92" />
                    <SPLIT distance="350" swimtime="00:05:03.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Gabriel Dalchau" birthdate="2014-08-27" gender="M" nation="BRA" license="402118" swrid="5661346" athleteid="1875" externalid="402118">
              <RESULTS>
                <RESULT eventid="1115" points="73" swimtime="00:00:59.63" resultid="1876" heatid="1986" lane="1" entrytime="00:01:02.11" entrycourse="SCM" />
                <RESULT eventid="1083" points="114" swimtime="00:03:24.54" resultid="1877" heatid="1971" lane="2" entrytime="00:03:29.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.77" />
                    <SPLIT distance="100" swimtime="00:01:38.53" />
                    <SPLIT distance="150" swimtime="00:02:33.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1239" points="91" swimtime="00:00:49.13" resultid="1878" heatid="2041" lane="3" entrytime="00:00:50.59" entrycourse="SCM" />
                <RESULT eventid="1207" points="78" swimtime="00:01:55.27" resultid="1879" heatid="2022" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marianna" lastname="Galvao Oliveira" birthdate="2014-03-18" gender="F" nation="BRA" license="390835" swrid="5596902" athleteid="1813" externalid="390835">
              <RESULTS>
                <RESULT eventid="1112" points="167" swimtime="00:00:51.49" resultid="1814" heatid="1984" lane="3" entrytime="00:00:49.35" entrycourse="SCM" />
                <RESULT eventid="1080" points="159" swimtime="00:03:23.34" resultid="1815" heatid="1970" lane="1" entrytime="00:03:38.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.40" />
                    <SPLIT distance="100" swimtime="00:01:36.55" />
                    <SPLIT distance="150" swimtime="00:02:31.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Flavia" lastname="De Metz" birthdate="2011-01-07" gender="F" nation="BRA" license="390846" swrid="5596887" athleteid="1841" externalid="390846">
              <RESULTS>
                <RESULT eventid="1140" points="321" swimtime="00:02:53.63" resultid="1842" heatid="1998" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.15" />
                    <SPLIT distance="100" swimtime="00:01:25.69" />
                    <SPLIT distance="150" swimtime="00:02:10.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="337" swimtime="00:11:25.44" resultid="1843" heatid="1990" lane="2" />
                <RESULT eventid="1060" points="374" swimtime="00:01:09.73" resultid="1844" heatid="1961" lane="3" entrytime="00:01:10.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="387" swimtime="00:02:31.35" resultid="1845" heatid="2029" lane="5" entrytime="00:02:32.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="100" swimtime="00:01:13.31" />
                    <SPLIT distance="150" swimtime="00:01:52.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="312" swimtime="00:06:21.38" resultid="1846" heatid="2011" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.94" />
                    <SPLIT distance="100" swimtime="00:01:37.17" />
                    <SPLIT distance="150" swimtime="00:02:24.55" />
                    <SPLIT distance="200" swimtime="00:03:11.56" />
                    <SPLIT distance="250" swimtime="00:04:04.69" />
                    <SPLIT distance="300" swimtime="00:04:59.15" />
                    <SPLIT distance="350" swimtime="00:05:40.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Danilo" lastname="Rodrigues" birthdate="2011-05-23" gender="M" nation="BRA" license="370763" swrid="5596934" athleteid="1726" externalid="370763">
              <RESULTS>
                <RESULT eventid="1132" points="330" swimtime="00:10:41.56" resultid="1727" heatid="1993" lane="5" />
                <RESULT eventid="1100" points="285" swimtime="00:03:02.48" resultid="1728" heatid="1978" lane="3" entrytime="00:03:25.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                    <SPLIT distance="100" swimtime="00:01:28.64" />
                    <SPLIT distance="150" swimtime="00:02:15.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="251" swimtime="00:02:49.34" resultid="1729" heatid="2045" lane="2" entrytime="00:03:05.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:21.16" />
                    <SPLIT distance="150" swimtime="00:02:06.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="310" swimtime="00:02:26.79" resultid="1730" heatid="2033" lane="4" entrytime="00:02:27.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                    <SPLIT distance="100" swimtime="00:01:11.99" />
                    <SPLIT distance="150" swimtime="00:01:50.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="319" swimtime="00:05:43.33" resultid="1731" heatid="2015" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:21.18" />
                    <SPLIT distance="150" swimtime="00:02:07.76" />
                    <SPLIT distance="200" swimtime="00:02:50.96" />
                    <SPLIT distance="250" swimtime="00:03:39.67" />
                    <SPLIT distance="300" swimtime="00:04:27.42" />
                    <SPLIT distance="350" swimtime="00:05:06.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Sehn Uren" birthdate="2009-10-15" gender="F" nation="BRA" license="357159" swrid="5596937" athleteid="1661" externalid="357159">
              <RESULTS>
                <RESULT eventid="1168" points="290" swimtime="00:01:21.63" resultid="1662" heatid="2005" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="313" swimtime="00:11:42.97" resultid="1663" heatid="1990" lane="3" />
                <RESULT eventid="1292" points="370" swimtime="00:01:26.81" resultid="1664" heatid="2062" lane="1" entrytime="00:01:29.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="374" swimtime="00:02:33.02" resultid="1665" heatid="2028" lane="1" entrytime="00:02:41.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                    <SPLIT distance="100" swimtime="00:01:15.57" />
                    <SPLIT distance="150" swimtime="00:01:55.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="377" swimtime="00:05:58.30" resultid="1666" heatid="2012" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.50" />
                    <SPLIT distance="100" swimtime="00:01:26.99" />
                    <SPLIT distance="150" swimtime="00:02:14.82" />
                    <SPLIT distance="200" swimtime="00:03:00.23" />
                    <SPLIT distance="250" swimtime="00:03:48.58" />
                    <SPLIT distance="300" swimtime="00:04:36.81" />
                    <SPLIT distance="350" swimtime="00:05:19.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Henrique Wiebbeling" birthdate="2003-08-06" gender="M" nation="BRA" license="290420" swrid="4471225" athleteid="1614" externalid="290420">
              <RESULTS>
                <RESULT eventid="1132" status="DNS" swimtime="00:00:00.00" resultid="1615" heatid="1996" lane="4" entrytime="00:09:08.94" entrycourse="SCM" />
                <RESULT eventid="1068" status="DNS" swimtime="00:00:00.00" resultid="1616" heatid="1963" lane="2" />
                <RESULT eventid="1272" points="340" swimtime="00:01:09.24" resultid="1617" heatid="2052" lane="5" entrytime="00:01:07.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="465" swimtime="00:02:08.24" resultid="1618" heatid="2036" lane="4" entrytime="00:02:03.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="100" swimtime="00:01:01.33" />
                    <SPLIT distance="150" swimtime="00:01:34.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13068" nation="BRA" region="PR" clubid="1900" swrid="93787" name="Sociedade Morgenau" shortname="Morgenau">
          <ATHLETES>
            <ATHLETE firstname="Heloisa" lastname="Nitz Costa" birthdate="2015-02-09" gender="F" nation="BRA" license="397328" swrid="5641773" athleteid="1901" externalid="397328">
              <RESULTS>
                <RESULT eventid="1280" points="111" swimtime="00:00:47.60" resultid="1902" heatid="2055" lane="2" entrytime="00:00:43.46" entrycourse="SCM" />
                <RESULT eventid="1204" points="141" swimtime="00:01:48.44" resultid="1903" heatid="2019" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13025" nation="BRA" region="PR" clubid="1419" swrid="93779" name="Instituto Desportos Aquáticos De Foz Do Iguaçu" shortname="Cataratas Natação">
          <ATHLETES>
            <ATHLETE firstname="Lucas" lastname="Marques Petry" birthdate="2008-01-08" gender="M" nation="BRA" license="392351" swrid="4711489" athleteid="1485" externalid="392351" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1176" points="220" swimtime="00:01:19.10" resultid="1486" heatid="2007" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="377" swimtime="00:10:13.41" resultid="1487" heatid="1995" lane="3" entrytime="00:11:20.41" entrycourse="SCM" />
                <RESULT eventid="1068" points="323" swimtime="00:01:05.33" resultid="1488" heatid="1966" lane="6" entrytime="00:01:05.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="184" swimtime="00:01:24.87" resultid="1489" heatid="2051" lane="4" entrytime="00:01:22.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="342" swimtime="00:02:22.05" resultid="1490" heatid="2033" lane="3" entrytime="00:02:25.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                    <SPLIT distance="100" swimtime="00:01:08.41" />
                    <SPLIT distance="150" swimtime="00:01:45.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Mattiello" birthdate="2009-04-11" gender="F" nation="BRA" license="367011" swrid="5596914" athleteid="1474" externalid="367011" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1124" points="371" swimtime="00:11:04.04" resultid="1475" heatid="1992" lane="1" entrytime="00:11:02.88" entrycourse="SCM" />
                <RESULT eventid="1060" points="378" swimtime="00:01:09.47" resultid="1476" heatid="1962" lane="1" entrytime="00:01:08.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="292" swimtime="00:01:22.69" resultid="1477" heatid="2049" lane="6" entrytime="00:01:21.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" status="DSQ" swimtime="00:02:28.97" resultid="1478" heatid="2029" lane="3" entrytime="00:02:31.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="100" swimtime="00:01:14.62" />
                    <SPLIT distance="150" swimtime="00:01:52.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Abraao" lastname="Felipe Oliveira" birthdate="2012-05-20" gender="M" nation="BRA" license="400457" swrid="5420917" athleteid="1561" externalid="400457" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1121" points="139" swimtime="00:01:26.36" resultid="1562" heatid="1989" lane="1" entrytime="00:01:26.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1089" status="DSQ" swimtime="00:03:45.97" resultid="1563" heatid="1973" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.20" />
                    <SPLIT distance="100" swimtime="00:01:48.59" />
                    <SPLIT distance="150" swimtime="00:02:56.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="125" swimtime="00:00:49.90" resultid="1564" heatid="2059" lane="3" entrytime="00:00:53.89" entrycourse="SCM" />
                <RESULT eventid="1245" points="75" swimtime="00:01:54.32" resultid="1565" heatid="2043" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benjamin" lastname="Perius Goncalves De Lima" birthdate="2016-06-09" gender="M" nation="BRA" license="407798" athleteid="1592" externalid="407798">
              <RESULTS>
                <RESULT eventid="1110" points="88" swimtime="00:00:49.54" resultid="1593" heatid="1982" lane="4" />
                <RESULT eventid="1234" points="95" swimtime="00:00:44.09" resultid="1594" heatid="2038" lane="3" />
                <RESULT eventid="1202" points="52" swimtime="00:01:06.62" resultid="1595" heatid="2018" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Ferrari Ghellere" birthdate="2014-07-01" gender="F" nation="BRA" license="372038" swrid="5596895" athleteid="1520" externalid="372038" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1156" points="119" swimtime="00:00:49.46" resultid="1521" heatid="2001" lane="2" entrytime="00:00:50.09" entrycourse="SCM" />
                <RESULT eventid="1080" points="218" swimtime="00:03:03.09" resultid="1522" heatid="1970" lane="4" entrytime="00:03:13.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                    <SPLIT distance="100" swimtime="00:01:27.66" />
                    <SPLIT distance="150" swimtime="00:02:15.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="145" swimtime="00:00:47.97" resultid="1523" heatid="2040" lane="3" entrytime="00:00:47.32" entrycourse="SCM" />
                <RESULT eventid="1204" points="172" swimtime="00:01:41.47" resultid="1524" heatid="2020" lane="3" entrytime="00:01:49.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaleo" lastname="Bruno Da Luz" birthdate="2014-03-11" gender="M" nation="BRA" license="406658" swrid="4740124" athleteid="1580" externalid="406658" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1115" points="15" swimtime="00:01:40.90" resultid="1581" heatid="1985" lane="3" />
                <RESULT eventid="1283" points="53" swimtime="00:00:53.39" resultid="1582" heatid="2057" lane="1" entrytime="00:01:07.30" entrycourse="SCM" />
                <RESULT eventid="1239" points="35" swimtime="00:01:07.06" resultid="1583" heatid="2041" lane="5" entrytime="00:01:18.70" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Lima Belo" birthdate="2012-10-07" gender="F" nation="BRA" license="407799" athleteid="1596" externalid="407799">
              <RESULTS>
                <RESULT eventid="1118" points="84" swimtime="00:01:54.73" resultid="1597" heatid="1987" lane="5" />
                <RESULT eventid="1242" points="76" swimtime="00:02:09.45" resultid="1598" heatid="2042" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Faisal" lastname="Basem Ghotme" birthdate="2010-12-18" gender="M" nation="BRA" license="390809" swrid="5596871" athleteid="1550" externalid="390809" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1148" points="341" swimtime="00:02:31.05" resultid="1551" heatid="2000" lane="6" entrytime="00:02:32.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:12.92" />
                    <SPLIT distance="150" swimtime="00:01:52.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="393" swimtime="00:01:01.19" resultid="1552" heatid="1966" lane="2" entrytime="00:01:03.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="228" swimtime="00:01:30.37" resultid="1553" heatid="2064" lane="3" entrytime="00:01:31.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="331" swimtime="00:01:09.81" resultid="1554" heatid="2052" lane="1" entrytime="00:01:08.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="343" swimtime="00:02:21.91" resultid="1555" heatid="2034" lane="6" entrytime="00:02:24.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:09.99" />
                    <SPLIT distance="150" swimtime="00:01:46.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Oliveira" birthdate="2003-07-16" gender="M" nation="BRA" license="295723" swrid="5596944" athleteid="1440" externalid="295723" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1176" points="423" swimtime="00:01:03.62" resultid="1441" heatid="2010" lane="5" entrytime="00:00:59.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="435" swimtime="00:02:19.33" resultid="1442" heatid="2000" lane="3" entrytime="00:02:15.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:06.78" />
                    <SPLIT distance="150" swimtime="00:01:42.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="474" swimtime="00:00:57.48" resultid="1443" heatid="1968" lane="5" entrytime="00:00:57.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="418" swimtime="00:01:04.61" resultid="1444" heatid="2053" lane="4" entrytime="00:01:00.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="480" swimtime="00:02:06.88" resultid="1445" heatid="2036" lane="5" entrytime="00:02:05.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                    <SPLIT distance="100" swimtime="00:01:03.12" />
                    <SPLIT distance="150" swimtime="00:01:35.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabrizzio" lastname="Paolo Cazzola" birthdate="2009-06-15" gender="M" nation="BRA" license="357168" swrid="5596922" athleteid="1479" externalid="357168" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1148" points="300" swimtime="00:02:37.67" resultid="1480" heatid="1999" lane="3" entrytime="00:02:37.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                    <SPLIT distance="100" swimtime="00:01:16.84" />
                    <SPLIT distance="150" swimtime="00:01:57.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="326" swimtime="00:01:05.12" resultid="1481" heatid="1965" lane="4" entrytime="00:01:08.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="220" swimtime="00:01:31.56" resultid="1482" heatid="2064" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="283" swimtime="00:01:13.56" resultid="1483" heatid="2052" lane="6" entrytime="00:01:11.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="329" swimtime="00:02:23.85" resultid="1484" heatid="2034" lane="1" entrytime="00:02:24.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                    <SPLIT distance="100" swimtime="00:01:11.43" />
                    <SPLIT distance="150" swimtime="00:01:48.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Rogge" birthdate="2008-09-02" gender="M" nation="BRA" license="383387" swrid="4883279" athleteid="1428" externalid="383387" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1148" points="272" swimtime="00:02:42.85" resultid="1429" heatid="1999" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                    <SPLIT distance="100" swimtime="00:01:21.41" />
                    <SPLIT distance="150" swimtime="00:02:03.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="418" swimtime="00:00:59.94" resultid="1430" heatid="1968" lane="6" entrytime="00:00:58.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="244" swimtime="00:01:28.42" resultid="1431" heatid="2063" lane="2" />
                <RESULT eventid="1272" points="311" swimtime="00:01:11.33" resultid="1432" heatid="2052" lane="2" entrytime="00:01:07.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="319" swimtime="00:02:25.43" resultid="1433" heatid="2034" lane="4" entrytime="00:02:18.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="100" swimtime="00:01:10.07" />
                    <SPLIT distance="150" swimtime="00:01:48.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Leticia Sbardelatti" birthdate="2011-07-28" gender="F" nation="BRA" license="403147" swrid="5676303" athleteid="1566" externalid="403147" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1060" points="193" swimtime="00:01:26.84" resultid="1567" heatid="1960" lane="1" entrytime="00:01:31.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="114" swimtime="00:01:53.18" resultid="1568" heatid="2047" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="155" swimtime="00:03:25.02" resultid="1569" heatid="2027" lane="1" entrytime="00:04:10.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.37" />
                    <SPLIT distance="100" swimtime="00:01:38.66" />
                    <SPLIT distance="150" swimtime="00:02:32.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Carolina Ghellere" birthdate="2007-06-05" gender="F" nation="BRA" license="312662" swrid="5596874" athleteid="1426" externalid="312662" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1092" points="397" swimtime="00:03:03.03" resultid="1427" heatid="1976" lane="3" entrytime="00:02:48.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.03" />
                    <SPLIT distance="100" swimtime="00:01:28.74" />
                    <SPLIT distance="150" swimtime="00:02:15.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agata" lastname="Zacarias" birthdate="2014-08-05" gender="F" nation="BRA" license="387660" swrid="5596950" athleteid="1540" externalid="387660" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1112" points="139" swimtime="00:00:54.64" resultid="1541" heatid="1984" lane="5" entrytime="00:01:03.16" entrycourse="SCM" />
                <RESULT eventid="1080" points="149" swimtime="00:03:27.65" resultid="1542" heatid="1970" lane="2" entrytime="00:03:23.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.83" />
                    <SPLIT distance="100" swimtime="00:01:37.28" />
                    <SPLIT distance="150" swimtime="00:02:32.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="150" swimtime="00:00:43.10" resultid="1543" heatid="2055" lane="4" entrytime="00:00:41.19" entrycourse="SCM" />
                <RESULT eventid="1204" points="148" swimtime="00:01:46.70" resultid="1544" heatid="2019" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Resende Ames" birthdate="2006-02-10" gender="M" nation="BRA" license="365657" swrid="5596931" athleteid="1446" externalid="365657" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1176" points="489" swimtime="00:01:00.63" resultid="1447" heatid="2010" lane="2" entrytime="00:00:59.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="450" swimtime="00:02:17.80" resultid="1448" heatid="1999" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:07.04" />
                    <SPLIT distance="150" swimtime="00:01:42.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="525" swimtime="00:00:55.57" resultid="1449" heatid="1968" lane="2" entrytime="00:00:54.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="334" swimtime="00:01:09.63" resultid="1450" heatid="2053" lane="6" entrytime="00:01:05.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="554" swimtime="00:02:10.08" resultid="1451" heatid="2046" lane="3" entrytime="00:02:10.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                    <SPLIT distance="100" swimtime="00:01:01.98" />
                    <SPLIT distance="150" swimtime="00:01:35.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Riam Nagorski De Lima" birthdate="2014-04-26" gender="M" nation="BRA" license="407802" athleteid="1606" externalid="407802">
              <RESULTS>
                <RESULT eventid="1115" points="36" swimtime="00:01:15.07" resultid="1607" heatid="1985" lane="2" />
                <RESULT eventid="1283" points="46" swimtime="00:00:56.21" resultid="1608" heatid="2056" lane="2" />
                <RESULT eventid="1239" points="37" swimtime="00:01:05.86" resultid="1609" heatid="2041" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrieli" lastname="Brietzke Sbardelatti" birthdate="2014-07-14" gender="F" nation="BRA" license="400456" swrid="4379861" athleteid="1556" externalid="400456" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1112" points="123" swimtime="00:00:56.93" resultid="1557" heatid="1984" lane="1" entrytime="00:01:03.92" entrycourse="SCM" />
                <RESULT eventid="1080" points="161" swimtime="00:03:22.61" resultid="1558" heatid="1970" lane="6" entrytime="00:03:40.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.00" />
                    <SPLIT distance="100" swimtime="00:01:36.10" />
                    <SPLIT distance="150" swimtime="00:02:32.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="156" swimtime="00:00:42.59" resultid="1559" heatid="2055" lane="6" entrytime="00:00:45.01" entrycourse="SCM" />
                <RESULT eventid="1204" points="140" swimtime="00:01:48.59" resultid="1560" heatid="2019" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Laura Lima Belo" birthdate="2015-07-09" gender="F" nation="BRA" license="407801" athleteid="1603" externalid="407801">
              <RESULTS>
                <RESULT eventid="1280" points="31" swimtime="00:01:12.23" resultid="1604" heatid="2054" lane="5" />
                <RESULT eventid="1236" points="37" swimtime="00:01:15.60" resultid="1605" heatid="2039" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Kasprzak" birthdate="2011-08-09" gender="F" nation="BRA" license="406659" swrid="5073376" athleteid="1584" externalid="406659" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1060" points="133" swimtime="00:01:38.38" resultid="1585" heatid="1960" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" points="140" swimtime="00:01:59.93" resultid="1586" heatid="2061" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="96" swimtime="00:01:59.76" resultid="1587" heatid="2048" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Christopher" lastname="De Araujo" birthdate="2008-08-09" gender="M" nation="BRA" license="366376" swrid="5596884" athleteid="1462" externalid="366376" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1176" points="362" swimtime="00:01:07.01" resultid="1463" heatid="2007" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="488" swimtime="00:09:23.16" resultid="1464" heatid="1995" lane="1" />
                <RESULT eventid="1100" points="406" swimtime="00:02:42.20" resultid="1465" heatid="1980" lane="3" entrytime="00:02:34.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                    <SPLIT distance="100" swimtime="00:01:17.78" />
                    <SPLIT distance="150" swimtime="00:01:59.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="455" swimtime="00:01:11.85" resultid="1466" heatid="2066" lane="4" entrytime="00:01:12.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="425" swimtime="00:05:12.29" resultid="1467" heatid="2017" lane="2" entrytime="00:04:53.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                    <SPLIT distance="100" swimtime="00:01:12.60" />
                    <SPLIT distance="150" swimtime="00:01:55.15" />
                    <SPLIT distance="200" swimtime="00:02:36.10" />
                    <SPLIT distance="250" swimtime="00:03:19.02" />
                    <SPLIT distance="300" swimtime="00:04:01.60" />
                    <SPLIT distance="350" swimtime="00:04:38.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katherine" lastname="Kotz" birthdate="2012-05-18" gender="F" nation="BRA" license="390810" swrid="5596907" athleteid="1509" externalid="390810" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1118" points="288" swimtime="00:01:16.04" resultid="1510" heatid="1987" lane="3" entrytime="00:01:17.01" entrycourse="SCM" />
                <RESULT eventid="1086" points="243" swimtime="00:03:15.05" resultid="1511" heatid="1972" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.51" />
                    <SPLIT distance="100" swimtime="00:01:35.22" />
                    <SPLIT distance="150" swimtime="00:02:31.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="235" swimtime="00:00:45.93" resultid="1512" heatid="2058" lane="3" entrytime="00:00:49.25" entrycourse="SCM" />
                <RESULT eventid="1210" points="256" swimtime="00:06:03.87" resultid="1513" heatid="2023" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Ioris Souza" birthdate="2015-09-10" gender="F" nation="BRA" license="406693" swrid="5042791" athleteid="1588" externalid="406693" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1112" points="89" swimtime="00:01:03.44" resultid="1589" heatid="1983" lane="3" entrytime="00:01:12.58" entrycourse="SCM" />
                <RESULT eventid="1280" points="80" swimtime="00:00:53.17" resultid="1590" heatid="2054" lane="4" entrytime="00:01:00.61" entrycourse="SCM" />
                <RESULT eventid="1236" points="76" swimtime="00:00:59.39" resultid="1591" heatid="2040" lane="2" entrytime="00:01:06.75" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Roza" birthdate="2013-06-05" gender="M" nation="BRA" license="374412" swrid="5588949" athleteid="1525" externalid="374412" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1165" points="164" swimtime="00:00:39.66" resultid="1526" heatid="2004" lane="3" entrytime="00:00:37.58" entrycourse="SCM" />
                <RESULT eventid="1121" points="214" swimtime="00:01:14.85" resultid="1527" heatid="1989" lane="4" entrytime="00:01:16.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1245" status="DSQ" swimtime="00:01:36.06" resultid="1528" heatid="2043" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="178" swimtime="00:06:16.64" resultid="1529" heatid="2025" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Resende Ames" birthdate="2010-02-02" gender="M" nation="BRA" license="365505" swrid="5588876" athleteid="1514" externalid="365505" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1176" points="272" swimtime="00:01:13.70" resultid="1515" heatid="2009" lane="1" entrytime="00:01:13.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="400" swimtime="00:02:23.28" resultid="1516" heatid="2000" lane="5" entrytime="00:02:25.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                    <SPLIT distance="100" swimtime="00:01:09.60" />
                    <SPLIT distance="150" swimtime="00:01:47.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" status="DSQ" swimtime="00:01:03.23" resultid="1517" heatid="1966" lane="4" entrytime="00:01:02.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="368" swimtime="00:01:07.39" resultid="1518" heatid="2052" lane="4" entrytime="00:01:06.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="343" swimtime="00:02:21.84" resultid="1519" heatid="2035" lane="5" entrytime="00:02:14.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="100" swimtime="00:01:08.45" />
                    <SPLIT distance="150" swimtime="00:01:45.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edward" lastname="Mikael De Lima" birthdate="2012-03-11" gender="M" nation="BRA" license="376445" swrid="5588816" athleteid="1530" externalid="376445" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1121" points="316" swimtime="00:01:05.83" resultid="1531" heatid="1988" lane="3" entrytime="00:01:28.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1089" points="252" swimtime="00:02:53.34" resultid="1532" heatid="1974" lane="3" entrytime="00:02:43.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:17.07" />
                    <SPLIT distance="150" swimtime="00:02:11.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1245" points="259" swimtime="00:01:15.76" resultid="1533" heatid="2043" lane="3" entrytime="00:01:19.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:05.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="358" swimtime="00:04:58.78" resultid="1534" heatid="2025" lane="3" entrytime="00:05:28.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Targat Pinheiro" birthdate="2008-09-04" gender="F" nation="BRA" license="331610" swrid="5596894" athleteid="1420" externalid="331610" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="1421" heatid="2006" lane="3" entrytime="00:01:12.03" entrycourse="SCM" />
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="1422" heatid="1992" lane="4" entrytime="00:10:21.73" entrycourse="SCM" />
                <RESULT eventid="1264" status="DNS" swimtime="00:00:00.00" resultid="1423" heatid="2049" lane="4" entrytime="00:01:15.44" entrycourse="SCM" />
                <RESULT eventid="1216" status="DNS" swimtime="00:00:00.00" resultid="1424" heatid="2030" lane="2" entrytime="00:02:24.50" entrycourse="SCM" />
                <RESULT eventid="1184" status="DNS" swimtime="00:00:00.00" resultid="1425" heatid="2013" lane="5" entrytime="00:05:45.57" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Gabriel Dreher" birthdate="2011-12-05" gender="M" nation="BRA" license="403148" swrid="5676302" athleteid="1570" externalid="403148" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1068" points="116" swimtime="00:01:31.80" resultid="1571" heatid="1964" lane="5" entrytime="00:01:35.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="83" swimtime="00:01:50.43" resultid="1572" heatid="2050" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="103" swimtime="00:03:31.93" resultid="1573" heatid="2032" lane="5" entrytime="00:03:44.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.46" />
                    <SPLIT distance="100" swimtime="00:01:46.59" />
                    <SPLIT distance="150" swimtime="00:02:43.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Luiz Martinazzo" birthdate="2006-05-16" gender="M" nation="BRA" license="345593" swrid="5596910" athleteid="1457" externalid="345593" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1148" points="378" swimtime="00:02:25.99" resultid="1458" heatid="2000" lane="2" entrytime="00:02:19.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                    <SPLIT distance="100" swimtime="00:01:10.21" />
                    <SPLIT distance="150" swimtime="00:01:48.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="475" swimtime="00:00:57.44" resultid="1459" heatid="1967" lane="3" entrytime="00:00:58.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="391" swimtime="00:01:06.08" resultid="1460" heatid="2053" lane="5" entrytime="00:01:03.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="483" swimtime="00:02:06.58" resultid="1461" heatid="2036" lane="2" entrytime="00:02:04.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                    <SPLIT distance="100" swimtime="00:01:02.02" />
                    <SPLIT distance="150" swimtime="00:01:34.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Axel" lastname="Ariel Giménez González" birthdate="2011-06-01" gender="M" nation="BRA" license="365755" swrid="5676299" athleteid="1574" externalid="365755" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1100" points="219" swimtime="00:03:19.34" resultid="1575" heatid="1977" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.54" />
                    <SPLIT distance="100" swimtime="00:01:39.63" />
                    <SPLIT distance="150" swimtime="00:02:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="281" swimtime="00:01:08.45" resultid="1576" heatid="1965" lane="2" entrytime="00:01:09.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="211" swimtime="00:01:32.75" resultid="1577" heatid="2063" lane="4" />
                <RESULT eventid="1272" points="193" swimtime="00:01:23.61" resultid="1578" heatid="2050" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="260" swimtime="00:02:35.54" resultid="1579" heatid="2033" lane="1" entrytime="00:02:40.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                    <SPLIT distance="100" swimtime="00:01:15.10" />
                    <SPLIT distance="150" swimtime="00:01:57.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="De Souza Tulio" birthdate="2006-06-23" gender="F" nation="BRA" license="342344" swrid="5030980" athleteid="1434" externalid="342344" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1140" points="460" swimtime="00:02:34.01" resultid="1435" heatid="1998" lane="3" entrytime="00:02:23.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                    <SPLIT distance="100" swimtime="00:01:13.03" />
                    <SPLIT distance="150" swimtime="00:01:53.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="517" swimtime="00:01:02.58" resultid="1436" heatid="1962" lane="3" entrytime="00:00:58.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1292" status="DSQ" swimtime="00:01:29.78" resultid="1437" heatid="2061" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="413" swimtime="00:01:13.66" resultid="1438" heatid="2049" lane="3" entrytime="00:01:05.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="534" swimtime="00:02:15.92" resultid="1439" heatid="2030" lane="3" entrytime="00:02:07.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:05.94" />
                    <SPLIT distance="150" swimtime="00:01:40.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ysadora" lastname="Bertoldo" birthdate="2010-04-09" gender="F" nation="BRA" license="376444" swrid="5588553" athleteid="1503" externalid="376444" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1168" points="236" swimtime="00:01:27.42" resultid="1504" heatid="2005" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="406" swimtime="00:10:44.68" resultid="1505" heatid="1992" lane="6" entrytime="00:11:12.78" entrycourse="SCM" />
                <RESULT eventid="1060" points="329" swimtime="00:01:12.73" resultid="1506" heatid="1961" lane="6" entrytime="00:01:13.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="274" swimtime="00:01:24.46" resultid="1507" heatid="2047" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="374" swimtime="00:02:33.05" resultid="1508" heatid="2028" lane="3" entrytime="00:02:34.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                    <SPLIT distance="100" swimtime="00:01:16.80" />
                    <SPLIT distance="150" swimtime="00:01:56.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="De Assis Santos" birthdate="2003-02-21" gender="M" nation="BRA" license="342496" swrid="5596885" athleteid="1452" externalid="342496" level="INTERNE/IT">
              <RESULTS>
                <RESULT eventid="1176" points="299" swimtime="00:01:11.45" resultid="1453" heatid="2009" lane="4" entrytime="00:01:07.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="386" swimtime="00:02:25.00" resultid="1454" heatid="2000" lane="4" entrytime="00:02:18.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:09.54" />
                    <SPLIT distance="150" swimtime="00:01:47.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="396" swimtime="00:01:05.80" resultid="1455" heatid="2053" lane="2" entrytime="00:01:02.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="384" swimtime="00:02:16.66" resultid="1456" heatid="2032" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="100" swimtime="00:01:05.14" />
                    <SPLIT distance="150" swimtime="00:01:41.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="De Souza" birthdate="2014-03-30" gender="M" nation="BRA" license="407800" athleteid="1599" externalid="407800">
              <RESULTS>
                <RESULT eventid="1115" points="109" swimtime="00:00:52.20" resultid="1600" heatid="1985" lane="4" />
                <RESULT eventid="1283" points="78" swimtime="00:00:47.16" resultid="1601" heatid="2056" lane="3" />
                <RESULT eventid="1239" points="63" swimtime="00:00:55.40" resultid="1602" heatid="2041" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Kaiser" birthdate="2014-06-02" gender="F" nation="BRA" license="407883" athleteid="1610" externalid="407883">
              <RESULTS>
                <RESULT eventid="1280" points="29" swimtime="00:01:14.62" resultid="1611" heatid="2054" lane="1" />
                <RESULT eventid="1236" points="49" swimtime="00:01:08.86" resultid="1612" heatid="2039" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Bailke" birthdate="2007-05-04" gender="M" nation="BRA" license="370566" swrid="5596869" athleteid="1468" externalid="370566" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1176" points="269" swimtime="00:01:13.98" resultid="1469" heatid="2009" lane="5" entrytime="00:01:12.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="359" swimtime="00:10:23.46" resultid="1470" heatid="1996" lane="6" entrytime="00:10:33.53" entrycourse="SCM" />
                <RESULT eventid="1068" points="370" swimtime="00:01:02.45" resultid="1471" heatid="1966" lane="3" entrytime="00:01:02.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="232" swimtime="00:02:53.80" resultid="1472" heatid="2046" lane="1" entrytime="00:02:51.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="100" swimtime="00:01:19.05" />
                    <SPLIT distance="150" swimtime="00:02:06.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="375" swimtime="00:02:17.75" resultid="1473" heatid="2035" lane="1" entrytime="00:02:15.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                    <SPLIT distance="100" swimtime="00:01:08.21" />
                    <SPLIT distance="150" swimtime="00:01:42.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Paulo Sales" birthdate="2007-11-07" gender="M" nation="BRA" license="390712" swrid="5596923" athleteid="1491" externalid="390712" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1176" points="220" swimtime="00:01:19.07" resultid="1492" heatid="2007" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="241" swimtime="00:03:13.08" resultid="1493" heatid="1979" lane="5" entrytime="00:03:11.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.35" />
                    <SPLIT distance="100" swimtime="00:01:30.97" />
                    <SPLIT distance="150" swimtime="00:02:21.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="314" swimtime="00:01:05.91" resultid="1494" heatid="1965" lane="3" entrytime="00:01:08.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="227" swimtime="00:01:30.61" resultid="1495" heatid="2065" lane="5" entrytime="00:01:28.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="278" swimtime="00:02:32.10" resultid="1496" heatid="2031" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                    <SPLIT distance="100" swimtime="00:01:14.50" />
                    <SPLIT distance="150" swimtime="00:01:53.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alessandro" lastname="Cazzola" birthdate="2014-09-15" gender="M" nation="PRY" license="390713" athleteid="1545" externalid="390713" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1115" points="145" swimtime="00:00:47.47" resultid="1546" heatid="1986" lane="3" entrytime="00:00:48.22" entrycourse="SCM" />
                <RESULT eventid="1083" points="143" swimtime="00:03:09.89" resultid="1547" heatid="1971" lane="4" entrytime="00:03:18.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                    <SPLIT distance="100" swimtime="00:01:30.09" />
                    <SPLIT distance="150" swimtime="00:02:19.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1283" points="150" swimtime="00:00:37.86" resultid="1548" heatid="2057" lane="4" entrytime="00:00:37.83" entrycourse="SCM" />
                <RESULT eventid="1207" points="140" swimtime="00:01:34.90" resultid="1549" heatid="2022" lane="4" entrytime="00:01:58.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joshua" lastname="Davalos Gimenez" birthdate="2013-10-22" gender="M" nation="PRY" license="380598" athleteid="1535" externalid="380598" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1121" points="207" swimtime="00:01:15.72" resultid="1536" heatid="1989" lane="2" entrytime="00:01:19.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1089" points="167" swimtime="00:03:18.69" resultid="1537" heatid="1974" lane="1" entrytime="00:03:19.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.93" />
                    <SPLIT distance="100" swimtime="00:01:42.30" />
                    <SPLIT distance="150" swimtime="00:02:36.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1289" points="173" swimtime="00:00:44.72" resultid="1538" heatid="2060" lane="4" entrytime="00:00:44.88" entrycourse="SCM" />
                <RESULT eventid="1213" points="214" swimtime="00:05:54.61" resultid="1539" heatid="2025" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Marques Petry" birthdate="2008-01-08" gender="M" nation="BRA" license="392352" swrid="4795316" athleteid="1497" externalid="392352" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1148" points="264" swimtime="00:02:44.53" resultid="1498" heatid="1999" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.59" />
                    <SPLIT distance="100" swimtime="00:01:21.75" />
                    <SPLIT distance="150" swimtime="00:02:04.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="270" swimtime="00:03:05.72" resultid="1499" heatid="1979" lane="4" entrytime="00:03:08.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                    <SPLIT distance="100" swimtime="00:01:29.78" />
                    <SPLIT distance="150" swimtime="00:02:18.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="361" swimtime="00:01:02.94" resultid="1500" heatid="1966" lane="5" entrytime="00:01:03.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1300" points="265" swimtime="00:01:25.96" resultid="1501" heatid="2065" lane="3" entrytime="00:01:24.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="351" swimtime="00:02:20.84" resultid="1502" heatid="2034" lane="2" entrytime="00:02:20.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:10.14" />
                    <SPLIT distance="150" swimtime="00:01:46.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
