<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.79911">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Cascavel" name="Torneio Regional da 3ª Região (Pré-Mirim/Sênior)" course="SCM" deadline="2024-07-22" entrystartdate="2024-07-16" entrytype="INVITATION" hostclub="Associação Atlética Comercial" hostclub.url="https://www.clubecomercial.net.br/" number="38315" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/newInterface/eventos/38315" startmethod="1" timing="AUTOMATIC" touchpad="ONESIDE" masters="F" withdrawuntil="2024-07-25" state="PR" nation="BRA">
      <AGEDATE value="2024-01-01" type="YEAR" />
      <POOL name="Associação Atlética Comercial" lanemin="1" lanemax="6" />
      <FACILITY city="Cascavel" name="Associação Atlética Comercial" nation="BRA" state="PR" street="Rua Recife, 2563" street2="Bairro Coqueiral" zip="85807-060" />
      <POINTTABLE pointtableid="3016" name="FINA Point Scoring" version="2023" />
      <QUALIFY from="2023-07-28" until="2024-07-27" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99233-1025" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99233-1025" street="Avenida do Batel, 1230" street2="Batel" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-07-28" daytime="09:10" endtime="12:52" number="1">
          <EVENTS>
            <EVENT eventid="1060" daytime="09:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1711" />
                    <RANKING order="2" place="2" resultid="1804" />
                    <RANKING order="3" place="3" resultid="1831" />
                    <RANKING order="4" place="4" resultid="1745" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1064" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1065" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1625" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1067" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1638" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2002" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2003" daytime="09:14" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1068" daytime="09:18" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1069" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1676" />
                    <RANKING order="2" place="2" resultid="1699" />
                    <RANKING order="3" place="3" resultid="1682" />
                    <RANKING order="4" place="4" resultid="1717" />
                    <RANKING order="5" place="5" resultid="1815" />
                    <RANKING order="6" place="-1" resultid="1778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1751" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1072" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1757" />
                    <RANKING order="2" place="2" resultid="1471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1445" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1449" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2004" daytime="09:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2005" daytime="09:22" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1076" daytime="09:26" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1077" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1599" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1480" />
                    <RANKING order="2" place="2" resultid="1799" />
                    <RANKING order="3" place="3" resultid="1874" />
                    <RANKING order="4" place="-1" resultid="1569" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2006" daytime="09:26" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1079" daytime="09:30" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1080" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1768" />
                    <RANKING order="2" place="2" resultid="1398" />
                    <RANKING order="3" place="3" resultid="1884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1826" />
                    <RANKING order="2" place="2" resultid="1688" />
                    <RANKING order="3" place="3" resultid="1437" />
                    <RANKING order="4" place="4" resultid="1810" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2007" daytime="09:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2008" daytime="09:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1082" daytime="09:36" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1083" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1406" />
                    <RANKING order="2" place="2" resultid="1560" />
                    <RANKING order="3" place="3" resultid="1928" />
                    <RANKING order="4" place="-1" resultid="1594" />
                    <RANKING order="5" place="-1" resultid="1784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1773" />
                    <RANKING order="2" place="2" resultid="1863" />
                    <RANKING order="3" place="3" resultid="1789" />
                    <RANKING order="4" place="4" resultid="1735" />
                    <RANKING order="5" place="5" resultid="1430" />
                    <RANKING order="6" place="6" resultid="1896" />
                    <RANKING order="7" place="7" resultid="1418" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2009" daytime="09:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2010" daytime="09:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1085" daytime="09:42" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1086" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1410" />
                    <RANKING order="2" place="2" resultid="1879" />
                    <RANKING order="3" place="3" resultid="1900" />
                    <RANKING order="4" place="4" resultid="1932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1573" />
                    <RANKING order="2" place="2" resultid="1740" />
                    <RANKING order="3" place="3" resultid="1905" />
                    <RANKING order="4" place="4" resultid="1853" />
                    <RANKING order="5" place="5" resultid="1581" />
                    <RANKING order="6" place="6" resultid="1892" />
                    <RANKING order="7" place="7" resultid="1910" />
                    <RANKING order="8" place="-1" resultid="1426" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2011" daytime="09:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2012" daytime="09:44" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1088" daytime="09:48" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1089" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1705" />
                    <RANKING order="2" place="2" resultid="1712" />
                    <RANKING order="3" place="3" resultid="1979" />
                    <RANKING order="4" place="4" resultid="1832" />
                    <RANKING order="5" place="5" resultid="1973" />
                    <RANKING order="6" place="6" resultid="1357" />
                    <RANKING order="7" place="7" resultid="1746" />
                    <RANKING order="8" place="8" resultid="1535" />
                    <RANKING order="9" place="9" resultid="1551" />
                    <RANKING order="10" place="10" resultid="1991" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1646" />
                    <RANKING order="2" place="2" resultid="1837" />
                    <RANKING order="3" place="3" resultid="1321" />
                    <RANKING order="4" place="4" resultid="1961" />
                    <RANKING order="5" place="5" resultid="1968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1361" />
                    <RANKING order="2" place="2" resultid="1633" />
                    <RANKING order="3" place="3" resultid="1464" />
                    <RANKING order="4" place="-1" resultid="1652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1092" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1325" />
                    <RANKING order="2" place="2" resultid="1949" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1621" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2013" daytime="09:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2014" daytime="09:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2015" daytime="09:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2016" daytime="09:54" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1096" daytime="09:58" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1097" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1677" />
                    <RANKING order="2" place="2" resultid="1683" />
                    <RANKING order="3" place="3" resultid="1546" />
                    <RANKING order="4" place="4" resultid="1779" />
                    <RANKING order="5" place="5" resultid="1530" />
                    <RANKING order="6" place="6" resultid="1378" />
                    <RANKING order="7" place="7" resultid="1816" />
                    <RANKING order="8" place="8" resultid="1402" />
                    <RANKING order="9" place="9" resultid="1394" />
                    <RANKING order="10" place="10" resultid="1997" />
                    <RANKING order="11" place="11" resultid="1414" />
                    <RANKING order="12" place="12" resultid="1914" />
                    <RANKING order="13" place="13" resultid="1540" />
                    <RANKING order="14" place="-1" resultid="1985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1658" />
                    <RANKING order="2" place="2" resultid="1510" />
                    <RANKING order="3" place="3" resultid="1752" />
                    <RANKING order="4" place="4" resultid="1664" />
                    <RANKING order="5" place="5" resultid="1868" />
                    <RANKING order="6" place="6" resultid="1919" />
                    <RANKING order="7" place="-1" resultid="1485" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1723" />
                    <RANKING order="2" place="2" resultid="1642" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1442" />
                    <RANKING order="2" place="2" resultid="1758" />
                    <RANKING order="3" place="3" resultid="1346" />
                    <RANKING order="4" place="4" resultid="1729" />
                    <RANKING order="5" place="5" resultid="1937" />
                    <RANKING order="6" place="6" resultid="1472" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1350" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1454" />
                    <RANKING order="2" place="2" resultid="1615" />
                    <RANKING order="3" place="3" resultid="1955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1336" />
                    <RANKING order="2" place="2" resultid="1329" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2017" daytime="09:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2018" daytime="10:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2019" daytime="10:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2020" daytime="10:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2021" daytime="10:06" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2022" daytime="10:08" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1104" daytime="10:10" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1105" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1373" />
                    <RANKING order="2" place="2" resultid="1589" />
                    <RANKING order="3" place="3" resultid="1858" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1481" />
                    <RANKING order="2" place="2" resultid="1794" />
                    <RANKING order="3" place="3" resultid="1570" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2023" daytime="10:10" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1107" daytime="10:18" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1108" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1495" />
                    <RANKING order="2" place="2" resultid="1556" />
                    <RANKING order="3" place="-1" resultid="1515" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1500" />
                    <RANKING order="2" place="2" resultid="1689" />
                    <RANKING order="3" place="3" resultid="1763" />
                    <RANKING order="4" place="4" resultid="1525" />
                    <RANKING order="5" place="5" resultid="1811" />
                    <RANKING order="6" place="6" resultid="1585" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2024" daytime="10:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2025" daytime="10:22" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1110" daytime="10:26" gender="F" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1111" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1407" />
                    <RANKING order="2" place="2" resultid="1561" />
                    <RANKING order="3" place="3" resultid="1578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1112" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1821" />
                    <RANKING order="2" place="2" resultid="1490" />
                    <RANKING order="3" place="3" resultid="1520" />
                    <RANKING order="4" place="4" resultid="1774" />
                    <RANKING order="5" place="5" resultid="1864" />
                    <RANKING order="6" place="6" resultid="1790" />
                    <RANKING order="7" place="7" resultid="1431" />
                    <RANKING order="8" place="8" resultid="1924" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2026" daytime="10:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2027" daytime="10:30" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1113" daytime="10:34" gender="M" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1114" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1848" />
                    <RANKING order="2" place="2" resultid="1880" />
                    <RANKING order="3" place="3" resultid="1411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1741" />
                    <RANKING order="2" place="2" resultid="1854" />
                    <RANKING order="3" place="3" resultid="1390" />
                    <RANKING order="4" place="4" resultid="1843" />
                    <RANKING order="5" place="5" resultid="1574" />
                    <RANKING order="6" place="6" resultid="1906" />
                    <RANKING order="7" place="7" resultid="1888" />
                    <RANKING order="8" place="8" resultid="1582" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2028" daytime="10:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2029" daytime="10:36" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1116" daytime="10:54" gender="F" number="13" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1117" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1805" />
                    <RANKING order="2" place="2" resultid="1974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1476" />
                    <RANKING order="2" place="2" resultid="1505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1120" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1343" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1122" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1123" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2030" daytime="10:54" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1124" daytime="11:18" gender="M" number="14" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1125" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1718" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1127" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1643" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1131" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1610" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2031" daytime="11:18" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1132" daytime="11:40" gender="F" number="15" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1133" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1358" />
                    <RANKING order="2" place="2" resultid="1992" />
                    <RANKING order="3" place="3" resultid="1552" />
                    <RANKING order="4" place="-1" resultid="1339" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1134" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1962" />
                    <RANKING order="2" place="2" resultid="1838" />
                    <RANKING order="3" place="3" resultid="1365" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1634" />
                    <RANKING order="2" place="2" resultid="1362" />
                    <RANKING order="3" place="-1" resultid="1653" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1137" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1138" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1326" />
                    <RANKING order="2" place="2" resultid="1950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1139" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1943" />
                    <RANKING order="2" place="2" resultid="1622" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2032" daytime="11:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2033" daytime="11:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2034" daytime="11:44" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1140" daytime="11:48" gender="M" number="16" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1141" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1678" />
                    <RANKING order="2" place="2" resultid="1379" />
                    <RANKING order="3" place="3" resultid="1541" />
                    <RANKING order="4" place="4" resultid="1998" />
                    <RANKING order="5" place="-1" resultid="1986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1659" />
                    <RANKING order="2" place="-1" resultid="1486" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1143" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1144" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1671" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1455" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1332" />
                    <RANKING order="2" place="2" resultid="1450" />
                    <RANKING order="3" place="3" resultid="1611" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2035" daytime="11:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2036" daytime="11:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2037" daytime="11:52" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1148" daytime="11:54" gender="F" number="17" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1149" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1600" />
                    <RANKING order="2" place="2" resultid="1374" />
                    <RANKING order="3" place="3" resultid="1590" />
                    <RANKING order="4" place="4" resultid="1386" />
                    <RANKING order="5" place="5" resultid="1859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1800" />
                    <RANKING order="2" place="2" resultid="1795" />
                    <RANKING order="3" place="3" resultid="1875" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2038" daytime="11:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2039" daytime="11:58" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1151" daytime="12:00" gender="M" number="18" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1152" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1769" />
                    <RANKING order="2" place="2" resultid="1382" />
                    <RANKING order="3" place="3" resultid="1557" />
                    <RANKING order="4" place="4" resultid="1399" />
                    <RANKING order="5" place="5" resultid="1885" />
                    <RANKING order="6" place="-1" resultid="1496" />
                    <RANKING order="7" place="-1" resultid="1516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1764" />
                    <RANKING order="2" place="2" resultid="1827" />
                    <RANKING order="3" place="3" resultid="1438" />
                    <RANKING order="4" place="4" resultid="1526" />
                    <RANKING order="5" place="5" resultid="1586" />
                    <RANKING order="6" place="6" resultid="1434" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2040" daytime="12:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2041" daytime="12:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2042" daytime="12:06" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1154" daytime="12:08" gender="F" number="19" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1155" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1929" />
                    <RANKING order="2" place="-1" resultid="1595" />
                    <RANKING order="3" place="-1" resultid="1785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1491" />
                    <RANKING order="2" place="2" resultid="1822" />
                    <RANKING order="3" place="3" resultid="1521" />
                    <RANKING order="4" place="4" resultid="1736" />
                    <RANKING order="5" place="5" resultid="1925" />
                    <RANKING order="6" place="6" resultid="1897" />
                    <RANKING order="7" place="7" resultid="1419" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2043" daytime="12:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2044" daytime="12:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1157" daytime="12:14" gender="M" number="20" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1158" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1849" />
                    <RANKING order="2" place="2" resultid="1901" />
                    <RANKING order="3" place="3" resultid="1933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1844" />
                    <RANKING order="2" place="2" resultid="1889" />
                    <RANKING order="3" place="3" resultid="1893" />
                    <RANKING order="4" place="4" resultid="1911" />
                    <RANKING order="5" place="-1" resultid="1427" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2045" daytime="12:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2046" daytime="12:16" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1160" daytime="12:18" gender="F" number="21" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1161" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1833" />
                    <RANKING order="2" place="2" resultid="1713" />
                    <RANKING order="3" place="3" resultid="1806" />
                    <RANKING order="4" place="4" resultid="1975" />
                    <RANKING order="5" place="5" resultid="1747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1162" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1647" />
                    <RANKING order="2" place="2" resultid="1369" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1163" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1164" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1165" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1167" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1944" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2047" daytime="12:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2048" daytime="12:22" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1168" daytime="12:24" gender="M" number="22" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1169" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1700" />
                    <RANKING order="2" place="2" resultid="1531" />
                    <RANKING order="3" place="3" resultid="1719" />
                    <RANKING order="4" place="4" resultid="1780" />
                    <RANKING order="5" place="5" resultid="1684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1753" />
                    <RANKING order="2" place="2" resultid="1665" />
                    <RANKING order="3" place="3" resultid="1511" />
                    <RANKING order="4" place="4" resultid="1869" />
                    <RANKING order="5" place="-1" resultid="1487" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1724" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1759" />
                    <RANKING order="2" place="2" resultid="1939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1174" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2049" daytime="12:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2050" daytime="12:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2051" daytime="12:30" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1176" daytime="12:32" gender="F" number="23" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1177" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1980" />
                    <RANKING order="2" place="2" resultid="1706" />
                    <RANKING order="3" place="3" resultid="1536" />
                    <RANKING order="4" place="4" resultid="1340" />
                    <RANKING order="5" place="5" resultid="1553" />
                    <RANKING order="6" place="6" resultid="1993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1969" />
                    <RANKING order="2" place="-1" resultid="1506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1180" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1181" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1182" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1183" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1639" />
                    <RANKING order="2" place="2" resultid="1945" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2052" daytime="12:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2053" daytime="12:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1184" daytime="12:36" gender="M" number="24" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1185" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1817" />
                    <RANKING order="2" place="2" resultid="1547" />
                    <RANKING order="3" place="3" resultid="1915" />
                    <RANKING order="4" place="4" resultid="1403" />
                    <RANKING order="5" place="5" resultid="1542" />
                    <RANKING order="6" place="6" resultid="1999" />
                    <RANKING order="7" place="-1" resultid="1987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1604" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1188" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1347" />
                    <RANKING order="2" place="2" resultid="1730" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1189" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1354" />
                    <RANKING order="2" place="2" resultid="1956" />
                    <RANKING order="3" place="3" resultid="1456" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2054" daytime="12:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2055" daytime="12:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2056" daytime="12:40" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-07-28" daytime="15:40" endtime="18:39" number="2">
          <EVENTS>
            <EVENT eventid="1192" daytime="15:40" gender="F" number="25" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1193" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1714" />
                    <RANKING order="2" place="2" resultid="1707" />
                    <RANKING order="3" place="3" resultid="1807" />
                    <RANKING order="4" place="4" resultid="1748" />
                    <RANKING order="5" place="5" resultid="1834" />
                    <RANKING order="6" place="6" resultid="1976" />
                    <RANKING order="7" place="7" resultid="1981" />
                    <RANKING order="8" place="8" resultid="1537" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1477" />
                    <RANKING order="2" place="2" resultid="1648" />
                    <RANKING order="3" place="3" resultid="1963" />
                    <RANKING order="4" place="4" resultid="1322" />
                    <RANKING order="5" place="5" resultid="1507" />
                    <RANKING order="6" place="6" resultid="1839" />
                    <RANKING order="7" place="7" resultid="1970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1635" />
                    <RANKING order="2" place="-1" resultid="1654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1196" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1695" />
                    <RANKING order="2" place="2" resultid="1344" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1197" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1628" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1199" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2057" daytime="15:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2058" daytime="15:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2059" daytime="15:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2060" daytime="16:02" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1200" daytime="16:08" gender="M" number="26" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1201" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1679" />
                    <RANKING order="2" place="2" resultid="1701" />
                    <RANKING order="3" place="3" resultid="1720" />
                    <RANKING order="4" place="4" resultid="1685" />
                    <RANKING order="5" place="5" resultid="1781" />
                    <RANKING order="6" place="6" resultid="1818" />
                    <RANKING order="7" place="7" resultid="1543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1660" />
                    <RANKING order="2" place="2" resultid="1754" />
                    <RANKING order="3" place="3" resultid="1666" />
                    <RANKING order="4" place="4" resultid="1870" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1203" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1644" />
                    <RANKING order="2" place="2" resultid="1725" />
                    <RANKING order="3" place="3" resultid="1605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1204" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1631" />
                    <RANKING order="2" place="2" resultid="1760" />
                    <RANKING order="3" place="3" resultid="1731" />
                    <RANKING order="4" place="4" resultid="1468" />
                    <RANKING order="5" place="5" resultid="1473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1205" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1673" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1206" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1617" />
                    <RANKING order="2" place="2" resultid="1457" />
                    <RANKING order="3" place="3" resultid="1446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1612" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2061" daytime="16:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2062" daytime="16:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2063" daytime="16:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2064" daytime="16:26" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1208" daytime="16:32" gender="F" number="27" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1209" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1210" daytime="16:32" gender="M" number="28" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1211" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1212" daytime="16:32" gender="F" number="29" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1213" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1562" />
                    <RANKING order="2" place="-1" resultid="1786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1492" />
                    <RANKING order="2" place="2" resultid="1823" />
                    <RANKING order="3" place="3" resultid="1522" />
                    <RANKING order="4" place="4" resultid="1775" />
                    <RANKING order="5" place="5" resultid="1737" />
                    <RANKING order="6" place="6" resultid="1865" />
                    <RANKING order="7" place="7" resultid="1791" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2065" daytime="16:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2066" daytime="16:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1215" daytime="16:38" gender="M" number="30" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1216" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1850" />
                    <RANKING order="2" place="2" resultid="1881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1742" />
                    <RANKING order="2" place="2" resultid="1855" />
                    <RANKING order="3" place="3" resultid="1391" />
                    <RANKING order="4" place="4" resultid="1907" />
                    <RANKING order="5" place="5" resultid="1845" />
                    <RANKING order="6" place="6" resultid="1575" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2067" daytime="16:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2068" daytime="16:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1218" daytime="16:42" gender="F" number="31" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1219" agemax="11" agemin="11" />
                <AGEGROUP agegroupid="1220" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1801" />
                    <RANKING order="2" place="2" resultid="1796" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2069" daytime="16:42" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1221" daytime="16:46" gender="M" number="32" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1222" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1223" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1501" />
                    <RANKING order="2" place="2" resultid="1690" />
                    <RANKING order="3" place="3" resultid="1765" />
                    <RANKING order="4" place="4" resultid="1812" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2070" daytime="16:46" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1224" daytime="16:50" gender="F" number="33" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1225" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1226" daytime="16:50" gender="M" number="34" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1227" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1565" />
                    <RANKING order="2" place="2" resultid="1422" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2071" daytime="16:50" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1228" daytime="16:52" gender="F" number="35" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1229" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1749" />
                    <RANKING order="2" place="2" resultid="1835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1232" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1696" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1234" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1235" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1640" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2072" daytime="16:52" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1236" daytime="16:54" gender="M" number="36" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1237" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1702" />
                    <RANKING order="2" place="2" resultid="1721" />
                    <RANKING order="3" place="3" resultid="1415" />
                    <RANKING order="4" place="4" resultid="2000" />
                    <RANKING order="5" place="-1" resultid="1548" />
                    <RANKING order="6" place="-1" resultid="1988" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1238" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1661" />
                    <RANKING order="2" place="2" resultid="1921" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1239" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1240" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1732" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1674" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1355" />
                    <RANKING order="2" place="2" resultid="1957" />
                    <RANKING order="3" place="3" resultid="1618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1243" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2073" daytime="16:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2074" daytime="16:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2075" daytime="17:00" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1244" daytime="17:18" gender="F" number="37" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1245" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1708" />
                    <RANKING order="2" place="2" resultid="1982" />
                    <RANKING order="3" place="3" resultid="1977" />
                    <RANKING order="4" place="4" resultid="1715" />
                    <RANKING order="5" place="-1" resultid="1994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1964" />
                    <RANKING order="2" place="2" resultid="1649" />
                    <RANKING order="3" place="3" resultid="1370" />
                    <RANKING order="4" place="4" resultid="1478" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1248" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1249" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1250" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1251" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1623" />
                    <RANKING order="2" place="2" resultid="1946" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2076" daytime="17:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2077" daytime="17:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2078" daytime="17:22" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1252" daytime="17:24" gender="M" number="38" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1253" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1532" />
                    <RANKING order="2" place="2" resultid="1819" />
                    <RANKING order="3" place="3" resultid="1395" />
                    <RANKING order="4" place="4" resultid="1916" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1254" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1667" />
                    <RANKING order="2" place="2" resultid="1871" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1255" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1726" />
                    <RANKING order="2" place="2" resultid="1606" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1256" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1940" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1257" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1351" />
                    <RANKING order="2" place="2" resultid="1461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1258" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1333" />
                    <RANKING order="2" place="2" resultid="1451" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2079" daytime="17:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2080" daytime="17:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2081" daytime="17:28" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1260" daytime="17:30" gender="F" number="39" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1261" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1262" daytime="17:30" gender="M" number="40" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1263" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1566" />
                    <RANKING order="2" place="2" resultid="1423" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2082" daytime="17:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1264" daytime="17:32" gender="F" number="41" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1265" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1601" />
                    <RANKING order="2" place="2" resultid="1375" />
                    <RANKING order="3" place="3" resultid="1387" />
                    <RANKING order="4" place="-1" resultid="1591" />
                    <RANKING order="5" place="-1" resultid="1860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1482" />
                    <RANKING order="2" place="2" resultid="1802" />
                    <RANKING order="3" place="3" resultid="1876" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2083" daytime="17:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2084" daytime="17:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1267" daytime="17:38" gender="M" number="42" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1268" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1770" />
                    <RANKING order="2" place="2" resultid="1383" />
                    <RANKING order="3" place="-1" resultid="1517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1269" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1502" />
                    <RANKING order="2" place="2" resultid="1527" />
                    <RANKING order="3" place="3" resultid="1828" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2085" daytime="17:38" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1270" daytime="17:42" gender="F" number="43" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1271" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1808" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1272" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1965" />
                    <RANKING order="2" place="2" resultid="1371" />
                    <RANKING order="3" place="3" resultid="1840" />
                    <RANKING order="4" place="4" resultid="1366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1273" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1274" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1275" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1276" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1327" />
                    <RANKING order="2" place="2" resultid="1952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2086" daytime="17:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2087" daytime="17:44" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1278" daytime="17:48" gender="M" number="44" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1279" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1686" />
                    <RANKING order="2" place="2" resultid="1703" />
                    <RANKING order="3" place="3" resultid="1782" />
                    <RANKING order="4" place="4" resultid="1533" />
                    <RANKING order="5" place="5" resultid="1544" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1512" />
                    <RANKING order="2" place="-1" resultid="1488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1282" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1941" />
                    <RANKING order="2" place="2" resultid="1761" />
                    <RANKING order="3" place="3" resultid="1469" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1283" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1284" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1458" />
                    <RANKING order="2" place="2" resultid="1619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1452" />
                    <RANKING order="2" place="-1" resultid="1334" />
                    <RANKING order="3" place="-1" resultid="1613" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2088" daytime="17:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2089" daytime="17:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2090" daytime="17:54" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1286" daytime="17:56" gender="F" number="45" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1287" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1288" daytime="17:56" gender="M" number="46" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1289" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1567" />
                    <RANKING order="2" place="2" resultid="1424" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2091" daytime="17:56" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1290" daytime="18:00" gender="F" number="47" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1291" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1408" />
                    <RANKING order="2" place="2" resultid="1563" />
                    <RANKING order="3" place="3" resultid="1579" />
                    <RANKING order="4" place="4" resultid="1930" />
                    <RANKING order="5" place="-1" resultid="1596" />
                    <RANKING order="6" place="-1" resultid="1787" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1824" />
                    <RANKING order="2" place="2" resultid="1493" />
                    <RANKING order="3" place="3" resultid="1776" />
                    <RANKING order="4" place="4" resultid="1738" />
                    <RANKING order="5" place="5" resultid="1866" />
                    <RANKING order="6" place="6" resultid="1523" />
                    <RANKING order="7" place="7" resultid="1792" />
                    <RANKING order="8" place="8" resultid="1432" />
                    <RANKING order="9" place="9" resultid="1926" />
                    <RANKING order="10" place="10" resultid="1898" />
                    <RANKING order="11" place="11" resultid="1420" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2092" daytime="18:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2093" daytime="18:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2094" daytime="18:04" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1293" daytime="18:06" gender="M" number="48" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1294" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1851" />
                    <RANKING order="2" place="2" resultid="1412" />
                    <RANKING order="3" place="3" resultid="1882" />
                    <RANKING order="4" place="4" resultid="1902" />
                    <RANKING order="5" place="5" resultid="1934" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1295" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1743" />
                    <RANKING order="2" place="2" resultid="1392" />
                    <RANKING order="3" place="3" resultid="1846" />
                    <RANKING order="4" place="4" resultid="1576" />
                    <RANKING order="5" place="5" resultid="1856" />
                    <RANKING order="6" place="6" resultid="1908" />
                    <RANKING order="7" place="7" resultid="1583" />
                    <RANKING order="8" place="8" resultid="1890" />
                    <RANKING order="9" place="9" resultid="1894" />
                    <RANKING order="10" place="10" resultid="1912" />
                    <RANKING order="11" place="-1" resultid="1428" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2095" daytime="18:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2096" daytime="18:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2097" daytime="18:10" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1296" daytime="18:12" gender="F" number="49" order="26" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1297" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1602" />
                    <RANKING order="2" place="2" resultid="1376" />
                    <RANKING order="3" place="3" resultid="1592" />
                    <RANKING order="4" place="4" resultid="1388" />
                    <RANKING order="5" place="5" resultid="1861" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1298" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1483" />
                    <RANKING order="2" place="2" resultid="1571" />
                    <RANKING order="3" place="3" resultid="1797" />
                    <RANKING order="4" place="4" resultid="1877" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2098" daytime="18:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2099" daytime="18:14" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1299" daytime="18:16" gender="M" number="50" order="27" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1300" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1498" />
                    <RANKING order="2" place="2" resultid="1771" />
                    <RANKING order="3" place="3" resultid="1400" />
                    <RANKING order="4" place="4" resultid="1558" />
                    <RANKING order="5" place="5" resultid="1384" />
                    <RANKING order="6" place="6" resultid="1886" />
                    <RANKING order="7" place="-1" resultid="1518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1301" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1503" />
                    <RANKING order="2" place="2" resultid="1766" />
                    <RANKING order="3" place="3" resultid="1691" />
                    <RANKING order="4" place="4" resultid="1528" />
                    <RANKING order="5" place="5" resultid="1829" />
                    <RANKING order="6" place="6" resultid="1587" />
                    <RANKING order="7" place="7" resultid="1439" />
                    <RANKING order="8" place="8" resultid="1813" />
                    <RANKING order="9" place="9" resultid="1435" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2100" daytime="18:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2101" daytime="18:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2102" daytime="18:20" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1302" daytime="18:22" gender="F" number="51" order="28" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1303" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1983" />
                    <RANKING order="2" place="2" resultid="1709" />
                    <RANKING order="3" place="3" resultid="1538" />
                    <RANKING order="4" place="4" resultid="1359" />
                    <RANKING order="5" place="5" resultid="1341" />
                    <RANKING order="6" place="6" resultid="1995" />
                    <RANKING order="7" place="7" resultid="1554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1304" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1508" />
                    <RANKING order="2" place="2" resultid="1650" />
                    <RANKING order="3" place="3" resultid="1841" />
                    <RANKING order="4" place="4" resultid="1323" />
                    <RANKING order="5" place="5" resultid="1367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1305" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1363" />
                    <RANKING order="2" place="2" resultid="1465" />
                    <RANKING order="3" place="-1" resultid="1656" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1306" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1307" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1308" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1309" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1947" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2103" daytime="18:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2104" daytime="18:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2105" daytime="18:26" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1310" daytime="18:28" gender="M" number="52" order="29" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1311" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1680" />
                    <RANKING order="2" place="2" resultid="1549" />
                    <RANKING order="3" place="3" resultid="1380" />
                    <RANKING order="4" place="4" resultid="1404" />
                    <RANKING order="5" place="5" resultid="1396" />
                    <RANKING order="6" place="6" resultid="1416" />
                    <RANKING order="7" place="7" resultid="2001" />
                    <RANKING order="8" place="8" resultid="1917" />
                    <RANKING order="9" place="-1" resultid="1989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1312" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1513" />
                    <RANKING order="2" place="2" resultid="1662" />
                    <RANKING order="3" place="3" resultid="1755" />
                    <RANKING order="4" place="4" resultid="1668" />
                    <RANKING order="5" place="5" resultid="1872" />
                    <RANKING order="6" place="6" resultid="1922" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1313" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1727" />
                    <RANKING order="2" place="2" resultid="1607" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1314" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1443" />
                    <RANKING order="2" place="2" resultid="1348" />
                    <RANKING order="3" place="3" resultid="1733" />
                    <RANKING order="4" place="4" resultid="1474" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1315" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1352" />
                    <RANKING order="2" place="2" resultid="1462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1316" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1447" />
                    <RANKING order="2" place="2" resultid="1959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1317" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1337" />
                    <RANKING order="2" place="2" resultid="1330" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2106" daytime="18:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2107" daytime="18:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2108" daytime="18:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2109" daytime="18:32" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2110" daytime="18:34" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="3501" nation="BRA" region="PR" clubid="1319" swrid="93752" name="Ortega &amp; De Souza Jesus" shortname="Aquafoz">
          <ATHLETES>
            <ATHLETE firstname="Mateus" lastname="Wirtti" birthdate="2011-01-14" gender="M" nation="BRA" license="383854" swrid="4917570" athleteid="1377" externalid="383854">
              <RESULTS>
                <RESULT eventid="1096" points="288" swimtime="00:01:07.89" resultid="1378" heatid="2019" lane="1" entrytime="00:01:09.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="217" swimtime="00:00:36.77" resultid="1379" heatid="2037" lane="1" entrytime="00:00:39.06" entrycourse="SCM" />
                <RESULT eventid="1310" points="294" swimtime="00:00:30.29" resultid="1380" heatid="2108" lane="2" entrytime="00:00:30.13" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Rorato" birthdate="2013-04-18" gender="F" nation="BRA" license="383851" swrid="5596936" athleteid="1372" externalid="383851">
              <RESULTS>
                <RESULT eventid="1104" points="221" swimtime="00:03:02.19" resultid="1373" heatid="2023" lane="4" entrytime="00:03:09.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.44" />
                    <SPLIT distance="100" swimtime="00:01:26.61" />
                    <SPLIT distance="150" swimtime="00:02:14.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="205" swimtime="00:00:42.82" resultid="1374" heatid="2039" lane="3" entrytime="00:00:43.65" entrycourse="SCM" />
                <RESULT eventid="1264" points="197" swimtime="00:01:37.06" resultid="1375" heatid="2084" lane="2" entrytime="00:01:41.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="246" swimtime="00:00:36.56" resultid="1376" heatid="2099" lane="2" entrytime="00:00:37.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauan" lastname="Matheus Cunha" birthdate="2011-01-31" gender="M" nation="BRA" license="392834" swrid="5641770" athleteid="1393" externalid="392834">
              <RESULTS>
                <RESULT eventid="1096" points="229" swimtime="00:01:13.19" resultid="1394" heatid="2018" lane="5" entrytime="00:01:20.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="205" swimtime="00:00:36.83" resultid="1395" heatid="2080" lane="1" />
                <RESULT eventid="1310" points="240" swimtime="00:00:32.42" resultid="1396" heatid="2108" lane="6" entrytime="00:00:34.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Benicio Martins" birthdate="2013-01-20" gender="M" nation="BRA" license="392831" swrid="5641752" athleteid="1381" externalid="392831">
              <RESULTS>
                <RESULT eventid="1151" points="98" swimtime="00:00:47.83" resultid="1382" heatid="2042" lane="1" entrytime="00:00:50.53" entrycourse="SCM" />
                <RESULT eventid="1267" points="74" swimtime="00:01:57.21" resultid="1383" heatid="2085" lane="2" entrytime="00:01:57.05" entrycourse="SCM" />
                <RESULT eventid="1299" points="90" swimtime="00:00:44.94" resultid="1384" heatid="2101" lane="6" entrytime="00:00:44.22" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Mehl Sarabia" birthdate="2013-03-27" gender="M" nation="BRA" license="392835" swrid="5641771" athleteid="1397" externalid="392835">
              <RESULTS>
                <RESULT eventid="1079" points="104" swimtime="00:01:57.45" resultid="1398" heatid="2007" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="69" swimtime="00:00:53.77" resultid="1399" heatid="2041" lane="2" entrytime="00:00:55.01" entrycourse="SCM" />
                <RESULT eventid="1299" points="108" swimtime="00:00:42.27" resultid="1400" heatid="2101" lane="1" entrytime="00:00:43.07" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="De Albuquerque" birthdate="2014-11-19" gender="F" nation="BRA" license="406648" swrid="4823632" athleteid="1417" externalid="406648">
              <RESULTS>
                <RESULT eventid="1082" points="64" swimtime="00:01:10.75" resultid="1418" heatid="2009" lane="2" entrytime="00:01:23.17" entrycourse="SCM" />
                <RESULT eventid="1154" points="52" swimtime="00:01:07.37" resultid="1419" heatid="2044" lane="6" entrytime="00:01:19.41" entrycourse="SCM" />
                <RESULT eventid="1290" points="61" swimtime="00:00:57.97" resultid="1420" heatid="2093" lane="6" entrytime="00:01:02.43" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julio" lastname="Heck" birthdate="1998-02-15" gender="M" nation="BRA" license="185880" swrid="5596906" athleteid="1335" externalid="185880">
              <RESULTS>
                <RESULT eventid="1096" points="606" swimtime="00:00:52.98" resultid="1336" heatid="2022" lane="3" entrytime="00:00:52.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="584" swimtime="00:00:24.11" resultid="1337" heatid="2110" lane="3" entrytime="00:00:23.75" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gino" lastname="Benicio Ciallella" birthdate="2012-05-21" gender="M" nation="ARG" license="406735" swrid="4492694" athleteid="1433" externalid="406735">
              <RESULTS>
                <RESULT eventid="1151" points="53" swimtime="00:00:58.63" resultid="1434" heatid="2041" lane="5" />
                <RESULT eventid="1299" points="61" swimtime="00:00:51.14" resultid="1435" heatid="2100" lane="4" entrytime="00:01:01.83" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ian" lastname="Peroni Ottomar" birthdate="2016-07-15" gender="M" nation="BRA" license="406653" swrid="5258754" athleteid="1421" externalid="406653">
              <RESULTS>
                <RESULT eventid="1226" points="69" swimtime="00:00:25.03" resultid="1422" heatid="2071" lane="3" entrytime="00:00:27.53" entrycourse="SCM" />
                <RESULT eventid="1262" points="45" swimtime="00:00:32.07" resultid="1423" heatid="2082" lane="3" />
                <RESULT eventid="1288" points="59" swimtime="00:00:23.31" resultid="1424" heatid="2091" lane="3" entrytime="00:00:29.22" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Franco" birthdate="2010-06-09" gender="F" nation="BRA" license="383849" swrid="5596896" athleteid="1320" externalid="383849">
              <RESULTS>
                <RESULT eventid="1088" points="380" swimtime="00:01:09.34" resultid="1321" heatid="2014" lane="3" entrytime="00:01:11.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="336" swimtime="00:05:32.59" resultid="1322" heatid="2059" lane="2" entrytime="00:05:23.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:18.45" />
                    <SPLIT distance="150" swimtime="00:02:01.19" />
                    <SPLIT distance="200" swimtime="00:02:44.23" />
                    <SPLIT distance="250" swimtime="00:03:27.36" />
                    <SPLIT distance="300" swimtime="00:04:09.75" />
                    <SPLIT distance="350" swimtime="00:04:52.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="357" swimtime="00:00:32.32" resultid="1323" heatid="2104" lane="4" entrytime="00:00:32.84" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="De Souza Tulio" birthdate="2006-06-23" gender="F" nation="BRA" license="342344" swrid="5030980" athleteid="1324" externalid="342344">
              <RESULTS>
                <RESULT eventid="1088" points="568" swimtime="00:01:00.65" resultid="1325" heatid="2016" lane="3" entrytime="00:00:58.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="520" swimtime="00:00:31.39" resultid="1326" heatid="2034" lane="3" entrytime="00:00:30.64" entrycourse="SCM" />
                <RESULT eventid="1270" points="498" swimtime="00:01:09.21" resultid="1327" heatid="2087" lane="3" entrytime="00:01:05.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Mussi" birthdate="2006-12-31" gender="M" nation="BRA" license="370567" swrid="5596917" athleteid="1353" externalid="370567">
              <RESULTS>
                <RESULT eventid="1184" points="467" swimtime="00:00:32.14" resultid="1354" heatid="2056" lane="3" entrytime="00:00:32.66" entrycourse="SCM" />
                <RESULT eventid="1236" points="443" swimtime="00:01:12.47" resultid="1355" heatid="2075" lane="5" entrytime="00:01:15.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Victoria Portela" birthdate="2009-12-04" gender="F" nation="BRA" license="383047" swrid="5596945" athleteid="1360" externalid="383047">
              <RESULTS>
                <RESULT eventid="1088" points="461" swimtime="00:01:05.03" resultid="1361" heatid="2016" lane="1" entrytime="00:01:06.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="298" swimtime="00:00:37.77" resultid="1362" heatid="2033" lane="1" />
                <RESULT eventid="1302" points="477" swimtime="00:00:29.33" resultid="1363" heatid="2105" lane="3" entrytime="00:00:30.06" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Pires" birthdate="2011-04-09" gender="F" nation="BRA" license="383853" swrid="5596927" athleteid="1338" externalid="383853">
              <RESULTS>
                <RESULT eventid="1132" status="DSQ" swimtime="00:00:44.64" resultid="1339" heatid="2033" lane="2" entrytime="00:00:45.69" entrycourse="SCM" />
                <RESULT eventid="1176" points="208" swimtime="00:00:47.87" resultid="1340" heatid="2053" lane="1" entrytime="00:00:49.08" entrycourse="SCM" />
                <RESULT eventid="1302" points="225" swimtime="00:00:37.65" resultid="1341" heatid="2104" lane="6" entrytime="00:00:36.93" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Varela" birthdate="2010-05-20" gender="F" nation="BRA" license="365503" swrid="5596942" athleteid="1364" externalid="365503">
              <RESULTS>
                <RESULT eventid="1132" points="173" swimtime="00:00:45.24" resultid="1365" heatid="2034" lane="6" entrytime="00:00:41.25" entrycourse="SCM" />
                <RESULT eventid="1270" points="167" swimtime="00:01:39.55" resultid="1366" heatid="2086" lane="2" entrytime="00:01:27.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="186" swimtime="00:00:40.14" resultid="1367" heatid="2104" lane="2" entrytime="00:00:34.77" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Helena Sousa" birthdate="2013-03-20" gender="F" nation="BRA" license="392832" swrid="5641765" athleteid="1385" externalid="392832">
              <RESULTS>
                <RESULT eventid="1148" points="181" swimtime="00:00:44.62" resultid="1386" heatid="2039" lane="2" entrytime="00:00:48.13" entrycourse="SCM" />
                <RESULT eventid="1264" points="137" swimtime="00:01:49.46" resultid="1387" heatid="2083" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="190" swimtime="00:00:39.86" resultid="1388" heatid="2099" lane="1" entrytime="00:00:41.48" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Geórgia" lastname="Adeli Jesus" birthdate="2008-03-27" gender="F" nation="BRA" license="312649" swrid="5596864" athleteid="1342" externalid="312649">
              <RESULTS>
                <RESULT eventid="1116" points="357" swimtime="00:21:19.63" resultid="1343" heatid="2030" lane="4" entrytime="00:21:25.63" entrycourse="SCM" />
                <RESULT eventid="1192" points="409" swimtime="00:05:11.47" resultid="1344" heatid="2059" lane="4" entrytime="00:05:14.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                    <SPLIT distance="100" swimtime="00:01:11.73" />
                    <SPLIT distance="150" swimtime="00:01:50.81" />
                    <SPLIT distance="200" swimtime="00:02:30.46" />
                    <SPLIT distance="250" swimtime="00:03:10.12" />
                    <SPLIT distance="300" swimtime="00:03:50.70" />
                    <SPLIT distance="350" swimtime="00:04:31.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Gustavo Cunha" birthdate="2011-01-31" gender="M" nation="BRA" license="392836" swrid="5641764" athleteid="1401" externalid="392836">
              <RESULTS>
                <RESULT eventid="1096" points="236" swimtime="00:01:12.50" resultid="1402" heatid="2018" lane="3" entrytime="00:01:13.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="187" swimtime="00:00:43.60" resultid="1403" heatid="2056" lane="6" entrytime="00:00:45.74" entrycourse="SCM" />
                <RESULT eventid="1310" points="248" swimtime="00:00:32.08" resultid="1404" heatid="2108" lane="1" entrytime="00:00:33.62" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karim" lastname="Maruan Jaber" birthdate="2014-11-19" gender="M" nation="BRA" license="392833" swrid="5627304" athleteid="1389" externalid="392833">
              <RESULTS>
                <RESULT eventid="1113" points="140" swimtime="00:01:26.20" resultid="1390" heatid="2029" lane="5" entrytime="00:01:34.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="89" swimtime="00:00:48.60" resultid="1391" heatid="2068" lane="5" entrytime="00:00:56.75" entrycourse="SCM" />
                <RESULT eventid="1293" points="146" swimtime="00:00:38.25" resultid="1392" heatid="2097" lane="5" entrytime="00:00:41.23" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="De Zanchet" birthdate="2015-09-16" gender="M" nation="BRA" license="392838" swrid="5641762" athleteid="1409" externalid="392838">
              <RESULTS>
                <RESULT eventid="1085" points="99" swimtime="00:00:53.91" resultid="1410" heatid="2012" lane="4" entrytime="00:00:52.63" entrycourse="SCM" />
                <RESULT eventid="1113" points="86" swimtime="00:01:41.41" resultid="1411" heatid="2028" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1293" points="112" swimtime="00:00:41.76" resultid="1412" heatid="2096" lane="3" entrytime="00:00:45.10" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emma" lastname="Raquel Nascimento" birthdate="2015-11-06" gender="F" nation="BRA" license="392837" swrid="5641775" athleteid="1405" externalid="392837">
              <RESULTS>
                <RESULT eventid="1082" points="175" swimtime="00:00:50.72" resultid="1406" heatid="2010" lane="4" entrytime="00:00:49.37" entrycourse="SCM" />
                <RESULT eventid="1110" points="139" swimtime="00:01:36.78" resultid="1407" heatid="2026" lane="5" />
                <RESULT eventid="1290" points="170" swimtime="00:00:41.39" resultid="1408" heatid="2094" lane="2" entrytime="00:00:40.35" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vicente" lastname="Duarte Martins" birthdate="2014-12-23" gender="M" nation="BRA" license="406654" swrid="4956741" athleteid="1425" externalid="406654">
              <RESULTS>
                <RESULT eventid="1085" status="DNS" swimtime="00:00:00.00" resultid="1426" heatid="2012" lane="6" entrytime="00:01:31.16" entrycourse="SCM" />
                <RESULT eventid="1157" status="DNS" swimtime="00:00:00.00" resultid="1427" heatid="2046" lane="1" />
                <RESULT eventid="1293" status="DNS" swimtime="00:00:00.00" resultid="1428" heatid="2096" lane="5" entrytime="00:01:04.88" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Dominguez Olivieski" birthdate="2011-04-27" gender="M" nation="BRA" license="405717" swrid="5664737" athleteid="1413" externalid="405717">
              <RESULTS>
                <RESULT eventid="1096" points="197" swimtime="00:01:17.04" resultid="1414" heatid="2018" lane="2" entrytime="00:01:17.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="211" swimtime="00:01:32.80" resultid="1415" heatid="2074" lane="5" entrytime="00:01:40.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="233" swimtime="00:00:32.76" resultid="1416" heatid="2107" lane="3" entrytime="00:00:35.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Mendes Portela" birthdate="2014-03-08" gender="F" nation="BRA" license="406656" swrid="5117156" athleteid="1429" externalid="406656">
              <RESULTS>
                <RESULT eventid="1082" points="87" swimtime="00:01:03.91" resultid="1430" heatid="2009" lane="4" entrytime="00:01:12.22" entrycourse="SCM" />
                <RESULT eventid="1110" points="94" swimtime="00:01:50.27" resultid="1431" heatid="2026" lane="3" />
                <RESULT eventid="1290" points="134" swimtime="00:00:44.76" resultid="1432" heatid="2093" lane="1" entrytime="00:00:53.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paulo" lastname="Antonio Sousa" birthdate="2012-03-17" gender="M" nation="BRA" license="407497" swrid="5721498" athleteid="1436" externalid="407497">
              <RESULTS>
                <RESULT eventid="1079" points="115" swimtime="00:01:53.53" resultid="1437" heatid="2008" lane="5" entrytime="00:01:55.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="101" swimtime="00:00:47.45" resultid="1438" heatid="2040" lane="2" />
                <RESULT eventid="1299" points="135" swimtime="00:00:39.29" resultid="1439" heatid="2101" lane="4" entrytime="00:00:38.23" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Afonso Proteti" birthdate="2002-03-19" gender="M" nation="BRA" license="190464" swrid="5596865" athleteid="1331" externalid="190464">
              <RESULTS>
                <RESULT eventid="1140" points="528" swimtime="00:00:27.35" resultid="1332" heatid="2037" lane="3" entrytime="00:00:26.72" entrycourse="SCM" />
                <RESULT eventid="1252" points="659" swimtime="00:00:24.99" resultid="1333" heatid="2081" lane="3" entrytime="00:00:25.45" entrycourse="SCM" />
                <RESULT eventid="1278" status="DSQ" swimtime="00:00:59.85" resultid="1334" heatid="2090" lane="3" entrytime="00:00:57.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Gabriel Serighelli" birthdate="1999-03-12" gender="M" nation="BRA" license="121253" swrid="5596899" athleteid="1328" externalid="121253">
              <RESULTS>
                <RESULT eventid="1096" points="536" swimtime="00:00:55.19" resultid="1329" heatid="2022" lane="4" entrytime="00:00:55.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="559" swimtime="00:00:24.46" resultid="1330" heatid="2110" lane="4" entrytime="00:00:24.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yago" lastname="Simon Pires" birthdate="2008-10-29" gender="M" nation="BRA" license="328942" swrid="5596939" athleteid="1345" externalid="328942">
              <RESULTS>
                <RESULT eventid="1096" points="451" swimtime="00:00:58.47" resultid="1346" heatid="2021" lane="2" entrytime="00:00:59.36" entrycourse="SCM" />
                <RESULT eventid="1184" points="405" swimtime="00:00:33.70" resultid="1347" heatid="2056" lane="2" entrytime="00:00:33.95" entrycourse="SCM" />
                <RESULT eventid="1310" points="424" swimtime="00:00:26.83" resultid="1348" heatid="2109" lane="3" entrytime="00:00:26.58" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Marques Lima" birthdate="2010-04-30" gender="F" nation="BRA" license="383051" swrid="5596913" athleteid="1368" externalid="383051">
              <RESULTS>
                <RESULT eventid="1160" points="279" swimtime="00:01:22.66" resultid="1369" heatid="2048" lane="1" entrytime="00:01:26.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1244" points="341" swimtime="00:00:34.88" resultid="1370" heatid="2078" lane="6" entrytime="00:00:37.40" entrycourse="SCM" />
                <RESULT eventid="1270" points="305" swimtime="00:01:21.53" resultid="1371" heatid="2086" lane="3" entrytime="00:01:19.83" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Otremba Rouver" birthdate="2007-04-25" gender="M" nation="BRA" license="342152" swrid="5596919" athleteid="1349" externalid="342152">
              <RESULTS>
                <RESULT eventid="1096" points="433" swimtime="00:00:59.24" resultid="1350" heatid="2022" lane="5" entrytime="00:00:56.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="447" swimtime="00:00:28.44" resultid="1351" heatid="2081" lane="4" entrytime="00:00:27.44" entrycourse="SCM" />
                <RESULT eventid="1310" points="403" swimtime="00:00:27.28" resultid="1352" heatid="2110" lane="1" entrytime="00:00:25.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Maguet" birthdate="2011-07-01" gender="F" nation="BRA" license="370568" swrid="5596911" athleteid="1356" externalid="370568">
              <RESULTS>
                <RESULT eventid="1088" points="275" swimtime="00:01:17.26" resultid="1357" heatid="2014" lane="1" entrytime="00:01:18.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="218" swimtime="00:00:41.92" resultid="1358" heatid="2033" lane="3" entrytime="00:00:43.15" entrycourse="SCM" />
                <RESULT eventid="1302" points="270" swimtime="00:00:35.46" resultid="1359" heatid="2104" lane="1" entrytime="00:00:36.04" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18151" nation="BRA" region="PR" clubid="1597" swrid="95180" name="Clube Uniao Recreativo Palmense" shortname="Clube União">
          <ATHLETES>
            <ATHLETE firstname="Luiza" lastname="Langaro Spaniol" birthdate="2013-06-18" gender="F" nation="BRA" license="406600" swrid="5074027" athleteid="1598" externalid="406600">
              <RESULTS>
                <RESULT eventid="1076" points="333" swimtime="00:01:29.90" resultid="1599" heatid="2006" lane="3" entrytime="00:01:30.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="306" swimtime="00:00:37.45" resultid="1600" heatid="2038" lane="4" />
                <RESULT eventid="1264" points="341" swimtime="00:01:20.86" resultid="1601" heatid="2083" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="364" swimtime="00:00:32.09" resultid="1602" heatid="2099" lane="3" entrytime="00:00:32.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lohan" lastname="Henrique Oliveira" birthdate="2009-03-13" gender="M" nation="BRA" license="410110" athleteid="1603" externalid="410110">
              <RESULTS>
                <RESULT eventid="1184" points="236" swimtime="00:00:40.35" resultid="1604" heatid="2055" lane="5" />
                <RESULT eventid="1200" points="180" swimtime="00:06:15.66" resultid="1605" heatid="2061" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:17.28" />
                    <SPLIT distance="150" swimtime="00:02:01.38" />
                    <SPLIT distance="200" swimtime="00:02:50.43" />
                    <SPLIT distance="250" swimtime="00:03:39.64" />
                    <SPLIT distance="300" swimtime="00:04:31.86" />
                    <SPLIT distance="350" swimtime="00:05:26.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="185" swimtime="00:00:38.15" resultid="1606" heatid="2080" lane="4" />
                <RESULT eventid="1310" points="241" swimtime="00:00:32.39" resultid="1607" heatid="2106" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="36" nation="BRA" region="PR" clubid="1608" swrid="93753" name="Associação Atlética Comercial" shortname="Comercial Cascavel">
          <ATHLETES>
            <ATHLETE firstname="João" lastname="Pedro Serafini" birthdate="2012-05-15" gender="M" nation="BRA" license="365488" swrid="5596924" athleteid="1762" externalid="365488">
              <RESULTS>
                <RESULT eventid="1107" points="213" swimtime="00:02:46.25" resultid="1763" heatid="2025" lane="4" entrytime="00:02:47.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:01:21.28" />
                    <SPLIT distance="150" swimtime="00:02:05.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="143" swimtime="00:00:42.24" resultid="1764" heatid="2042" lane="2" entrytime="00:00:44.34" entrycourse="SCM" />
                <RESULT eventid="1221" points="131" swimtime="00:01:34.07" resultid="1765" heatid="2070" lane="2" entrytime="00:01:38.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="204" swimtime="00:00:34.21" resultid="1766" heatid="2101" lane="3" entrytime="00:00:36.93" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luann" lastname="Miguel Mazur" birthdate="2007-01-10" gender="M" nation="BRA" license="365682" swrid="5596915" athleteid="1669" externalid="365682">
              <RESULTS>
                <RESULT eventid="1068" points="473" swimtime="00:02:20.63" resultid="1670" heatid="2005" lane="4" entrytime="00:02:21.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="100" swimtime="00:01:07.80" />
                    <SPLIT distance="150" swimtime="00:01:47.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="285" swimtime="00:00:33.59" resultid="1671" heatid="2036" lane="2" />
                <RESULT eventid="1184" points="414" swimtime="00:00:33.46" resultid="1672" heatid="2054" lane="4" />
                <RESULT eventid="1200" points="493" swimtime="00:04:28.65" resultid="1673" heatid="2063" lane="1" entrytime="00:04:36.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                    <SPLIT distance="100" swimtime="00:01:05.36" />
                    <SPLIT distance="150" swimtime="00:01:39.80" />
                    <SPLIT distance="200" swimtime="00:02:14.06" />
                    <SPLIT distance="250" swimtime="00:02:48.95" />
                    <SPLIT distance="300" swimtime="00:03:24.11" />
                    <SPLIT distance="350" swimtime="00:03:55.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="472" swimtime="00:01:10.95" resultid="1674" heatid="2075" lane="4" entrytime="00:01:11.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raul" lastname="Bonamigo" birthdate="2010-12-01" gender="M" nation="BRA" license="344397" swrid="5588559" athleteid="1750" externalid="344397">
              <RESULTS>
                <RESULT eventid="1068" points="396" swimtime="00:02:29.24" resultid="1751" heatid="2005" lane="1" entrytime="00:02:28.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                    <SPLIT distance="100" swimtime="00:01:09.47" />
                    <SPLIT distance="150" swimtime="00:01:55.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="380" swimtime="00:01:01.90" resultid="1752" heatid="2020" lane="2" entrytime="00:01:01.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="335" swimtime="00:01:08.77" resultid="1753" heatid="2050" lane="5" entrytime="00:01:15.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="448" swimtime="00:04:37.25" resultid="1754" heatid="2063" lane="5" entrytime="00:04:35.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                    <SPLIT distance="100" swimtime="00:01:06.21" />
                    <SPLIT distance="150" swimtime="00:01:41.03" />
                    <SPLIT distance="200" swimtime="00:02:15.94" />
                    <SPLIT distance="250" swimtime="00:02:51.11" />
                    <SPLIT distance="300" swimtime="00:03:26.91" />
                    <SPLIT distance="350" swimtime="00:04:02.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="344" swimtime="00:00:28.77" resultid="1755" heatid="2108" lane="4" entrytime="00:00:30.09" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Mariotti De Castro" birthdate="2008-06-27" gender="M" nation="BRA" license="329200" swrid="5596912" athleteid="1630" externalid="329200">
              <RESULTS>
                <RESULT eventid="1200" points="599" swimtime="00:04:11.69" resultid="1631" heatid="2064" lane="3" entrytime="00:04:03.58" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Danilo" lastname="Rodrigues" birthdate="2011-05-23" gender="M" nation="BRA" license="370763" swrid="5596934" athleteid="1716" externalid="370763">
              <RESULTS>
                <RESULT eventid="1068" points="336" swimtime="00:02:37.59" resultid="1717" heatid="2004" lane="1" entrytime="00:02:47.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                    <SPLIT distance="100" swimtime="00:01:16.51" />
                    <SPLIT distance="150" swimtime="00:02:02.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="401" swimtime="00:19:08.39" resultid="1718" heatid="2031" lane="5" entrytime="00:19:47.68" entrycourse="SCM" />
                <RESULT eventid="1168" points="265" swimtime="00:01:14.38" resultid="1719" heatid="2050" lane="2" entrytime="00:01:14.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="385" swimtime="00:04:51.61" resultid="1720" heatid="2061" lane="3" entrytime="00:05:17.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:09.48" />
                    <SPLIT distance="150" swimtime="00:01:46.74" />
                    <SPLIT distance="200" swimtime="00:02:23.69" />
                    <SPLIT distance="250" swimtime="00:03:01.10" />
                    <SPLIT distance="300" swimtime="00:03:38.57" />
                    <SPLIT distance="350" swimtime="00:04:16.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="300" swimtime="00:01:22.52" resultid="1721" heatid="2074" lane="4" entrytime="00:01:28.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Queiroz Da Costa" birthdate="2014-05-30" gender="F" nation="BRA" license="406698" swrid="5335148" athleteid="1862" externalid="406698">
              <RESULTS>
                <RESULT eventid="1082" points="177" swimtime="00:00:50.46" resultid="1863" heatid="2009" lane="3" entrytime="00:01:03.99" entrycourse="SCM" />
                <RESULT eventid="1110" points="160" swimtime="00:01:32.51" resultid="1864" heatid="2027" lane="2" entrytime="00:01:29.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="102" swimtime="00:00:52.05" resultid="1865" heatid="2066" lane="5" entrytime="00:00:52.29" entrycourse="SCM" />
                <RESULT eventid="1290" points="183" swimtime="00:00:40.36" resultid="1866" heatid="2094" lane="3" entrytime="00:00:39.65" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Souza Garute Da Silva" birthdate="2009-01-07" gender="F" nation="BRA" license="329307" swrid="5596940" athleteid="1632" externalid="329307">
              <RESULTS>
                <RESULT eventid="1088" points="453" swimtime="00:01:05.40" resultid="1633" heatid="2013" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="391" swimtime="00:00:34.53" resultid="1634" heatid="2032" lane="3" />
                <RESULT eventid="1192" points="437" swimtime="00:05:04.77" resultid="1635" heatid="2060" lane="3" entrytime="00:04:47.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                    <SPLIT distance="100" swimtime="00:01:10.94" />
                    <SPLIT distance="150" swimtime="00:01:48.94" />
                    <SPLIT distance="200" swimtime="00:02:27.76" />
                    <SPLIT distance="250" swimtime="00:03:06.77" />
                    <SPLIT distance="300" swimtime="00:03:46.61" />
                    <SPLIT distance="350" swimtime="00:04:26.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="396" swimtime="00:01:14.70" resultid="1636" heatid="2087" lane="2" entrytime="00:01:13.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Kupicki" birthdate="2004-03-02" gender="F" nation="BRA" license="311897" swrid="5624094" athleteid="1620" externalid="311897">
              <RESULTS>
                <RESULT eventid="1088" points="346" swimtime="00:01:11.55" resultid="1621" heatid="2016" lane="2" entrytime="00:01:06.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="278" swimtime="00:00:38.66" resultid="1622" heatid="2032" lane="2" />
                <RESULT eventid="1244" points="336" swimtime="00:00:35.05" resultid="1623" heatid="2076" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benicio" lastname="Hermisdorff Bruning" birthdate="2015-06-22" gender="M" nation="BRA" license="414000" athleteid="1878" externalid="414000">
              <RESULTS>
                <RESULT eventid="1085" points="74" swimtime="00:00:59.40" resultid="1879" heatid="2011" lane="2" />
                <RESULT eventid="1113" points="93" swimtime="00:01:38.86" resultid="1880" heatid="2028" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="63" swimtime="00:00:54.57" resultid="1881" heatid="2067" lane="2" />
                <RESULT eventid="1293" points="100" swimtime="00:00:43.35" resultid="1882" heatid="2095" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Alves Serafini" birthdate="2008-04-15" gender="M" nation="BRA" license="351644" swrid="5596867" athleteid="1756" externalid="351644">
              <RESULTS>
                <RESULT eventid="1068" points="416" swimtime="00:02:26.76" resultid="1757" heatid="2005" lane="2" entrytime="00:02:25.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                    <SPLIT distance="100" swimtime="00:01:07.64" />
                    <SPLIT distance="150" swimtime="00:01:53.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="454" swimtime="00:00:58.31" resultid="1758" heatid="2022" lane="6" entrytime="00:00:57.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="470" swimtime="00:01:01.44" resultid="1759" heatid="2051" lane="4" entrytime="00:01:01.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="504" swimtime="00:04:26.69" resultid="1760" heatid="2063" lane="3" entrytime="00:04:29.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                    <SPLIT distance="100" swimtime="00:01:03.50" />
                    <SPLIT distance="150" swimtime="00:01:37.04" />
                    <SPLIT distance="200" swimtime="00:02:10.79" />
                    <SPLIT distance="250" swimtime="00:02:44.30" />
                    <SPLIT distance="300" swimtime="00:03:18.72" />
                    <SPLIT distance="350" swimtime="00:03:52.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="344" swimtime="00:01:08.94" resultid="1761" heatid="2088" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Breno" lastname="Zanella Janke" birthdate="2011-04-26" gender="M" nation="BRA" license="365697" swrid="5588970" athleteid="1698" externalid="365697">
              <RESULTS>
                <RESULT eventid="1068" points="378" swimtime="00:02:31.56" resultid="1699" heatid="2005" lane="5" entrytime="00:02:28.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.31" />
                    <SPLIT distance="100" swimtime="00:01:12.51" />
                    <SPLIT distance="150" swimtime="00:01:55.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="298" swimtime="00:01:11.52" resultid="1700" heatid="2051" lane="5" entrytime="00:01:09.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="423" swimtime="00:04:42.73" resultid="1701" heatid="2062" lane="3" entrytime="00:04:42.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="100" swimtime="00:01:07.78" />
                    <SPLIT distance="150" swimtime="00:01:43.94" />
                    <SPLIT distance="200" swimtime="00:02:21.09" />
                    <SPLIT distance="250" swimtime="00:02:55.87" />
                    <SPLIT distance="300" swimtime="00:03:31.45" />
                    <SPLIT distance="350" swimtime="00:04:06.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="341" swimtime="00:01:19.12" resultid="1702" heatid="2074" lane="3" entrytime="00:01:18.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="294" swimtime="00:01:12.68" resultid="1703" heatid="2089" lane="1" entrytime="00:01:18.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maite" lastname="Poglia Brenner" birthdate="2014-05-13" gender="F" nation="BRA" license="414004" athleteid="1895" externalid="414004">
              <RESULTS>
                <RESULT eventid="1082" points="67" swimtime="00:01:09.63" resultid="1896" heatid="2009" lane="1" />
                <RESULT eventid="1154" points="59" swimtime="00:01:04.50" resultid="1897" heatid="2043" lane="4" />
                <RESULT eventid="1290" points="77" swimtime="00:00:53.68" resultid="1898" heatid="2092" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marianna" lastname="Galvao Oliveira" birthdate="2014-03-18" gender="F" nation="BRA" license="390835" swrid="5596902" athleteid="1772" externalid="390835">
              <RESULTS>
                <RESULT eventid="1082" points="207" swimtime="00:00:47.92" resultid="1773" heatid="2010" lane="3" entrytime="00:00:47.11" entrycourse="SCM" />
                <RESULT eventid="1110" points="181" swimtime="00:01:28.68" resultid="1774" heatid="2027" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="142" swimtime="00:00:46.64" resultid="1775" heatid="2066" lane="4" entrytime="00:00:50.00" entrycourse="SCM" />
                <RESULT eventid="1290" points="223" swimtime="00:00:37.78" resultid="1776" heatid="2094" lane="4" entrytime="00:00:39.95" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Bortoli Da Silva" birthdate="2010-09-30" gender="M" nation="BRA" license="365500" athleteid="1867" externalid="365500">
              <RESULTS>
                <RESULT eventid="1096" points="277" swimtime="00:01:08.74" resultid="1868" heatid="2017" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="208" swimtime="00:01:20.59" resultid="1869" heatid="2049" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="290" swimtime="00:05:20.60" resultid="1870" heatid="2061" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:01:14.35" />
                    <SPLIT distance="150" swimtime="00:01:55.14" />
                    <SPLIT distance="200" swimtime="00:02:35.89" />
                    <SPLIT distance="250" swimtime="00:03:18.49" />
                    <SPLIT distance="300" swimtime="00:04:00.48" />
                    <SPLIT distance="350" swimtime="00:04:41.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="219" swimtime="00:00:36.03" resultid="1871" heatid="2079" lane="3" />
                <RESULT eventid="1310" points="236" swimtime="00:00:32.61" resultid="1872" heatid="2107" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Gaio" birthdate="2014-08-27" gender="F" nation="BRA" license="390841" swrid="5596900" athleteid="1788" externalid="390841">
              <RESULTS>
                <RESULT eventid="1082" points="150" swimtime="00:00:53.31" resultid="1789" heatid="2010" lane="5" entrytime="00:00:52.96" entrycourse="SCM" />
                <RESULT eventid="1110" points="130" swimtime="00:01:39.05" resultid="1790" heatid="2027" lane="1" entrytime="00:01:49.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="92" swimtime="00:00:53.91" resultid="1791" heatid="2066" lane="1" entrytime="00:00:52.73" entrycourse="SCM" />
                <RESULT eventid="1290" points="140" swimtime="00:00:44.12" resultid="1792" heatid="2093" lane="3" entrytime="00:00:44.06" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Douglas" lastname="Dos Santos Luz" birthdate="2013-12-10" gender="M" nation="BRA" license="414001" athleteid="1883" externalid="414001">
              <RESULTS>
                <RESULT eventid="1079" points="38" swimtime="00:02:43.94" resultid="1884" heatid="2007" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="45" swimtime="00:01:01.95" resultid="1885" heatid="2040" lane="3" />
                <RESULT eventid="1299" points="36" swimtime="00:01:00.69" resultid="1886" heatid="2100" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jordana" lastname="Rinaldini" birthdate="2004-09-13" gender="F" nation="BRA" license="342426" swrid="5596933" athleteid="1637" externalid="342426">
              <RESULTS>
                <RESULT eventid="1060" points="370" swimtime="00:02:49.71" resultid="1638" heatid="2003" lane="4" entrytime="00:02:50.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="100" swimtime="00:01:18.02" />
                    <SPLIT distance="150" swimtime="00:02:08.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="383" swimtime="00:00:39.06" resultid="1639" heatid="2053" lane="4" entrytime="00:00:39.15" entrycourse="SCM" />
                <RESULT eventid="1228" points="427" swimtime="00:01:22.78" resultid="1640" heatid="2072" lane="4" entrytime="00:01:24.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laisa" lastname="Bernardini" birthdate="2012-06-25" gender="F" nation="BRA" license="390843" swrid="5596872" athleteid="1798" externalid="390843">
              <RESULTS>
                <RESULT eventid="1076" points="219" swimtime="00:01:43.40" resultid="1799" heatid="2006" lane="2" entrytime="00:01:46.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="203" swimtime="00:00:42.91" resultid="1800" heatid="2038" lane="2" />
                <RESULT eventid="1218" points="169" swimtime="00:01:37.76" resultid="1801" heatid="2069" lane="3" entrytime="00:01:45.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="242" swimtime="00:01:30.61" resultid="1802" heatid="2084" lane="4" entrytime="00:01:39.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Michelsen Vidal" birthdate="2015-11-29" gender="M" nation="BRA" license="414005" athleteid="1899" externalid="414005">
              <RESULTS>
                <RESULT eventid="1085" points="66" swimtime="00:01:01.64" resultid="1900" heatid="2011" lane="4" />
                <RESULT eventid="1157" points="72" swimtime="00:00:53.03" resultid="1901" heatid="2046" lane="5" />
                <RESULT eventid="1293" points="95" swimtime="00:00:44.17" resultid="1902" heatid="2095" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia" lastname="Oliveira Faria" birthdate="2013-10-04" gender="F" nation="BRA" license="406697" swrid="5227019" athleteid="1857" externalid="406697">
              <RESULTS>
                <RESULT eventid="1104" points="150" swimtime="00:03:27.19" resultid="1858" heatid="2023" lane="5" entrytime="00:04:09.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.38" />
                    <SPLIT distance="100" swimtime="00:01:37.82" />
                    <SPLIT distance="150" swimtime="00:02:33.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="133" swimtime="00:00:49.35" resultid="1859" heatid="2039" lane="1" entrytime="00:00:59.39" entrycourse="SCM" />
                <RESULT eventid="1264" status="DSQ" swimtime="00:01:50.15" resultid="1860" heatid="2084" lane="5" entrytime="00:02:12.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="182" swimtime="00:00:40.39" resultid="1861" heatid="2098" lane="4" entrytime="00:00:48.76" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Bertelli Weirich" birthdate="2011-03-18" gender="F" nation="BRA" license="369534" swrid="5588552" athleteid="1704" externalid="369534">
              <RESULTS>
                <RESULT eventid="1088" points="404" swimtime="00:01:07.95" resultid="1705" heatid="2015" lane="3" entrytime="00:01:07.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="336" swimtime="00:00:40.77" resultid="1706" heatid="2052" lane="2" />
                <RESULT eventid="1192" points="433" swimtime="00:05:05.72" resultid="1707" heatid="2060" lane="5" entrytime="00:05:01.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                    <SPLIT distance="100" swimtime="00:01:11.70" />
                    <SPLIT distance="150" swimtime="00:01:49.90" />
                    <SPLIT distance="200" swimtime="00:02:28.57" />
                    <SPLIT distance="250" swimtime="00:03:07.70" />
                    <SPLIT distance="300" swimtime="00:03:47.43" />
                    <SPLIT distance="350" swimtime="00:04:26.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1244" points="336" swimtime="00:00:35.05" resultid="1708" heatid="2078" lane="5" entrytime="00:00:35.58" entrycourse="SCM" />
                <RESULT eventid="1302" points="365" swimtime="00:00:32.08" resultid="1709" heatid="2103" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ramirez Vasconcelos" birthdate="2011-04-06" gender="M" nation="BRA" license="392013" swrid="4863662" athleteid="1814" externalid="392013">
              <RESULTS>
                <RESULT eventid="1068" points="305" swimtime="00:02:42.84" resultid="1815" heatid="2004" lane="6" entrytime="00:02:53.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                    <SPLIT distance="100" swimtime="00:01:19.24" />
                    <SPLIT distance="150" swimtime="00:02:05.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="286" swimtime="00:01:08.00" resultid="1816" heatid="2019" lane="2" entrytime="00:01:08.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="283" swimtime="00:00:37.99" resultid="1817" heatid="2056" lane="5" entrytime="00:00:38.91" entrycourse="SCM" />
                <RESULT eventid="1200" points="319" swimtime="00:05:10.32" resultid="1818" heatid="2061" lane="2" entrytime="00:05:24.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                    <SPLIT distance="100" swimtime="00:01:14.08" />
                    <SPLIT distance="150" swimtime="00:01:54.30" />
                    <SPLIT distance="200" swimtime="00:02:34.99" />
                    <SPLIT distance="250" swimtime="00:03:15.14" />
                    <SPLIT distance="300" swimtime="00:03:55.31" />
                    <SPLIT distance="350" swimtime="00:04:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="254" swimtime="00:00:34.32" resultid="1819" heatid="2080" lane="3" entrytime="00:00:38.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Do Prado Martins" birthdate="2008-10-17" gender="F" nation="BRA" license="369419" swrid="5596893" athleteid="1692" externalid="369419">
              <RESULTS>
                <RESULT eventid="1088" points="476" swimtime="00:01:04.33" resultid="1693" heatid="2016" lane="5" entrytime="00:01:06.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="489" swimtime="00:00:36.00" resultid="1694" heatid="2052" lane="5" />
                <RESULT eventid="1192" points="491" swimtime="00:04:53.13" resultid="1695" heatid="2060" lane="4" entrytime="00:04:56.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:09.09" />
                    <SPLIT distance="150" swimtime="00:01:45.81" />
                    <SPLIT distance="200" swimtime="00:02:22.76" />
                    <SPLIT distance="250" swimtime="00:03:00.36" />
                    <SPLIT distance="300" swimtime="00:03:38.44" />
                    <SPLIT distance="350" swimtime="00:04:16.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="485" swimtime="00:01:19.32" resultid="1696" heatid="2072" lane="3" entrytime="00:01:19.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="416" swimtime="00:00:30.71" resultid="1697" heatid="2103" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Bonamigo" birthdate="2013-06-25" gender="M" nation="BRA" license="365484" swrid="5588558" athleteid="1767" externalid="365484">
              <RESULTS>
                <RESULT eventid="1079" points="239" swimtime="00:01:28.99" resultid="1768" heatid="2008" lane="3" entrytime="00:01:28.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="191" swimtime="00:00:38.39" resultid="1769" heatid="2040" lane="4" />
                <RESULT eventid="1267" points="205" swimtime="00:01:23.57" resultid="1770" heatid="2085" lane="3" entrytime="00:01:25.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="236" swimtime="00:00:32.60" resultid="1771" heatid="2102" lane="2" entrytime="00:00:33.62" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Luis Lottermann" birthdate="2014-10-08" gender="M" nation="BRA" license="382237" swrid="5596908" athleteid="1739" externalid="382237">
              <RESULTS>
                <RESULT eventid="1085" points="127" swimtime="00:00:49.53" resultid="1740" heatid="2012" lane="5" entrytime="00:00:53.06" entrycourse="SCM" />
                <RESULT eventid="1113" points="192" swimtime="00:01:17.64" resultid="1741" heatid="2029" lane="3" entrytime="00:01:16.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="152" swimtime="00:00:40.71" resultid="1742" heatid="2068" lane="4" entrytime="00:00:45.02" entrycourse="SCM" />
                <RESULT eventid="1293" points="168" swimtime="00:00:36.51" resultid="1743" heatid="2097" lane="3" entrytime="00:00:35.50" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Gabriel Dalchau" birthdate="2014-08-27" gender="M" nation="BRA" license="402118" swrid="5661346" athleteid="1842" externalid="402118">
              <RESULTS>
                <RESULT eventid="1113" points="140" swimtime="00:01:26.21" resultid="1843" heatid="2029" lane="2" entrytime="00:01:32.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="117" swimtime="00:00:45.20" resultid="1844" heatid="2046" lane="4" entrytime="00:00:47.58" entrycourse="SCM" />
                <RESULT eventid="1215" points="66" swimtime="00:00:53.71" resultid="1845" heatid="2067" lane="3" />
                <RESULT eventid="1293" points="139" swimtime="00:00:38.87" resultid="1846" heatid="2097" lane="6" entrytime="00:00:42.49" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Livia" lastname="De Oliveira" birthdate="2012-02-07" gender="F" nation="BRA" license="413999" athleteid="1873" externalid="413999">
              <RESULTS>
                <RESULT eventid="1076" points="90" swimtime="00:02:18.82" resultid="1874" heatid="2006" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="73" swimtime="00:01:00.32" resultid="1875" heatid="2038" lane="3" />
                <RESULT eventid="1264" points="96" swimtime="00:02:03.04" resultid="1876" heatid="2083" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="101" swimtime="00:00:49.22" resultid="1877" heatid="2098" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Vitoria Gugel" birthdate="2011-12-08" gender="F" nation="BRA" license="365490" swrid="5588960" athleteid="1830" externalid="365490">
              <RESULTS>
                <RESULT eventid="1060" points="337" swimtime="00:02:55.04" resultid="1831" heatid="2003" lane="5" entrytime="00:02:55.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.46" />
                    <SPLIT distance="100" swimtime="00:01:23.13" />
                    <SPLIT distance="150" swimtime="00:02:13.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="340" swimtime="00:01:11.93" resultid="1832" heatid="2014" lane="2" entrytime="00:01:15.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="303" swimtime="00:01:20.44" resultid="1833" heatid="2048" lane="5" entrytime="00:01:24.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="340" swimtime="00:05:31.15" resultid="1834" heatid="2058" lane="4" entrytime="00:05:38.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                    <SPLIT distance="100" swimtime="00:01:17.19" />
                    <SPLIT distance="150" swimtime="00:01:58.24" />
                    <SPLIT distance="200" swimtime="00:02:39.75" />
                    <SPLIT distance="250" swimtime="00:03:20.81" />
                    <SPLIT distance="300" swimtime="00:04:03.68" />
                    <SPLIT distance="350" swimtime="00:04:47.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="301" swimtime="00:01:32.96" resultid="1835" heatid="2072" lane="5" entrytime="00:01:37.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Flavia" lastname="De Metz" birthdate="2011-01-07" gender="F" nation="BRA" license="390846" swrid="5596887" athleteid="1803" externalid="390846">
              <RESULTS>
                <RESULT eventid="1060" points="343" swimtime="00:02:53.95" resultid="1804" heatid="2002" lane="4" entrytime="00:03:03.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:01:22.60" />
                    <SPLIT distance="150" swimtime="00:02:16.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="338" swimtime="00:21:42.84" resultid="1805" heatid="2030" lane="1" />
                <RESULT eventid="1160" points="223" swimtime="00:01:29.05" resultid="1806" heatid="2047" lane="4" entrytime="00:01:37.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="405" swimtime="00:05:12.58" resultid="1807" heatid="2059" lane="5" entrytime="00:05:24.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.69" />
                    <SPLIT distance="100" swimtime="00:01:12.21" />
                    <SPLIT distance="150" swimtime="00:01:50.86" />
                    <SPLIT distance="200" swimtime="00:02:31.18" />
                    <SPLIT distance="250" swimtime="00:03:11.24" />
                    <SPLIT distance="300" swimtime="00:03:51.79" />
                    <SPLIT distance="350" swimtime="00:04:32.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="307" swimtime="00:01:21.30" resultid="1808" heatid="2087" lane="1" entrytime="00:01:19.25" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabelle" lastname="Cordeiro Silva" birthdate="2015-06-14" gender="F" nation="BRA" license="390839" swrid="5596878" athleteid="1783" externalid="390839">
              <RESULTS>
                <RESULT eventid="1082" status="DNS" swimtime="00:00:00.00" resultid="1784" heatid="2010" lane="2" entrytime="00:00:52.45" entrycourse="SCM" />
                <RESULT eventid="1154" status="DNS" swimtime="00:00:00.00" resultid="1785" heatid="2044" lane="5" entrytime="00:00:51.43" entrycourse="SCM" />
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="1786" heatid="2066" lane="6" entrytime="00:00:53.12" entrycourse="SCM" />
                <RESULT eventid="1290" status="DNS" swimtime="00:00:00.00" resultid="1787" heatid="2093" lane="2" entrytime="00:00:45.44" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Tolentino Smarczewski" birthdate="2008-09-01" gender="M" nation="BRA" license="378818" swrid="5596941" athleteid="1728" externalid="378818">
              <RESULTS>
                <RESULT eventid="1096" points="435" swimtime="00:00:59.14" resultid="1729" heatid="2021" lane="4" entrytime="00:00:59.21" entrycourse="SCM" />
                <RESULT eventid="1184" points="320" swimtime="00:00:36.47" resultid="1730" heatid="2055" lane="1" />
                <RESULT eventid="1200" points="470" swimtime="00:04:32.88" resultid="1731" heatid="2063" lane="2" entrytime="00:04:32.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                    <SPLIT distance="150" swimtime="00:01:40.31" />
                    <SPLIT distance="200" swimtime="00:02:15.65" />
                    <SPLIT distance="250" swimtime="00:02:50.28" />
                    <SPLIT distance="300" swimtime="00:03:24.57" />
                    <SPLIT distance="350" swimtime="00:03:58.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="335" swimtime="00:01:19.59" resultid="1732" heatid="2075" lane="1" entrytime="00:01:15.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="355" swimtime="00:00:28.45" resultid="1733" heatid="2109" lane="5" entrytime="00:00:28.14" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Claudio" lastname="Rohnelt" birthdate="2010-03-08" gender="M" nation="BRA" license="357954" swrid="5596935" athleteid="1663" externalid="357954">
              <RESULTS>
                <RESULT eventid="1096" points="332" swimtime="00:01:04.73" resultid="1664" heatid="2019" lane="5" entrytime="00:01:09.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="299" swimtime="00:01:11.39" resultid="1665" heatid="2050" lane="3" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="338" swimtime="00:05:04.47" resultid="1666" heatid="2062" lane="2" entrytime="00:04:59.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                    <SPLIT distance="100" swimtime="00:01:08.55" />
                    <SPLIT distance="150" swimtime="00:01:46.59" />
                    <SPLIT distance="200" swimtime="00:02:25.68" />
                    <SPLIT distance="250" swimtime="00:03:05.15" />
                    <SPLIT distance="300" swimtime="00:03:45.09" />
                    <SPLIT distance="350" swimtime="00:04:25.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="262" swimtime="00:00:33.96" resultid="1667" heatid="2081" lane="6" entrytime="00:00:33.63" entrycourse="SCM" />
                <RESULT eventid="1310" points="309" swimtime="00:00:29.80" resultid="1668" heatid="2108" lane="5" entrytime="00:00:30.71" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Henrique Marca Dos Santos" birthdate="2015-03-28" gender="M" nation="BRA" license="406695" swrid="4991165" athleteid="1847" externalid="406695">
              <RESULTS>
                <RESULT eventid="1113" points="121" swimtime="00:01:30.46" resultid="1848" heatid="2029" lane="1" entrytime="00:02:02.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="119" swimtime="00:00:44.85" resultid="1849" heatid="2046" lane="3" entrytime="00:00:42.73" entrycourse="SCM" />
                <RESULT eventid="1215" points="133" swimtime="00:00:42.56" resultid="1850" heatid="2068" lane="2" entrytime="00:00:47.73" entrycourse="SCM" />
                <RESULT eventid="1293" points="143" swimtime="00:00:38.53" resultid="1851" heatid="2097" lane="4" entrytime="00:00:37.21" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Luisa Lottermann" birthdate="2011-08-26" gender="F" nation="BRA" license="382238" swrid="5596909" athleteid="1744" externalid="382238">
              <RESULTS>
                <RESULT eventid="1060" points="331" swimtime="00:02:56.00" resultid="1745" heatid="2002" lane="3" entrytime="00:03:01.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.78" />
                    <SPLIT distance="100" swimtime="00:01:31.31" />
                    <SPLIT distance="150" swimtime="00:02:16.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="248" swimtime="00:01:19.98" resultid="1746" heatid="2013" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="214" swimtime="00:01:30.36" resultid="1747" heatid="2047" lane="2" entrytime="00:01:40.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="365" swimtime="00:05:23.58" resultid="1748" heatid="2058" lane="5" entrytime="00:05:53.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:01:17.84" />
                    <SPLIT distance="150" swimtime="00:01:58.92" />
                    <SPLIT distance="200" swimtime="00:02:40.49" />
                    <SPLIT distance="250" swimtime="00:03:21.21" />
                    <SPLIT distance="300" swimtime="00:04:01.78" />
                    <SPLIT distance="350" swimtime="00:04:42.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="327" swimtime="00:01:30.46" resultid="1749" heatid="2072" lane="2" entrytime="00:01:28.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Gamero Prado" birthdate="2007-05-16" gender="F" nation="BRA" license="305973" swrid="5596903" athleteid="1624" externalid="305973">
              <RESULTS>
                <RESULT eventid="1060" points="334" swimtime="00:02:55.47" resultid="1625" heatid="2003" lane="2" entrytime="00:02:50.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                    <SPLIT distance="100" swimtime="00:01:19.42" />
                    <SPLIT distance="150" swimtime="00:02:14.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="386" swimtime="00:01:08.98" resultid="1626" heatid="2016" lane="4" entrytime="00:01:06.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="354" swimtime="00:01:16.36" resultid="1627" heatid="2048" lane="3" entrytime="00:01:14.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="459" swimtime="00:04:59.68" resultid="1628" heatid="2060" lane="2" entrytime="00:05:00.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:10.56" />
                    <SPLIT distance="150" swimtime="00:01:48.49" />
                    <SPLIT distance="200" swimtime="00:02:26.43" />
                    <SPLIT distance="250" swimtime="00:03:04.48" />
                    <SPLIT distance="300" swimtime="00:03:42.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1244" points="384" swimtime="00:00:33.54" resultid="1629" heatid="2076" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Sehn Uren" birthdate="2009-10-15" gender="F" nation="BRA" license="357159" swrid="5596937" athleteid="1651" externalid="357159">
              <RESULTS>
                <RESULT eventid="1088" status="DNS" swimtime="00:00:00.00" resultid="1652" heatid="2015" lane="1" entrytime="00:01:10.03" entrycourse="SCM" />
                <RESULT eventid="1132" status="DNS" swimtime="00:00:00.00" resultid="1653" heatid="2034" lane="1" entrytime="00:00:37.26" entrycourse="SCM" />
                <RESULT eventid="1192" status="DNS" swimtime="00:00:00.00" resultid="1654" heatid="2058" lane="3" entrytime="00:05:35.98" entrycourse="SCM" />
                <RESULT eventid="1244" status="DNS" swimtime="00:00:00.00" resultid="1655" heatid="2078" lane="2" entrytime="00:00:35.07" entrycourse="SCM" />
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="1656" heatid="2104" lane="3" entrytime="00:00:32.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Vieira Rohnelt" birthdate="2012-05-03" gender="M" nation="BRA" license="365692" swrid="5588952" athleteid="1687" externalid="365692">
              <RESULTS>
                <RESULT eventid="1079" points="171" swimtime="00:01:39.58" resultid="1688" heatid="2008" lane="4" entrytime="00:01:41.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="217" swimtime="00:02:45.25" resultid="1689" heatid="2025" lane="5" entrytime="00:02:51.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:01:20.27" />
                    <SPLIT distance="150" swimtime="00:02:04.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1221" points="143" swimtime="00:01:31.27" resultid="1690" heatid="2070" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="196" swimtime="00:00:34.70" resultid="1691" heatid="2102" lane="6" entrytime="00:00:36.49" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Vargas Moreira" birthdate="2014-03-09" gender="F" nation="BRA" license="392014" swrid="4904290" athleteid="1820" externalid="392014">
              <RESULTS>
                <RESULT eventid="1110" points="275" swimtime="00:01:17.27" resultid="1821" heatid="2027" lane="4" entrytime="00:01:21.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1154" points="169" swimtime="00:00:45.65" resultid="1822" heatid="2044" lane="4" entrytime="00:00:47.45" entrycourse="SCM" />
                <RESULT eventid="1212" points="156" swimtime="00:00:45.25" resultid="1823" heatid="2066" lane="2" entrytime="00:00:51.09" entrycourse="SCM" />
                <RESULT eventid="1290" points="255" swimtime="00:00:36.15" resultid="1824" heatid="2094" lane="1" entrytime="00:00:40.59" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Henrique Wiebbeling" birthdate="2003-08-06" gender="M" nation="BRA" license="290420" swrid="4471225" athleteid="1609" externalid="290420">
              <RESULTS>
                <RESULT eventid="1124" points="477" swimtime="00:18:03.22" resultid="1610" heatid="2031" lane="4" entrytime="00:17:34.10" entrycourse="SCM" />
                <RESULT eventid="1140" points="335" swimtime="00:00:31.82" resultid="1611" heatid="2035" lane="3" />
                <RESULT eventid="1200" points="478" swimtime="00:04:31.40" resultid="1612" heatid="2064" lane="5" entrytime="00:04:21.56" entrycourse="SCM" />
                <RESULT eventid="1278" status="DNS" swimtime="00:00:00.00" resultid="1613" heatid="2090" lane="6" entrytime="00:01:07.46" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Gaio" birthdate="2012-11-13" gender="F" nation="BRA" license="390842" swrid="5596901" athleteid="1793" externalid="390842">
              <RESULTS>
                <RESULT eventid="1104" points="114" swimtime="00:03:47.42" resultid="1794" heatid="2023" lane="1" entrytime="00:04:24.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.37" />
                    <SPLIT distance="100" swimtime="00:01:50.00" />
                    <SPLIT distance="150" swimtime="00:02:51.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="80" swimtime="00:00:58.36" resultid="1795" heatid="2039" lane="5" entrytime="00:00:55.99" entrycourse="SCM" />
                <RESULT eventid="1218" points="72" swimtime="00:02:09.73" resultid="1796" heatid="2069" lane="4" entrytime="00:02:34.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="125" swimtime="00:00:45.83" resultid="1797" heatid="2098" lane="3" entrytime="00:00:44.93" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hendrik" lastname="Alteiro Groenwold" birthdate="2011-03-23" gender="M" nation="BRA" license="365756" swrid="5588520" athleteid="1675" externalid="365756">
              <RESULTS>
                <RESULT eventid="1068" points="385" swimtime="00:02:30.58" resultid="1676" heatid="2004" lane="3" entrytime="00:02:38.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:10.61" />
                    <SPLIT distance="150" swimtime="00:01:57.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="391" swimtime="00:01:01.29" resultid="1677" heatid="2020" lane="6" entrytime="00:01:04.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="302" swimtime="00:00:32.94" resultid="1678" heatid="2036" lane="5" />
                <RESULT eventid="1200" points="424" swimtime="00:04:42.48" resultid="1679" heatid="2062" lane="4" entrytime="00:04:43.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="100" swimtime="00:01:07.29" />
                    <SPLIT distance="150" swimtime="00:01:42.39" />
                    <SPLIT distance="200" swimtime="00:02:18.80" />
                    <SPLIT distance="250" swimtime="00:02:55.43" />
                    <SPLIT distance="300" swimtime="00:03:31.54" />
                    <SPLIT distance="350" swimtime="00:04:07.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="350" swimtime="00:00:28.58" resultid="1680" heatid="2106" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Borille Busetti" birthdate="2010-02-17" gender="F" nation="BRA" license="392830" swrid="5622263" athleteid="1836" externalid="392830">
              <RESULTS>
                <RESULT eventid="1088" points="394" swimtime="00:01:08.51" resultid="1837" heatid="2015" lane="2" entrytime="00:01:08.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="293" swimtime="00:00:37.99" resultid="1838" heatid="2033" lane="5" />
                <RESULT eventid="1192" points="324" swimtime="00:05:36.43" resultid="1839" heatid="2059" lane="6" entrytime="00:05:33.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                    <SPLIT distance="100" swimtime="00:01:17.77" />
                    <SPLIT distance="150" swimtime="00:02:00.82" />
                    <SPLIT distance="200" swimtime="00:02:43.59" />
                    <SPLIT distance="250" swimtime="00:03:27.48" />
                    <SPLIT distance="300" swimtime="00:04:11.57" />
                    <SPLIT distance="350" swimtime="00:04:54.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1270" points="283" swimtime="00:01:23.52" resultid="1840" heatid="2086" lane="4" entrytime="00:01:25.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="384" swimtime="00:00:31.52" resultid="1841" heatid="2103" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Kloeckner Feracin" birthdate="2014-03-21" gender="M" nation="BRA" license="414002" athleteid="1887" externalid="414002">
              <RESULTS>
                <RESULT eventid="1113" points="85" swimtime="00:01:41.90" resultid="1888" heatid="2029" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1157" points="79" swimtime="00:00:51.42" resultid="1889" heatid="2045" lane="3" />
                <RESULT eventid="1293" points="77" swimtime="00:00:47.19" resultid="1890" heatid="2096" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gael" lastname="Vicenzo Pereira" birthdate="2012-09-18" gender="M" nation="BRA" license="390847" swrid="5596943" athleteid="1809" externalid="390847">
              <RESULTS>
                <RESULT eventid="1079" points="52" swimtime="00:02:27.86" resultid="1810" heatid="2007" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="98" swimtime="00:03:35.17" resultid="1811" heatid="2024" lane="3" entrytime="00:03:57.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.64" />
                    <SPLIT distance="100" swimtime="00:01:41.92" />
                    <SPLIT distance="150" swimtime="00:02:37.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1221" points="47" swimtime="00:02:11.64" resultid="1812" heatid="2070" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="127" swimtime="00:00:40.09" resultid="1813" heatid="2100" lane="3" entrytime="00:00:48.04" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose" lastname="Eliziario Filho" birthdate="2014-03-27" gender="M" nation="BRA" license="406696" swrid="4979701" athleteid="1852" externalid="406696">
              <RESULTS>
                <RESULT eventid="1085" points="92" swimtime="00:00:55.22" resultid="1853" heatid="2011" lane="6" />
                <RESULT eventid="1113" points="150" swimtime="00:01:24.33" resultid="1854" heatid="2029" lane="4" entrytime="00:01:26.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="127" swimtime="00:00:43.20" resultid="1855" heatid="2068" lane="3" entrytime="00:00:41.60" entrycourse="SCM" />
                <RESULT eventid="1293" points="125" swimtime="00:00:40.30" resultid="1856" heatid="2097" lane="2" entrytime="00:00:39.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Rinaldini" birthdate="2009-04-09" gender="M" nation="BRA" license="348289" swrid="5596932" athleteid="1641" externalid="348289">
              <RESULTS>
                <RESULT eventid="1096" points="459" swimtime="00:00:58.10" resultid="1642" heatid="2021" lane="3" entrytime="00:00:59.05" entrycourse="SCM" />
                <RESULT eventid="1124" points="545" swimtime="00:17:16.78" resultid="1643" heatid="2031" lane="3" entrytime="00:17:23.57" entrycourse="SCM" />
                <RESULT eventid="1200" points="551" swimtime="00:04:18.86" resultid="1644" heatid="2064" lane="1" entrytime="00:04:22.48" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Balduíno" birthdate="2009-06-24" gender="M" nation="BRA" license="370764" swrid="5596870" athleteid="1722" externalid="370764">
              <RESULTS>
                <RESULT eventid="1096" points="465" swimtime="00:00:57.87" resultid="1723" heatid="2017" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="444" swimtime="00:01:02.61" resultid="1724" heatid="2051" lane="2" entrytime="00:01:04.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="471" swimtime="00:04:32.74" resultid="1725" heatid="2063" lane="6" entrytime="00:04:41.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:05.69" />
                    <SPLIT distance="150" swimtime="00:01:40.28" />
                    <SPLIT distance="200" swimtime="00:02:14.93" />
                    <SPLIT distance="250" swimtime="00:02:49.76" />
                    <SPLIT distance="300" swimtime="00:03:24.65" />
                    <SPLIT distance="350" swimtime="00:03:59.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="451" swimtime="00:00:28.36" resultid="1726" heatid="2080" lane="2" />
                <RESULT eventid="1310" points="251" swimtime="00:00:31.95" resultid="1727" heatid="2107" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Macedo Medeiros" birthdate="2012-05-12" gender="M" nation="BRA" license="392015" swrid="4697574" athleteid="1825" externalid="392015">
              <RESULTS>
                <RESULT eventid="1079" points="182" swimtime="00:01:37.52" resultid="1826" heatid="2008" lane="2" entrytime="00:01:55.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="119" swimtime="00:00:44.86" resultid="1827" heatid="2041" lane="3" entrytime="00:00:52.14" entrycourse="SCM" />
                <RESULT eventid="1267" points="140" swimtime="00:01:34.71" resultid="1828" heatid="2085" lane="4" entrytime="00:01:39.06" entrycourse="SCM" />
                <RESULT eventid="1299" points="165" swimtime="00:00:36.72" resultid="1829" heatid="2100" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Colaco Da Conceicao" birthdate="2011-05-25" gender="F" nation="BRA" license="369535" swrid="5588601" athleteid="1710" externalid="369535">
              <RESULTS>
                <RESULT eventid="1060" points="382" swimtime="00:02:47.86" resultid="1711" heatid="2003" lane="3" entrytime="00:02:47.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                    <SPLIT distance="100" swimtime="00:01:22.61" />
                    <SPLIT distance="150" swimtime="00:02:11.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="399" swimtime="00:01:08.20" resultid="1712" heatid="2013" lane="4" />
                <RESULT eventid="1160" points="278" swimtime="00:01:22.77" resultid="1713" heatid="2047" lane="3" entrytime="00:01:29.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="471" swimtime="00:04:57.27" resultid="1714" heatid="2060" lane="6" entrytime="00:05:02.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                    <SPLIT distance="100" swimtime="00:01:11.54" />
                    <SPLIT distance="150" swimtime="00:01:49.19" />
                    <SPLIT distance="200" swimtime="00:02:27.01" />
                    <SPLIT distance="250" swimtime="00:03:04.09" />
                    <SPLIT distance="300" swimtime="00:03:42.28" />
                    <SPLIT distance="350" swimtime="00:04:19.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1244" points="260" swimtime="00:00:38.18" resultid="1715" heatid="2077" lane="4" entrytime="00:00:40.06" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emanuel" lastname="Ranieri" birthdate="2011-01-24" gender="M" nation="BRA" license="390838" swrid="5596930" athleteid="1777" externalid="390838">
              <RESULTS>
                <RESULT eventid="1068" status="DSQ" swimtime="00:02:38.77" resultid="1778" heatid="2004" lane="2" entrytime="00:02:44.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                    <SPLIT distance="100" swimtime="00:01:15.90" />
                    <SPLIT distance="150" swimtime="00:02:03.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="338" swimtime="00:01:04.32" resultid="1779" heatid="2019" lane="4" entrytime="00:01:05.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="218" swimtime="00:01:19.27" resultid="1780" heatid="2049" lane="3" entrytime="00:01:32.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="344" swimtime="00:05:02.75" resultid="1781" heatid="2061" lane="4" entrytime="00:05:19.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                    <SPLIT distance="100" swimtime="00:01:12.65" />
                    <SPLIT distance="150" swimtime="00:01:51.62" />
                    <SPLIT distance="200" swimtime="00:02:30.14" />
                    <SPLIT distance="250" swimtime="00:03:09.24" />
                    <SPLIT distance="300" swimtime="00:03:48.21" />
                    <SPLIT distance="350" swimtime="00:04:26.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="230" swimtime="00:01:18.83" resultid="1782" heatid="2089" lane="5" entrytime="00:01:17.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Zimmermann" birthdate="2010-01-19" gender="M" nation="BRA" license="357160" swrid="5588977" athleteid="1657" externalid="357160">
              <RESULTS>
                <RESULT eventid="1096" points="473" swimtime="00:00:57.52" resultid="1658" heatid="2021" lane="6" entrytime="00:00:59.63" entrycourse="SCM" />
                <RESULT eventid="1140" points="364" swimtime="00:00:30.96" resultid="1659" heatid="2035" lane="4" />
                <RESULT eventid="1200" points="516" swimtime="00:04:24.47" resultid="1660" heatid="2064" lane="2" entrytime="00:04:20.92" entrycourse="SCM" />
                <RESULT eventid="1236" points="352" swimtime="00:01:18.23" resultid="1661" heatid="2075" lane="6" entrytime="00:01:17.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="411" swimtime="00:00:27.11" resultid="1662" heatid="2109" lane="2" entrytime="00:00:27.71" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Menegazzi Daga" birthdate="2014-12-05" gender="M" nation="BRA" license="414003" athleteid="1891" externalid="414003">
              <RESULTS>
                <RESULT eventid="1085" points="63" swimtime="00:01:02.48" resultid="1892" heatid="2011" lane="1" />
                <RESULT eventid="1157" points="53" swimtime="00:00:58.51" resultid="1893" heatid="2045" lane="4" />
                <RESULT eventid="1293" points="63" swimtime="00:00:50.46" resultid="1894" heatid="2095" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Stein Duarte" birthdate="2010-10-03" gender="F" nation="BRA" license="351635" swrid="5588923" athleteid="1645" externalid="351635">
              <RESULTS>
                <RESULT eventid="1088" points="439" swimtime="00:01:06.10" resultid="1646" heatid="2015" lane="6" entrytime="00:01:10.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="328" swimtime="00:01:18.31" resultid="1647" heatid="2048" lane="2" entrytime="00:01:23.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="425" swimtime="00:05:07.47" resultid="1648" heatid="2059" lane="3" entrytime="00:05:09.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="100" swimtime="00:01:12.32" />
                    <SPLIT distance="150" swimtime="00:01:50.74" />
                    <SPLIT distance="200" swimtime="00:02:30.03" />
                    <SPLIT distance="250" swimtime="00:03:09.04" />
                    <SPLIT distance="300" swimtime="00:03:48.38" />
                    <SPLIT distance="350" swimtime="00:04:28.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1244" points="341" swimtime="00:00:34.87" resultid="1649" heatid="2077" lane="5" />
                <RESULT eventid="1302" points="392" swimtime="00:00:31.33" resultid="1650" heatid="2103" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Paese Worm" birthdate="2014-07-23" gender="F" nation="BRA" license="380655" swrid="5596920" athleteid="1734" externalid="380655">
              <RESULTS>
                <RESULT eventid="1082" points="119" swimtime="00:00:57.61" resultid="1735" heatid="2010" lane="1" entrytime="00:00:55.57" entrycourse="SCM" />
                <RESULT eventid="1154" points="121" swimtime="00:00:51.01" resultid="1736" heatid="2044" lane="2" entrytime="00:00:48.30" entrycourse="SCM" />
                <RESULT eventid="1212" points="109" swimtime="00:00:50.97" resultid="1737" heatid="2065" lane="2" />
                <RESULT eventid="1290" points="187" swimtime="00:00:40.07" resultid="1738" heatid="2093" lane="4" entrytime="00:00:45.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Paiz Ribeiro" birthdate="2006-02-17" gender="M" nation="BRA" license="297583" swrid="5596921" athleteid="1614" externalid="297583">
              <RESULTS>
                <RESULT eventid="1096" points="455" swimtime="00:00:58.28" resultid="1615" heatid="2017" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="480" swimtime="00:01:01.00" resultid="1616" heatid="2051" lane="3" entrytime="00:01:00.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="510" swimtime="00:04:25.56" resultid="1617" heatid="2063" lane="4" entrytime="00:04:30.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.02" />
                    <SPLIT distance="100" swimtime="00:01:02.89" />
                    <SPLIT distance="150" swimtime="00:01:36.10" />
                    <SPLIT distance="200" swimtime="00:02:09.81" />
                    <SPLIT distance="250" swimtime="00:02:43.49" />
                    <SPLIT distance="300" swimtime="00:03:17.96" />
                    <SPLIT distance="350" swimtime="00:03:52.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="400" swimtime="00:01:15.02" resultid="1618" heatid="2075" lane="2" entrytime="00:01:12.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="343" swimtime="00:01:08.99" resultid="1619" heatid="2089" lane="4" entrytime="00:01:09.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Dillenburg Benetti" birthdate="2011-03-10" gender="M" nation="BRA" license="368119" swrid="5588656" athleteid="1681" externalid="368119">
              <RESULTS>
                <RESULT eventid="1068" points="340" swimtime="00:02:37.04" resultid="1682" heatid="2004" lane="4" entrytime="00:02:38.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="100" swimtime="00:01:15.88" />
                    <SPLIT distance="150" swimtime="00:02:03.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="347" swimtime="00:01:03.75" resultid="1683" heatid="2019" lane="3" entrytime="00:01:05.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="205" swimtime="00:01:20.98" resultid="1684" heatid="2050" lane="1" entrytime="00:01:23.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="383" swimtime="00:04:52.07" resultid="1685" heatid="2062" lane="6" entrytime="00:05:10.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:09.97" />
                    <SPLIT distance="150" swimtime="00:01:46.15" />
                    <SPLIT distance="200" swimtime="00:02:23.20" />
                    <SPLIT distance="250" swimtime="00:03:01.11" />
                    <SPLIT distance="300" swimtime="00:03:38.39" />
                    <SPLIT distance="350" swimtime="00:04:15.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="302" swimtime="00:01:11.97" resultid="1686" heatid="2089" lane="2" entrytime="00:01:10.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="1903" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Felipe" lastname="Arend Fiedler" birthdate="2015-06-26" gender="M" nation="BRA" license="414195" athleteid="1931" externalid="414195">
              <RESULTS>
                <RESULT eventid="1085" points="33" swimtime="00:01:17.75" resultid="1932" heatid="2011" lane="5" />
                <RESULT eventid="1157" points="46" swimtime="00:01:01.69" resultid="1933" heatid="2045" lane="2" />
                <RESULT eventid="1293" points="31" swimtime="00:01:04.09" resultid="1934" heatid="2095" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Schneider Paz" birthdate="2011-07-03" gender="M" nation="BRA" license="412899" athleteid="1913" externalid="412899">
              <RESULTS>
                <RESULT eventid="1096" points="183" swimtime="00:01:18.97" resultid="1914" heatid="2017" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="194" swimtime="00:00:43.03" resultid="1915" heatid="2054" lane="3" />
                <RESULT eventid="1252" points="175" swimtime="00:00:38.83" resultid="1916" heatid="2080" lane="5" />
                <RESULT eventid="1310" points="206" swimtime="00:00:34.09" resultid="1917" heatid="2107" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Laura Oliveira" birthdate="2014-05-19" gender="F" nation="BRA" license="414179" athleteid="1923" externalid="414179">
              <RESULTS>
                <RESULT eventid="1110" points="93" swimtime="00:01:50.53" resultid="1924" heatid="2026" lane="2" />
                <RESULT eventid="1154" points="87" swimtime="00:00:56.86" resultid="1925" heatid="2043" lane="2" />
                <RESULT eventid="1290" points="117" swimtime="00:00:46.77" resultid="1926" heatid="2092" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiggi" lastname="Frasson Abreu" birthdate="2014-07-16" gender="M" nation="BRA" license="411413" athleteid="1909" externalid="411413">
              <RESULTS>
                <RESULT eventid="1085" points="60" swimtime="00:01:03.66" resultid="1910" heatid="2011" lane="3" />
                <RESULT eventid="1157" points="41" swimtime="00:01:04.12" resultid="1911" heatid="2046" lane="2" />
                <RESULT eventid="1293" points="47" swimtime="00:00:55.76" resultid="1912" heatid="2096" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Schneider Paz" birthdate="2010-04-21" gender="M" nation="BRA" license="412900" athleteid="1918" externalid="412900">
              <RESULTS>
                <RESULT eventid="1096" points="152" swimtime="00:01:24.00" resultid="1919" heatid="2018" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="168" swimtime="00:00:45.19" resultid="1920" heatid="2055" lane="2" />
                <RESULT eventid="1236" points="142" swimtime="00:01:45.77" resultid="1921" heatid="2073" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="159" swimtime="00:00:37.21" resultid="1922" heatid="2107" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Vitoria Loh" birthdate="2015-08-31" gender="F" nation="BRA" license="414180" athleteid="1927" externalid="414180">
              <RESULTS>
                <RESULT eventid="1082" points="51" swimtime="00:01:16.23" resultid="1928" heatid="2009" lane="5" />
                <RESULT eventid="1154" points="69" swimtime="00:01:01.29" resultid="1929" heatid="2043" lane="5" />
                <RESULT eventid="1290" points="55" swimtime="00:01:00.08" resultid="1930" heatid="2092" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Voltarelli Souza" birthdate="2014-07-26" gender="M" nation="BRA" license="410202" swrid="5748710" athleteid="1904" externalid="410202">
              <RESULTS>
                <RESULT eventid="1085" points="101" swimtime="00:00:53.53" resultid="1905" heatid="2012" lane="2" entrytime="00:00:52.90" entrycourse="SCM" />
                <RESULT eventid="1113" points="88" swimtime="00:01:40.67" resultid="1906" heatid="2028" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="84" swimtime="00:00:49.48" resultid="1907" heatid="2067" lane="4" />
                <RESULT eventid="1293" points="107" swimtime="00:00:42.34" resultid="1908" heatid="2097" lane="1" entrytime="00:00:41.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3133" nation="BRA" region="PR" clubid="1935" swrid="93768" name="Associação Toledo Natação" shortname="Toledo Natação">
          <ATHLETES>
            <ATHLETE firstname="Gabriel" lastname="Marafon" birthdate="2006-06-17" gender="M" nation="BRA" license="380288" swrid="5622291" athleteid="1954" externalid="380288">
              <RESULTS>
                <RESULT eventid="1096" points="414" swimtime="00:01:00.15" resultid="1955" heatid="2021" lane="1" entrytime="00:00:59.58" entrycourse="SCM" />
                <RESULT eventid="1184" points="441" swimtime="00:00:32.77" resultid="1956" heatid="2056" lane="4" entrytime="00:00:32.77" entrycourse="SCM" />
                <RESULT eventid="1236" points="441" swimtime="00:01:12.59" resultid="1957" heatid="2075" lane="3" entrytime="00:01:11.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="277" swimtime="00:00:33.33" resultid="1958" heatid="2079" lane="4" />
                <RESULT eventid="1310" points="402" swimtime="00:00:27.31" resultid="1959" heatid="2109" lane="4" entrytime="00:00:26.99" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giullia" lastname="Lagni" birthdate="2006-11-22" gender="F" nation="BRA" license="337671" swrid="5622285" athleteid="1948" externalid="337671">
              <RESULTS>
                <RESULT eventid="1088" points="328" swimtime="00:01:12.83" resultid="1949" heatid="2015" lane="5" entrytime="00:01:09.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="282" swimtime="00:00:38.49" resultid="1950" heatid="2034" lane="2" entrytime="00:00:36.28" entrycourse="SCM" />
                <RESULT eventid="1244" points="233" swimtime="00:00:39.59" resultid="1951" heatid="2077" lane="1" />
                <RESULT eventid="1270" points="283" swimtime="00:01:23.54" resultid="1952" heatid="2087" lane="5" entrytime="00:01:16.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="313" swimtime="00:00:33.75" resultid="1953" heatid="2105" lane="1" entrytime="00:00:31.62" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Torres Romancini" birthdate="2010-05-28" gender="F" nation="BRA" license="347218" swrid="5622309" athleteid="1960" externalid="347218">
              <RESULTS>
                <RESULT eventid="1088" points="370" swimtime="00:01:09.94" resultid="1961" heatid="2014" lane="4" entrytime="00:01:12.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="420" swimtime="00:00:33.71" resultid="1962" heatid="2034" lane="4" entrytime="00:00:33.68" entrycourse="SCM" />
                <RESULT eventid="1192" points="356" swimtime="00:05:26.19" resultid="1963" heatid="2057" lane="2" />
                <RESULT eventid="1244" points="378" swimtime="00:00:33.71" resultid="1964" heatid="2078" lane="3" entrytime="00:00:33.64" entrycourse="SCM" />
                <RESULT eventid="1270" points="382" swimtime="00:01:15.59" resultid="1965" heatid="2087" lane="4" entrytime="00:01:13.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Fernando Braga Da Silva" birthdate="2011-01-10" gender="M" nation="BRA" license="380291" swrid="5453344" athleteid="1984" externalid="380291">
              <RESULTS>
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="1985" heatid="2018" lane="4" entrytime="00:01:17.56" entrycourse="SCM" />
                <RESULT eventid="1140" status="DNS" swimtime="00:00:00.00" resultid="1986" heatid="2037" lane="6" entrytime="00:00:40.33" entrycourse="SCM" />
                <RESULT eventid="1184" status="DNS" swimtime="00:00:00.00" resultid="1987" heatid="2055" lane="3" entrytime="00:00:49.94" entrycourse="SCM" />
                <RESULT eventid="1236" status="DNS" swimtime="00:00:00.00" resultid="1988" heatid="2073" lane="4" />
                <RESULT eventid="1310" status="DNS" swimtime="00:00:00.00" resultid="1989" heatid="2107" lane="4" entrytime="00:00:35.71" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Marafon" birthdate="2011-03-23" gender="F" nation="BRA" license="380287" swrid="5652623" athleteid="1978" externalid="380287">
              <RESULTS>
                <RESULT eventid="1088" points="357" swimtime="00:01:10.81" resultid="1979" heatid="2015" lane="4" entrytime="00:01:07.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="371" swimtime="00:00:39.48" resultid="1980" heatid="2053" lane="3" entrytime="00:00:38.58" entrycourse="SCM" />
                <RESULT eventid="1192" points="323" swimtime="00:05:36.78" resultid="1981" heatid="2057" lane="4" />
                <RESULT eventid="1244" points="302" swimtime="00:00:36.32" resultid="1982" heatid="2077" lane="2" entrytime="00:00:40.33" entrycourse="SCM" />
                <RESULT eventid="1302" points="374" swimtime="00:00:31.82" resultid="1983" heatid="2105" lane="2" entrytime="00:00:30.93" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lavinia" lastname="Martins Paludo" birthdate="2010-09-30" gender="F" nation="BRA" license="347217" swrid="5652624" athleteid="1966" externalid="347217">
              <RESULTS>
                <RESULT eventid="1060" points="195" swimtime="00:03:29.84" resultid="1967" heatid="2002" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.16" />
                    <SPLIT distance="100" swimtime="00:01:44.13" />
                    <SPLIT distance="150" swimtime="00:02:40.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="225" swimtime="00:01:22.53" resultid="1968" heatid="2014" lane="5" entrytime="00:01:15.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="221" swimtime="00:00:46.88" resultid="1969" heatid="2053" lane="5" entrytime="00:00:44.97" entrycourse="SCM" />
                <RESULT eventid="1192" points="217" swimtime="00:06:24.69" resultid="1970" heatid="2057" lane="3" />
                <RESULT eventid="1228" points="214" swimtime="00:01:44.17" resultid="1971" heatid="2072" lane="1" entrytime="00:01:38.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Feder" birthdate="2008-11-13" gender="M" nation="BRA" license="347224" swrid="5622278" athleteid="1936" externalid="347224">
              <RESULTS>
                <RESULT eventid="1096" points="379" swimtime="00:01:01.92" resultid="1937" heatid="2020" lane="3" entrytime="00:00:59.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="398" swimtime="00:00:30.04" resultid="1938" heatid="2037" lane="2" entrytime="00:00:29.80" entrycourse="SCM" />
                <RESULT eventid="1168" points="290" swimtime="00:01:12.11" resultid="1939" heatid="2051" lane="1" entrytime="00:01:10.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="427" swimtime="00:00:28.87" resultid="1940" heatid="2081" lane="2" entrytime="00:00:30.32" entrycourse="SCM" />
                <RESULT eventid="1278" points="388" swimtime="00:01:06.24" resultid="1941" heatid="2090" lane="1" entrytime="00:01:05.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Pauly Follmann" birthdate="2011-04-19" gender="F" nation="BRA" license="413886" athleteid="1990" externalid="413886">
              <RESULTS>
                <RESULT eventid="1088" points="150" swimtime="00:01:34.43" resultid="1991" heatid="2013" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="181" swimtime="00:00:44.59" resultid="1992" heatid="2033" lane="4" entrytime="00:00:45.04" entrycourse="SCM" />
                <RESULT eventid="1176" points="177" swimtime="00:00:50.48" resultid="1993" heatid="2052" lane="1" />
                <RESULT eventid="1244" status="DSQ" swimtime="00:00:51.80" resultid="1994" heatid="2076" lane="2" />
                <RESULT eventid="1302" points="191" swimtime="00:00:39.77" resultid="1995" heatid="2103" lane="4" entrytime="00:00:43.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Welter Levandowski" birthdate="2011-05-06" gender="F" nation="BRA" license="380286" swrid="5652626" athleteid="1972" externalid="380286">
              <RESULTS>
                <RESULT eventid="1088" points="313" swimtime="00:01:13.98" resultid="1973" heatid="2013" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="298" swimtime="00:22:39.38" resultid="1974" heatid="2030" lane="2" />
                <RESULT eventid="1160" points="218" swimtime="00:01:29.78" resultid="1975" heatid="2048" lane="6" entrytime="00:01:26.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="330" swimtime="00:05:34.57" resultid="1976" heatid="2059" lane="1" entrytime="00:05:26.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.52" />
                    <SPLIT distance="100" swimtime="00:01:17.11" />
                    <SPLIT distance="150" swimtime="00:01:59.31" />
                    <SPLIT distance="200" swimtime="00:02:42.29" />
                    <SPLIT distance="250" swimtime="00:03:25.65" />
                    <SPLIT distance="300" swimtime="00:04:09.62" />
                    <SPLIT distance="350" swimtime="00:04:52.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1244" points="278" swimtime="00:00:37.35" resultid="1977" heatid="2078" lane="1" entrytime="00:00:35.82" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Marafon Duarte" birthdate="2011-08-18" gender="M" nation="BRA" license="414184" athleteid="1996" externalid="414184">
              <RESULTS>
                <RESULT eventid="1096" points="205" swimtime="00:01:15.93" resultid="1997" heatid="2017" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="125" swimtime="00:00:44.11" resultid="1998" heatid="2036" lane="4" />
                <RESULT eventid="1184" points="108" swimtime="00:00:52.28" resultid="1999" heatid="2054" lane="2" />
                <RESULT eventid="1236" points="143" swimtime="00:01:45.61" resultid="2000" heatid="2073" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="212" swimtime="00:00:33.78" resultid="2001" heatid="2106" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrielly" lastname="Luiza Horn" birthdate="2004-04-03" gender="F" nation="BRA" license="315145" swrid="5622288" athleteid="1942" externalid="315145">
              <RESULTS>
                <RESULT eventid="1132" points="346" swimtime="00:00:35.96" resultid="1943" heatid="2034" lane="5" entrytime="00:00:36.32" entrycourse="SCM" />
                <RESULT eventid="1160" points="253" swimtime="00:01:25.36" resultid="1944" heatid="2048" lane="4" entrytime="00:01:20.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="242" swimtime="00:00:45.52" resultid="1945" heatid="2053" lane="2" entrytime="00:00:40.16" entrycourse="SCM" />
                <RESULT eventid="1244" points="327" swimtime="00:00:35.37" resultid="1946" heatid="2078" lane="4" entrytime="00:00:33.69" entrycourse="SCM" />
                <RESULT eventid="1302" points="335" swimtime="00:00:32.99" resultid="1947" heatid="2105" lane="6" entrytime="00:00:32.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13025" nation="BRA" region="PR" clubid="1440" swrid="93779" name="Instituto Desportos Aquáticos De Foz Do Iguaçu" shortname="Cataratas Natação">
          <ATHLETES>
            <ATHLETE firstname="Benjamin" lastname="Perius Goncalves De Lima" birthdate="2016-06-09" gender="M" nation="BRA" license="407798" swrid="5721506" athleteid="1564" externalid="407798">
              <RESULTS>
                <RESULT eventid="1226" points="89" swimtime="00:00:23.01" resultid="1565" heatid="2071" lane="4" />
                <RESULT eventid="1262" points="88" swimtime="00:00:25.76" resultid="1566" heatid="2082" lane="4" />
                <RESULT eventid="1288" points="120" swimtime="00:00:18.39" resultid="1567" heatid="2091" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mayumi" lastname="Napole" birthdate="2010-02-01" gender="F" nation="BRA" license="376446" swrid="5596918" athleteid="1504" externalid="376446" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1116" points="271" swimtime="00:23:22.37" resultid="1505" heatid="2030" lane="5" />
                <RESULT eventid="1176" status="DNS" swimtime="00:00:00.00" resultid="1506" heatid="2052" lane="4" />
                <RESULT eventid="1192" points="329" swimtime="00:05:34.78" resultid="1507" heatid="2058" lane="2" entrytime="00:05:40.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                    <SPLIT distance="100" swimtime="00:01:17.95" />
                    <SPLIT distance="150" swimtime="00:02:00.08" />
                    <SPLIT distance="200" swimtime="00:02:43.25" />
                    <SPLIT distance="250" swimtime="00:03:26.14" />
                    <SPLIT distance="300" swimtime="00:04:09.88" />
                    <SPLIT distance="350" swimtime="00:04:52.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="392" swimtime="00:00:31.32" resultid="1508" heatid="2105" lane="5" entrytime="00:00:31.09" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Marques Petry" birthdate="2008-01-08" gender="M" nation="BRA" license="392352" swrid="4795316" athleteid="1470" externalid="392352" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1068" points="300" swimtime="00:02:43.72" resultid="1471" heatid="2004" lane="5" entrytime="00:02:45.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                    <SPLIT distance="100" swimtime="00:01:20.62" />
                    <SPLIT distance="150" swimtime="00:02:07.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="378" swimtime="00:01:01.99" resultid="1472" heatid="2020" lane="5" entrytime="00:01:02.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="342" swimtime="00:05:03.43" resultid="1473" heatid="2062" lane="1" entrytime="00:05:07.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                    <SPLIT distance="150" swimtime="00:01:47.64" />
                    <SPLIT distance="200" swimtime="00:02:26.28" />
                    <SPLIT distance="250" swimtime="00:03:05.82" />
                    <SPLIT distance="300" swimtime="00:03:45.48" />
                    <SPLIT distance="350" swimtime="00:04:25.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="341" swimtime="00:00:28.83" resultid="1474" heatid="2109" lane="1" entrytime="00:00:29.12" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Riam Nagorski De Lima" birthdate="2014-04-26" gender="M" nation="BRA" license="407802" swrid="5721507" athleteid="1580" externalid="407802">
              <RESULTS>
                <RESULT eventid="1085" points="67" swimtime="00:01:01.24" resultid="1581" heatid="2012" lane="1" entrytime="00:01:15.07" entrycourse="SCM" />
                <RESULT eventid="1113" points="83" swimtime="00:01:42.79" resultid="1582" heatid="2028" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1293" points="86" swimtime="00:00:45.53" resultid="1583" heatid="2096" lane="2" entrytime="00:00:56.21" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Laura Lima Belo" birthdate="2015-07-09" gender="F" nation="BRA" license="407801" swrid="5721501" athleteid="1577" externalid="407801">
              <RESULTS>
                <RESULT eventid="1110" points="49" swimtime="00:02:16.90" resultid="1578" heatid="2026" lane="4" />
                <RESULT eventid="1290" points="62" swimtime="00:00:57.85" resultid="1579" heatid="2092" lane="3" entrytime="00:01:12.23" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Carvalho Carelli" birthdate="2011-10-15" gender="M" nation="BRA" license="403146" swrid="5676300" athleteid="1529" externalid="403146" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1096" points="304" swimtime="00:01:06.65" resultid="1530" heatid="2019" lane="6" entrytime="00:01:09.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="282" swimtime="00:01:12.82" resultid="1531" heatid="2051" lane="6" entrytime="00:01:11.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1252" points="283" swimtime="00:00:33.11" resultid="1532" heatid="2081" lane="5" entrytime="00:00:32.78" entrycourse="SCM" />
                <RESULT eventid="1278" points="221" swimtime="00:01:19.84" resultid="1533" heatid="2088" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Abraao" lastname="Felipe Oliveira" birthdate="2012-05-20" gender="M" nation="BRA" license="400457" swrid="5420917" athleteid="1524" externalid="400457" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1107" points="146" swimtime="00:03:08.68" resultid="1525" heatid="2025" lane="6" entrytime="00:03:14.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.05" />
                    <SPLIT distance="100" swimtime="00:01:32.49" />
                    <SPLIT distance="150" swimtime="00:02:21.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="78" swimtime="00:00:51.62" resultid="1526" heatid="2042" lane="5" entrytime="00:00:48.15" entrycourse="SCM" />
                <RESULT eventid="1267" points="146" swimtime="00:01:33.44" resultid="1527" heatid="2085" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="189" swimtime="00:00:35.10" resultid="1528" heatid="2102" lane="5" entrytime="00:00:34.26" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Roza" birthdate="2013-06-05" gender="M" nation="BRA" license="374412" swrid="5588949" athleteid="1494" externalid="374412" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1107" points="233" swimtime="00:02:41.40" resultid="1495" heatid="2025" lane="2" entrytime="00:02:48.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:15.61" />
                    <SPLIT distance="150" swimtime="00:01:59.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" status="DSQ" swimtime="00:00:38.89" resultid="1496" heatid="2042" lane="3" entrytime="00:00:41.28" entrycourse="SCM" />
                <RESULT eventid="1221" points="160" swimtime="00:01:27.88" resultid="1497" heatid="2070" lane="4" entrytime="00:01:23.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="250" swimtime="00:00:32.00" resultid="1498" heatid="2102" lane="4" entrytime="00:00:31.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ayla" lastname="Corazza Boncompanho" birthdate="2015-10-13" gender="F" nation="BRA" license="414175" athleteid="1593" externalid="414175">
              <RESULTS>
                <RESULT eventid="1082" status="DNS" swimtime="00:00:00.00" resultid="1594" heatid="2009" lane="6" />
                <RESULT eventid="1154" status="DNS" swimtime="00:00:00.00" resultid="1595" heatid="2043" lane="3" />
                <RESULT eventid="1290" status="DNS" swimtime="00:00:00.00" resultid="1596" heatid="2092" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Ioris Souza" birthdate="2015-09-10" gender="F" nation="BRA" license="406693" swrid="5042791" athleteid="1559" externalid="406693" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1082" points="139" swimtime="00:00:54.69" resultid="1560" heatid="2010" lane="6" entrytime="00:01:03.44" entrycourse="SCM" />
                <RESULT eventid="1110" points="116" swimtime="00:01:42.93" resultid="1561" heatid="2026" lane="1" />
                <RESULT eventid="1212" points="120" swimtime="00:00:49.35" resultid="1562" heatid="2065" lane="4" />
                <RESULT eventid="1290" points="119" swimtime="00:00:46.60" resultid="1563" heatid="2093" lane="5" entrytime="00:00:53.17" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Kasprzak" birthdate="2011-08-09" gender="F" nation="BRA" license="406659" swrid="5073376" athleteid="1550" externalid="406659" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1088" points="154" swimtime="00:01:33.70" resultid="1551" heatid="2013" lane="3" entrytime="00:01:31.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="167" swimtime="00:00:45.81" resultid="1552" heatid="2032" lane="4" />
                <RESULT eventid="1176" points="182" swimtime="00:00:50.00" resultid="1553" heatid="2052" lane="3" entrytime="00:01:00.08" entrycourse="SCM" />
                <RESULT eventid="1302" points="169" swimtime="00:00:41.44" resultid="1554" heatid="2103" lane="3" entrytime="00:00:39.67" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Katherine" lastname="Kotz" birthdate="2012-05-18" gender="F" nation="BRA" license="390810" swrid="5596907" athleteid="1479" externalid="390810" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1076" points="244" swimtime="00:01:39.71" resultid="1480" heatid="2006" lane="4" entrytime="00:01:42.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="282" swimtime="00:02:48.08" resultid="1481" heatid="2023" lane="3" entrytime="00:02:45.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:01:24.19" />
                    <SPLIT distance="150" swimtime="00:02:08.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="251" swimtime="00:01:29.51" resultid="1482" heatid="2084" lane="3" entrytime="00:01:32.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="326" swimtime="00:00:33.29" resultid="1483" heatid="2099" lane="4" entrytime="00:00:32.56" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Bailke" birthdate="2007-05-04" gender="M" nation="BRA" license="370566" swrid="5596869" athleteid="1459" externalid="370566" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1124" points="314" swimtime="00:20:44.98" resultid="1460" heatid="2031" lane="1" entrytime="00:20:20.71" entrycourse="SCM" />
                <RESULT eventid="1252" points="319" swimtime="00:00:31.81" resultid="1461" heatid="2081" lane="1" entrytime="00:00:33.00" entrycourse="SCM" />
                <RESULT eventid="1310" points="360" swimtime="00:00:28.32" resultid="1462" heatid="2108" lane="3" entrytime="00:00:29.62" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Resende Ames" birthdate="2006-02-10" gender="M" nation="BRA" license="365657" swrid="5596931" athleteid="1444" externalid="365657" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1068" points="499" swimtime="00:02:18.20" resultid="1445" heatid="2005" lane="3" entrytime="00:02:20.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.21" />
                    <SPLIT distance="100" swimtime="00:01:02.91" />
                    <SPLIT distance="150" swimtime="00:01:48.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1200" points="249" swimtime="00:05:37.07" resultid="1446" heatid="2064" lane="4" entrytime="00:04:16.49" entrycourse="SCM" />
                <RESULT eventid="1310" points="484" swimtime="00:00:25.67" resultid="1447" heatid="2110" lane="2" entrytime="00:00:25.49" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Luiz Martinazzo" birthdate="2006-05-16" gender="M" nation="BRA" license="345593" swrid="5596910" athleteid="1453" externalid="345593" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1096" points="490" swimtime="00:00:56.84" resultid="1454" heatid="2022" lane="2" entrytime="00:00:56.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="372" swimtime="00:00:30.72" resultid="1455" heatid="2037" lane="4" entrytime="00:00:29.70" entrycourse="SCM" />
                <RESULT eventid="1184" points="321" swimtime="00:00:36.42" resultid="1456" heatid="2055" lane="6" />
                <RESULT eventid="1200" points="449" swimtime="00:04:37.01" resultid="1457" heatid="2064" lane="6" entrytime="00:04:28.15" entrycourse="SCM" />
                <RESULT eventid="1278" points="351" swimtime="00:01:08.49" resultid="1458" heatid="2090" lane="2" entrytime="00:01:03.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Ferrari Ghellere" birthdate="2014-07-01" gender="F" nation="BRA" license="372038" swrid="5596895" athleteid="1489" externalid="372038" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1110" points="256" swimtime="00:01:19.13" resultid="1490" heatid="2027" lane="3" entrytime="00:01:20.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1154" points="179" swimtime="00:00:44.75" resultid="1491" heatid="2044" lane="3" entrytime="00:00:45.03" entrycourse="SCM" />
                <RESULT eventid="1212" points="187" swimtime="00:00:42.61" resultid="1492" heatid="2066" lane="3" entrytime="00:00:41.03" entrycourse="SCM" />
                <RESULT eventid="1290" points="227" swimtime="00:00:37.56" resultid="1493" heatid="2094" lane="5" entrytime="00:00:40.46" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Lima Belo" birthdate="2012-10-07" gender="F" nation="BRA" license="407799" swrid="5721502" athleteid="1568" externalid="407799">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="1569" heatid="2006" lane="1" />
                <RESULT eventid="1104" points="113" swimtime="00:03:47.72" resultid="1570" heatid="2023" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.62" />
                    <SPLIT distance="100" swimtime="00:01:48.34" />
                    <SPLIT distance="150" swimtime="00:02:47.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="138" swimtime="00:00:44.28" resultid="1571" heatid="2099" lane="6" entrytime="00:00:42.58" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edward" lastname="Mikael De Lima" birthdate="2012-03-11" gender="M" nation="BRA" license="376445" swrid="5588816" athleteid="1499" externalid="376445" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1107" points="365" swimtime="00:02:19.01" resultid="1500" heatid="2025" lane="3" entrytime="00:02:18.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                    <SPLIT distance="100" swimtime="00:01:08.25" />
                    <SPLIT distance="150" swimtime="00:01:43.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1221" points="250" swimtime="00:01:15.79" resultid="1501" heatid="2070" lane="3" entrytime="00:01:15.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="289" swimtime="00:01:14.49" resultid="1502" heatid="2085" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="351" swimtime="00:00:28.56" resultid="1503" heatid="2102" lane="3" entrytime="00:00:27.35" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Resende Ames" birthdate="2010-02-02" gender="M" nation="BRA" license="365505" swrid="5588876" athleteid="1484" externalid="365505" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="1485" heatid="2021" lane="5" entrytime="00:00:59.51" entrycourse="SCM" />
                <RESULT eventid="1140" status="DNS" swimtime="00:00:00.00" resultid="1486" heatid="2037" lane="5" entrytime="00:00:31.15" entrycourse="SCM" />
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="1487" heatid="2050" lane="4" entrytime="00:01:13.05" entrycourse="SCM" />
                <RESULT eventid="1278" status="DNS" swimtime="00:00:00.00" resultid="1488" heatid="2090" lane="5" entrytime="00:01:05.13" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Marcio Peixoto" birthdate="2012-10-22" gender="M" nation="BRA" license="411994" swrid="5740013" athleteid="1584" externalid="411994">
              <RESULTS>
                <RESULT eventid="1107" points="98" swimtime="00:03:35.23" resultid="1585" heatid="2024" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.70" />
                    <SPLIT distance="100" swimtime="00:01:30.93" />
                    <SPLIT distance="150" swimtime="00:02:30.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="66" swimtime="00:00:54.44" resultid="1586" heatid="2042" lane="6" entrytime="00:00:51.48" entrycourse="SCM" />
                <RESULT eventid="1299" points="137" swimtime="00:00:39.03" resultid="1587" heatid="2101" lane="2" entrytime="00:00:39.70" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="De Souza" birthdate="2014-03-30" gender="M" nation="BRA" license="407800" swrid="5721499" athleteid="1572" externalid="407800">
              <RESULTS>
                <RESULT eventid="1085" points="140" swimtime="00:00:47.96" resultid="1573" heatid="2012" lane="3" entrytime="00:00:52.20" entrycourse="SCM" />
                <RESULT eventid="1113" points="125" swimtime="00:01:29.58" resultid="1574" heatid="2028" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="60" swimtime="00:00:55.40" resultid="1575" heatid="2068" lane="1" />
                <RESULT eventid="1293" points="128" swimtime="00:00:39.91" resultid="1576" heatid="2096" lane="4" entrytime="00:00:47.16" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Faisal" lastname="Basem Ghotme" birthdate="2010-12-18" gender="M" nation="BRA" license="390809" swrid="5596871" athleteid="1509" externalid="390809" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1096" points="452" swimtime="00:00:58.39" resultid="1510" heatid="2020" lane="4" entrytime="00:01:01.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="261" swimtime="00:01:14.74" resultid="1511" heatid="2049" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="359" swimtime="00:01:08.00" resultid="1512" heatid="2089" lane="3" entrytime="00:01:08.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="449" swimtime="00:00:26.32" resultid="1513" heatid="2110" lane="6" entrytime="00:00:26.52" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paula" lastname="Palma Fornarolli" birthdate="2013-08-07" gender="F" nation="BRA" license="411995" swrid="5740016" athleteid="1588" externalid="411995">
              <RESULTS>
                <RESULT eventid="1104" points="199" swimtime="00:03:08.89" resultid="1589" heatid="2023" lane="2" entrytime="00:03:33.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:27.40" />
                    <SPLIT distance="150" swimtime="00:02:20.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="202" swimtime="00:00:43.03" resultid="1590" heatid="2039" lane="4" entrytime="00:00:45.94" entrycourse="SCM" />
                <RESULT eventid="1264" status="DSQ" swimtime="00:01:43.67" resultid="1591" heatid="2084" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="226" swimtime="00:00:37.64" resultid="1592" heatid="2099" lane="5" entrytime="00:00:37.69" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marlon" lastname="Antonio Junior" birthdate="2013-05-12" gender="M" nation="BRA" license="397300" swrid="5641751" athleteid="1514" externalid="397300" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1107" status="DNS" swimtime="00:00:00.00" resultid="1515" heatid="2025" lane="1" entrytime="00:03:11.82" entrycourse="SCM" />
                <RESULT eventid="1151" status="DNS" swimtime="00:00:00.00" resultid="1516" heatid="2042" lane="4" entrytime="00:00:44.24" entrycourse="SCM" />
                <RESULT eventid="1267" status="DNS" swimtime="00:00:00.00" resultid="1517" heatid="2085" lane="1" />
                <RESULT eventid="1299" status="DNS" swimtime="00:00:00.00" resultid="1518" heatid="2102" lane="1" entrytime="00:00:35.46" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Mattiello" birthdate="2009-04-11" gender="F" nation="BRA" license="367011" swrid="5596914" athleteid="1463" externalid="367011" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1088" points="409" swimtime="00:01:07.68" resultid="1464" heatid="2016" lane="6" entrytime="00:01:07.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="402" swimtime="00:00:31.05" resultid="1465" heatid="2105" lane="4" entrytime="00:00:30.48" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Gabriel Dreher" birthdate="2011-12-05" gender="M" nation="BRA" license="403148" swrid="5676302" athleteid="1539" externalid="403148" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1096" points="153" swimtime="00:01:23.68" resultid="1540" heatid="2018" lane="1" entrytime="00:01:21.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="149" swimtime="00:00:41.66" resultid="1541" heatid="2036" lane="3" entrytime="00:00:47.84" entrycourse="SCM" />
                <RESULT eventid="1184" points="130" swimtime="00:00:49.18" resultid="1542" heatid="2055" lane="4" entrytime="00:00:56.95" entrycourse="SCM" />
                <RESULT eventid="1200" points="198" swimtime="00:06:04.06" resultid="1543" heatid="2061" lane="5" entrytime="00:06:02.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                    <SPLIT distance="100" swimtime="00:01:25.78" />
                    <SPLIT distance="150" swimtime="00:02:09.89" />
                    <SPLIT distance="200" swimtime="00:02:55.88" />
                    <SPLIT distance="250" swimtime="00:03:44.62" />
                    <SPLIT distance="300" swimtime="00:04:31.28" />
                    <SPLIT distance="350" swimtime="00:05:18.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="140" swimtime="00:01:33.07" resultid="1544" heatid="2088" lane="3" entrytime="00:01:28.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Rogge" birthdate="2008-09-02" gender="M" nation="BRA" license="383387" swrid="4883279" athleteid="1441" externalid="383387" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1096" points="481" swimtime="00:00:57.22" resultid="1442" heatid="2022" lane="1" entrytime="00:00:56.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="484" swimtime="00:00:25.67" resultid="1443" heatid="2110" lane="5" entrytime="00:00:25.81" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="De Assis Santos" birthdate="2003-02-21" gender="M" nation="BRA" license="342496" swrid="5596885" athleteid="1448" externalid="342496" level="INTERNE/IT">
              <RESULTS>
                <RESULT eventid="1068" points="415" swimtime="00:02:26.95" resultid="1449" heatid="2005" lane="6" entrytime="00:02:32.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                    <SPLIT distance="100" swimtime="00:01:05.12" />
                    <SPLIT distance="150" swimtime="00:01:51.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="435" swimtime="00:00:29.17" resultid="1450" heatid="2035" lane="2" />
                <RESULT eventid="1252" points="431" swimtime="00:00:28.78" resultid="1451" heatid="2079" lane="2" />
                <RESULT eventid="1278" points="440" swimtime="00:01:03.50" resultid="1452" heatid="2090" lane="4" entrytime="00:01:02.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Leticia Sbardelatti" birthdate="2011-07-28" gender="F" nation="BRA" license="403147" swrid="5676303" athleteid="1534" externalid="403147" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1088" points="245" swimtime="00:01:20.26" resultid="1535" heatid="2014" lane="6" entrytime="00:01:22.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="229" swimtime="00:00:46.32" resultid="1536" heatid="2053" lane="6" entrytime="00:00:49.97" entrycourse="SCM" />
                <RESULT eventid="1192" points="215" swimtime="00:06:25.94" resultid="1537" heatid="2058" lane="1" entrytime="00:06:15.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                    <SPLIT distance="100" swimtime="00:01:33.66" />
                    <SPLIT distance="150" swimtime="00:02:22.28" />
                    <SPLIT distance="200" swimtime="00:03:11.94" />
                    <SPLIT distance="250" swimtime="00:04:02.08" />
                    <SPLIT distance="300" swimtime="00:04:51.79" />
                    <SPLIT distance="350" swimtime="00:05:41.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="276" swimtime="00:00:35.18" resultid="1538" heatid="2104" lane="5" entrytime="00:00:35.73" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jeronimo" lastname="Pujato Flores" birthdate="2013-12-28" gender="M" nation="BRA" license="392839" swrid="5652625" athleteid="1555" externalid="392839" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1107" points="101" swimtime="00:03:33.18" resultid="1556" heatid="2024" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.20" />
                    <SPLIT distance="100" swimtime="00:01:42.69" />
                    <SPLIT distance="150" swimtime="00:02:38.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="93" swimtime="00:00:48.64" resultid="1557" heatid="2041" lane="4" entrytime="00:00:52.42" entrycourse="SCM" />
                <RESULT eventid="1299" points="103" swimtime="00:00:42.90" resultid="1558" heatid="2101" lane="5" entrytime="00:00:42.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ysadora" lastname="Bertoldo" birthdate="2010-04-09" gender="F" nation="BRA" license="376444" swrid="5588553" athleteid="1475" externalid="376444" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1116" points="420" swimtime="00:20:12.44" resultid="1476" heatid="2030" lane="3" entrytime="00:19:50.99" entrycourse="SCM" />
                <RESULT eventid="1192" points="432" swimtime="00:05:05.93" resultid="1477" heatid="2060" lane="1" entrytime="00:05:01.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="100" swimtime="00:01:14.14" />
                    <SPLIT distance="150" swimtime="00:01:53.46" />
                    <SPLIT distance="200" swimtime="00:02:32.56" />
                    <SPLIT distance="250" swimtime="00:03:12.01" />
                    <SPLIT distance="300" swimtime="00:03:50.49" />
                    <SPLIT distance="350" swimtime="00:04:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1244" points="332" swimtime="00:00:35.18" resultid="1478" heatid="2077" lane="3" entrytime="00:00:38.35" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrieli" lastname="Brietzke Sbardelatti" birthdate="2014-07-14" gender="F" nation="BRA" license="400456" swrid="4379861" athleteid="1519" externalid="400456" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1110" points="205" swimtime="00:01:25.11" resultid="1520" heatid="2027" lane="5" entrytime="00:01:39.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1154" points="163" swimtime="00:00:46.22" resultid="1521" heatid="2044" lane="1" entrytime="00:00:53.84" entrycourse="SCM" />
                <RESULT eventid="1212" points="155" swimtime="00:00:45.37" resultid="1522" heatid="2065" lane="3" entrytime="00:00:55.83" entrycourse="SCM" />
                <RESULT eventid="1290" points="167" swimtime="00:00:41.61" resultid="1523" heatid="2094" lane="6" entrytime="00:00:42.59" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Marques Petry" birthdate="2008-01-08" gender="M" nation="BRA" license="392351" swrid="4711489" athleteid="1466" externalid="392351" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1124" points="404" swimtime="00:19:05.50" resultid="1467" heatid="2031" lane="2" entrytime="00:19:25.84" entrycourse="SCM" />
                <RESULT eventid="1200" points="423" swimtime="00:04:42.67" resultid="1468" heatid="2062" lane="5" entrytime="00:05:00.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                    <SPLIT distance="100" swimtime="00:01:06.68" />
                    <SPLIT distance="150" swimtime="00:01:42.15" />
                    <SPLIT distance="200" swimtime="00:02:18.58" />
                    <SPLIT distance="250" swimtime="00:02:55.52" />
                    <SPLIT distance="300" swimtime="00:03:31.81" />
                    <SPLIT distance="350" swimtime="00:04:07.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1278" points="197" swimtime="00:01:22.96" resultid="1469" heatid="2089" lane="6" entrytime="00:01:22.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Axel" lastname="Ariel Giménez González" birthdate="2011-06-01" gender="M" nation="BRA" license="365755" swrid="5676299" athleteid="1545" externalid="365755" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1096" points="342" swimtime="00:01:04.06" resultid="1546" heatid="2020" lane="1" entrytime="00:01:04.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="268" swimtime="00:00:38.67" resultid="1547" heatid="2056" lane="1" entrytime="00:00:39.21" entrycourse="SCM" />
                <RESULT eventid="1236" status="DSQ" swimtime="00:01:23.83" resultid="1548" heatid="2074" lane="2" entrytime="00:01:32.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="335" swimtime="00:00:29.00" resultid="1549" heatid="2109" lane="6" entrytime="00:00:29.16" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
