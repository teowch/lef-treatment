<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.79911">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Guarapuava" name="63º Jogos Universitários do Paraná 2024" course="SCM" entrytype="INVITATION" hostclub="Prefeitura Municipal de Guarapuava" hostclub.url="https://guarapuava.pr.gov.br/" number="38310" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/newInterface/eventos/38310" startmethod="1" timing="AUTOMATIC" touchpad="ONESIDE" masters="F" withdrawuntil="2024-06-28" state="PR" nation="BRA">
      <AGEDATE value="2024-07-06" type="YEAR" />
      <POOL name="AquaCentro" lanemin="1" lanemax="5" />
      <FACILITY city="Guarapuava" name="AquaCentro" nation="BRA" state="PR" street="Rua Barão de Capanema, 788" street2="Santa Cruz" zip="85015-420" />
      <POINTTABLE pointtableid="3124" name="FINA Master Point Scoring" version="2024" />
      <QUALIFY from="2023-07-06" until="2024-07-05" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99233-1025" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99233-1025" street="Avenida do Batel, 1230" street2="Batel" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-07-06" daytime="15:30" endtime="18:49" number="1" officialmeeting="15:00" warmupfrom="14:30" warmupuntil="15:20">
          <EVENTS>
            <EVENT eventid="1074" daytime="15:30" gender="M" number="2" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2111" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1837" />
                    <RANKING order="2" place="2" resultid="1798" />
                    <RANKING order="3" place="3" resultid="1617" />
                    <RANKING order="4" place="4" resultid="1535" />
                    <RANKING order="5" place="5" resultid="1727" />
                    <RANKING order="6" place="6" resultid="1574" />
                    <RANKING order="7" place="7" resultid="1983" />
                    <RANKING order="8" place="-1" resultid="1904" />
                    <RANKING order="9" place="-1" resultid="1689" />
                    <RANKING order="10" place="-1" resultid="1612" />
                    <RANKING order="11" place="-1" resultid="1709" />
                    <RANKING order="12" place="-1" resultid="1927" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2153" daytime="15:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2154" daytime="15:34" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2155" daytime="15:38" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1087" daytime="15:42" gender="F" number="3" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2112" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1538" />
                    <RANKING order="2" place="2" resultid="1909" />
                    <RANKING order="3" place="3" resultid="1804" />
                    <RANKING order="4" place="-1" resultid="1832" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2156" daytime="15:42" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1100" daytime="15:46" gender="M" number="4" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2114" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1883" />
                    <RANKING order="2" place="2" resultid="1841" />
                    <RANKING order="3" place="3" resultid="1872" />
                    <RANKING order="4" place="4" resultid="1922" />
                    <RANKING order="5" place="5" resultid="2238" />
                    <RANKING order="6" place="6" resultid="1675" />
                    <RANKING order="7" place="7" resultid="1671" />
                    <RANKING order="8" place="8" resultid="1950" />
                    <RANKING order="9" place="9" resultid="1781" />
                    <RANKING order="10" place="10" resultid="1734" />
                    <RANKING order="11" place="11" resultid="1700" />
                    <RANKING order="12" place="-1" resultid="1613" />
                    <RANKING order="13" place="-1" resultid="1590" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2157" daytime="15:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2158" daytime="15:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2159" daytime="15:52" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1113" daytime="15:54" gender="F" number="5" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2115" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1570" />
                    <RANKING order="2" place="2" resultid="1856" />
                    <RANKING order="3" place="3" resultid="1808" />
                    <RANKING order="4" place="4" resultid="1978" />
                    <RANKING order="5" place="5" resultid="1623" />
                    <RANKING order="6" place="6" resultid="1940" />
                    <RANKING order="7" place="7" resultid="1602" />
                    <RANKING order="8" place="8" resultid="1635" />
                    <RANKING order="9" place="9" resultid="1594" />
                    <RANKING order="10" place="10" resultid="1632" />
                    <RANKING order="11" place="11" resultid="1775" />
                    <RANKING order="12" place="-1" resultid="1767" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2160" daytime="15:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2161" daytime="15:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2162" daytime="15:58" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1126" daytime="16:14" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2116" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1934" />
                    <RANKING order="2" place="2" resultid="1562" />
                    <RANKING order="3" place="3" resultid="1815" />
                    <RANKING order="4" place="4" resultid="1578" />
                    <RANKING order="5" place="5" resultid="1528" />
                    <RANKING order="6" place="6" resultid="1652" />
                    <RANKING order="7" place="7" resultid="1646" />
                    <RANKING order="8" place="8" resultid="1887" />
                    <RANKING order="9" place="9" resultid="1733" />
                    <RANKING order="10" place="10" resultid="1769" />
                    <RANKING order="11" place="11" resultid="1667" />
                    <RANKING order="12" place="12" resultid="1949" />
                    <RANKING order="13" place="13" resultid="1780" />
                    <RANKING order="14" place="14" resultid="1982" />
                    <RANKING order="15" place="-1" resultid="1790" />
                    <RANKING order="16" place="-1" resultid="1703" />
                    <RANKING order="17" place="-1" resultid="1714" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2163" daytime="16:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2164" daytime="16:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2165" daytime="16:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2166" daytime="16:20" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1139" daytime="16:24" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2117" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1908" />
                    <RANKING order="2" place="2" resultid="1661" />
                    <RANKING order="3" place="3" resultid="1860" />
                    <RANKING order="4" place="4" resultid="1803" />
                    <RANKING order="5" place="5" resultid="1586" />
                    <RANKING order="6" place="6" resultid="1598" />
                    <RANKING order="7" place="7" resultid="1977" />
                    <RANKING order="8" place="8" resultid="1971" />
                    <RANKING order="9" place="9" resultid="1738" />
                    <RANKING order="10" place="10" resultid="1939" />
                    <RANKING order="11" place="11" resultid="1774" />
                    <RANKING order="12" place="-1" resultid="1639" />
                    <RANKING order="13" place="-1" resultid="1766" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2167" daytime="16:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2168" daytime="16:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2169" daytime="16:28" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1152" daytime="16:30" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2118" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1797" />
                    <RANKING order="2" place="2" resultid="1876" />
                    <RANKING order="3" place="3" resultid="1534" />
                    <RANKING order="4" place="4" resultid="1656" />
                    <RANKING order="5" place="-1" resultid="1849" />
                    <RANKING order="6" place="-1" resultid="1921" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2170" daytime="16:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2171" daytime="16:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1165" daytime="16:40" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2119" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1891" />
                    <RANKING order="2" place="2" resultid="1743" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2172" daytime="16:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1178" daytime="16:44" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2120" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1550" />
                    <RANKING order="2" place="2" resultid="1554" />
                    <RANKING order="3" place="3" resultid="1852" />
                    <RANKING order="4" place="4" resultid="2148" />
                    <RANKING order="5" place="5" resultid="1846" />
                    <RANKING order="6" place="6" resultid="1755" />
                    <RANKING order="7" place="7" resultid="1618" />
                    <RANKING order="8" place="8" resultid="1529" />
                    <RANKING order="9" place="9" resultid="1935" />
                    <RANKING order="10" place="10" resultid="1728" />
                    <RANKING order="11" place="11" resultid="1647" />
                    <RANKING order="12" place="12" resultid="1984" />
                    <RANKING order="13" place="13" resultid="1644" />
                    <RANKING order="14" place="-1" resultid="1710" />
                    <RANKING order="15" place="-1" resultid="1717" />
                    <RANKING order="16" place="-1" resultid="1747" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2173" daytime="16:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2174" daytime="16:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2175" daytime="16:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2176" daytime="16:48" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1191" daytime="16:52" gender="F" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2121" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1809" />
                    <RANKING order="2" place="2" resultid="1761" />
                    <RANKING order="3" place="3" resultid="1805" />
                    <RANKING order="4" place="4" resultid="1861" />
                    <RANKING order="5" place="5" resultid="1739" />
                    <RANKING order="6" place="6" resultid="1558" />
                    <RANKING order="7" place="7" resultid="1972" />
                    <RANKING order="8" place="8" resultid="1599" />
                    <RANKING order="9" place="9" resultid="1776" />
                    <RANKING order="10" place="10" resultid="1633" />
                    <RANKING order="11" place="-1" resultid="1640" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2177" daytime="16:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2178" daytime="16:52" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1061" daytime="16:56" gender="F" number="1" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1073" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1819" />
                    <RANKING order="2" place="2" resultid="1662" />
                    <RANKING order="3" place="3" resultid="1827" />
                    <RANKING order="4" place="4" resultid="1965" />
                    <RANKING order="5" place="5" resultid="1960" />
                    <RANKING order="6" place="6" resultid="1546" />
                    <RANKING order="7" place="7" resultid="1744" />
                    <RANKING order="8" place="-1" resultid="1823" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2151" daytime="16:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2152" daytime="17:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1204" daytime="17:24" gender="M" number="12" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2123" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1518" />
                    <RANKING order="2" place="2" resultid="1796" />
                    <RANKING order="3" place="3" resultid="1871" />
                    <RANKING order="4" place="4" resultid="1542" />
                    <RANKING order="5" place="5" resultid="1954" />
                    <RANKING order="6" place="6" resultid="1566" />
                    <RANKING order="7" place="7" resultid="1866" />
                    <RANKING order="8" place="8" resultid="1685" />
                    <RANKING order="9" place="-1" resultid="1524" />
                    <RANKING order="10" place="-1" resultid="1920" />
                    <RANKING order="11" place="-1" resultid="1704" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2179" daytime="17:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2180" daytime="17:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2181" daytime="18:10" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1217" daytime="18:50" gender="F" number="13" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1218" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1912" />
                    <RANKING order="2" place="2" resultid="1604" />
                    <RANKING order="3" place="3" resultid="1985" />
                    <RANKING order="4" place="4" resultid="1783" />
                    <RANKING order="5" place="5" resultid="1692" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2182" daytime="18:50" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1219" daytime="18:56" gender="M" number="14" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1220" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1915" />
                    <RANKING order="2" place="2" resultid="1607" />
                    <RANKING order="3" place="3" resultid="1695" />
                    <RANKING order="4" place="4" resultid="1786" />
                    <RANKING order="5" place="5" resultid="1988" />
                    <RANKING order="6" place="-1" resultid="2245" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2183" daytime="18:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2184" daytime="19:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-07-07" daytime="09:00" endtime="11:42" number="2" officialmeeting="08:30" warmupfrom="08:00" warmupuntil="08:50">
          <EVENTS>
            <EVENT eventid="1221" daytime="09:00" gender="F" number="15" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2124" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1820" />
                    <RANKING order="2" place="2" resultid="1910" />
                    <RANKING order="3" place="3" resultid="1829" />
                    <RANKING order="4" place="4" resultid="1966" />
                    <RANKING order="5" place="5" resultid="1752" />
                    <RANKING order="6" place="6" resultid="1961" />
                    <RANKING order="7" place="7" resultid="1547" />
                    <RANKING order="8" place="8" resultid="1973" />
                    <RANKING order="9" place="9" resultid="1624" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2185" daytime="09:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2186" daytime="09:06" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1234" daytime="09:14" gender="M" number="16" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2125" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1543" />
                    <RANKING order="2" place="2" resultid="1955" />
                    <RANKING order="3" place="3" resultid="1888" />
                    <RANKING order="4" place="4" resultid="1575" />
                    <RANKING order="5" place="5" resultid="1677" />
                    <RANKING order="6" place="6" resultid="1658" />
                    <RANKING order="7" place="7" resultid="1567" />
                    <RANKING order="8" place="8" resultid="1867" />
                    <RANKING order="9" place="9" resultid="1686" />
                    <RANKING order="10" place="-1" resultid="1520" />
                    <RANKING order="11" place="-1" resultid="1525" />
                    <RANKING order="12" place="-1" resultid="1928" />
                    <RANKING order="13" place="-1" resultid="1931" />
                    <RANKING order="14" place="-1" resultid="1799" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2187" daytime="09:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2188" daytime="09:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2189" daytime="09:26" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1247" daytime="09:34" gender="F" number="17" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2126" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1810" />
                    <RANKING order="2" place="2" resultid="1762" />
                    <RANKING order="3" place="3" resultid="1862" />
                    <RANKING order="4" place="4" resultid="1893" />
                    <RANKING order="5" place="5" resultid="1559" />
                    <RANKING order="6" place="-1" resultid="1777" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2190" daytime="09:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2191" daytime="09:38" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1260" daytime="09:44" gender="M" number="18" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2127" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2150" />
                    <RANKING order="2" place="2" resultid="1551" />
                    <RANKING order="3" place="3" resultid="1853" />
                    <RANKING order="4" place="4" resultid="1619" />
                    <RANKING order="5" place="5" resultid="1879" />
                    <RANKING order="6" place="6" resultid="1582" />
                    <RANKING order="7" place="7" resultid="1729" />
                    <RANKING order="8" place="8" resultid="1648" />
                    <RANKING order="9" place="9" resultid="1628" />
                    <RANKING order="10" place="-1" resultid="1711" />
                    <RANKING order="11" place="-1" resultid="1748" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2192" daytime="09:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2193" daytime="09:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2194" daytime="09:50" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1273" daytime="09:56" gender="F" number="19" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2128" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1911" />
                    <RANKING order="2" place="2" resultid="1663" />
                    <RANKING order="3" place="3" resultid="1539" />
                    <RANKING order="4" place="4" resultid="1857" />
                    <RANKING order="5" place="5" resultid="1763" />
                    <RANKING order="6" place="6" resultid="1588" />
                    <RANKING order="7" place="7" resultid="1979" />
                    <RANKING order="8" place="8" resultid="1863" />
                    <RANKING order="9" place="9" resultid="1967" />
                    <RANKING order="10" place="10" resultid="1740" />
                    <RANKING order="11" place="11" resultid="1962" />
                    <RANKING order="12" place="12" resultid="1595" />
                    <RANKING order="13" place="13" resultid="1636" />
                    <RANKING order="14" place="14" resultid="1778" />
                    <RANKING order="15" place="-1" resultid="1941" />
                    <RANKING order="16" place="-1" resultid="1641" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2195" daytime="09:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2196" daytime="09:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2197" daytime="09:58" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1286" daytime="10:00" gender="M" number="20" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2129" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1555" />
                    <RANKING order="2" place="2" resultid="1936" />
                    <RANKING order="3" place="3" resultid="1906" />
                    <RANKING order="4" place="4" resultid="1816" />
                    <RANKING order="5" place="5" resultid="1946" />
                    <RANKING order="6" place="6" resultid="1579" />
                    <RANKING order="7" place="7" resultid="1530" />
                    <RANKING order="8" place="8" resultid="1756" />
                    <RANKING order="9" place="9" resultid="1956" />
                    <RANKING order="10" place="10" resultid="1880" />
                    <RANKING order="11" place="11" resultid="1771" />
                    <RANKING order="12" place="12" resultid="1668" />
                    <RANKING order="13" place="13" resultid="1951" />
                    <RANKING order="14" place="14" resultid="1735" />
                    <RANKING order="15" place="15" resultid="1681" />
                    <RANKING order="16" place="16" resultid="1629" />
                    <RANKING order="17" place="-1" resultid="1706" />
                    <RANKING order="18" place="-1" resultid="1715" />
                    <RANKING order="19" place="-1" resultid="1721" />
                    <RANKING order="20" place="-1" resultid="1792" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2198" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2199" daytime="10:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2200" daytime="10:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2201" daytime="10:06" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1299" daytime="10:22" gender="F" number="21" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2130" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1751" />
                    <RANKING order="2" place="2" resultid="1828" />
                    <RANKING order="3" place="3" resultid="1600" />
                    <RANKING order="4" place="-1" resultid="1833" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2202" daytime="10:22" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1312" daytime="10:26" gender="M" number="22" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2131" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1884" />
                    <RANKING order="2" place="2" resultid="1842" />
                    <RANKING order="3" place="3" resultid="1873" />
                    <RANKING order="4" place="4" resultid="1676" />
                    <RANKING order="5" place="5" resultid="1672" />
                    <RANKING order="6" place="-1" resultid="1519" />
                    <RANKING order="7" place="-1" resultid="1614" />
                    <RANKING order="8" place="-1" resultid="1705" />
                    <RANKING order="9" place="-1" resultid="1923" />
                    <RANKING order="10" place="-1" resultid="1591" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2203" daytime="10:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2204" daytime="10:30" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1325" daytime="10:34" gender="F" number="23" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2132" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1892" />
                    <RANKING order="2" place="2" resultid="1587" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2205" daytime="10:34" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1338" daytime="10:38" gender="M" number="24" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2136" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1838" />
                    <RANKING order="2" place="2" resultid="1905" />
                    <RANKING order="3" place="3" resultid="1877" />
                    <RANKING order="4" place="4" resultid="1563" />
                    <RANKING order="5" place="5" resultid="1536" />
                    <RANKING order="6" place="6" resultid="1770" />
                    <RANKING order="7" place="7" resultid="1657" />
                    <RANKING order="8" place="8" resultid="1653" />
                    <RANKING order="9" place="9" resultid="1690" />
                    <RANKING order="10" place="-1" resultid="1791" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2206" daytime="10:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2207" daytime="10:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1351" daytime="10:42" gender="F" number="25" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2135" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1811" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2208" daytime="10:42" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1364" daytime="10:50" gender="M" number="26" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2134" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1800" />
                    <RANKING order="2" place="2" resultid="1843" />
                    <RANKING order="3" place="3" resultid="1945" />
                    <RANKING order="4" place="4" resultid="1620" />
                    <RANKING order="5" place="5" resultid="1924" />
                    <RANKING order="6" place="6" resultid="1868" />
                    <RANKING order="7" place="-1" resultid="1615" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2209" daytime="10:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2210" daytime="10:56" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1377" daytime="11:20" gender="F" number="27" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1378" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1913" />
                    <RANKING order="2" place="2" resultid="1605" />
                    <RANKING order="3" place="3" resultid="1986" />
                    <RANKING order="4" place="4" resultid="1784" />
                    <RANKING order="5" place="-1" resultid="1693" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2211" daytime="11:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1379" daytime="11:30" gender="M" number="28" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1380" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1916" />
                    <RANKING order="2" place="2" resultid="1608" />
                    <RANKING order="3" place="3" resultid="1696" />
                    <RANKING order="4" place="4" resultid="1989" />
                    <RANKING order="5" place="-1" resultid="1723" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2212" daytime="11:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-07-07" daytime="15:30" endtime="17:49" number="3" officialmeeting="15:00" warmupfrom="14:30" warmupuntil="15:20">
          <EVENTS>
            <EVENT eventid="1381" daytime="15:30" gender="M" number="29" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2147" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1544" />
                    <RANKING order="2" place="2" resultid="1958" />
                    <RANKING order="3" place="3" resultid="1679" />
                    <RANKING order="4" place="4" resultid="1568" />
                    <RANKING order="5" place="5" resultid="1869" />
                    <RANKING order="6" place="6" resultid="1687" />
                    <RANKING order="7" place="-1" resultid="1521" />
                    <RANKING order="8" place="-1" resultid="1526" />
                    <RANKING order="9" place="-1" resultid="1707" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2213" daytime="15:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2214" daytime="15:42" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1394" daytime="15:56" gender="F" number="30" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2146" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1571" />
                    <RANKING order="2" place="2" resultid="1664" />
                    <RANKING order="3" place="3" resultid="1753" />
                    <RANKING order="4" place="4" resultid="1812" />
                    <RANKING order="5" place="5" resultid="1548" />
                    <RANKING order="6" place="6" resultid="1625" />
                    <RANKING order="7" place="7" resultid="1637" />
                    <RANKING order="8" place="8" resultid="1596" />
                    <RANKING order="9" place="-1" resultid="1942" />
                    <RANKING order="10" place="-1" resultid="1834" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2215" daytime="15:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2216" daytime="15:58" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1407" daytime="16:02" gender="M" number="31" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2144" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1885" />
                    <RANKING order="2" place="2" resultid="1844" />
                    <RANKING order="3" place="3" resultid="1874" />
                    <RANKING order="4" place="4" resultid="1678" />
                    <RANKING order="5" place="5" resultid="1673" />
                    <RANKING order="6" place="6" resultid="1782" />
                    <RANKING order="7" place="7" resultid="1682" />
                    <RANKING order="8" place="-1" resultid="1701" />
                    <RANKING order="9" place="-1" resultid="1592" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2217" daytime="16:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2218" daytime="16:04" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1420" daytime="16:08" gender="F" number="32" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2143" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1665" />
                    <RANKING order="2" place="2" resultid="1806" />
                    <RANKING order="3" place="3" resultid="1969" />
                    <RANKING order="4" place="4" resultid="1980" />
                    <RANKING order="5" place="5" resultid="1975" />
                    <RANKING order="6" place="-1" resultid="1825" />
                    <RANKING order="7" place="-1" resultid="1835" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2219" daytime="16:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2220" daytime="16:12" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1433" daytime="16:16" gender="M" number="33" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2142" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1817" />
                    <RANKING order="2" place="2" resultid="1564" />
                    <RANKING order="3" place="3" resultid="1947" />
                    <RANKING order="4" place="4" resultid="1957" />
                    <RANKING order="5" place="5" resultid="1584" />
                    <RANKING order="6" place="6" resultid="1889" />
                    <RANKING order="7" place="7" resultid="1576" />
                    <RANKING order="8" place="8" resultid="1731" />
                    <RANKING order="9" place="9" resultid="1650" />
                    <RANKING order="10" place="10" resultid="1669" />
                    <RANKING order="11" place="11" resultid="1630" />
                    <RANKING order="12" place="-1" resultid="1850" />
                    <RANKING order="13" place="-1" resultid="1929" />
                    <RANKING order="14" place="-1" resultid="1932" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2221" daytime="16:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2222" daytime="16:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2223" daytime="16:24" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1446" daytime="16:42" gender="F" number="34" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2141" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1572" />
                    <RANKING order="2" place="2" resultid="1858" />
                    <RANKING order="3" place="3" resultid="1896" />
                    <RANKING order="4" place="4" resultid="1626" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2224" daytime="16:42" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1459" daytime="16:44" gender="M" number="35" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2140" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1556" />
                    <RANKING order="2" place="2" resultid="1839" />
                    <RANKING order="3" place="3" resultid="1847" />
                    <RANKING order="4" place="4" resultid="1531" />
                    <RANKING order="5" place="5" resultid="1772" />
                    <RANKING order="6" place="6" resultid="1654" />
                    <RANKING order="7" place="7" resultid="1580" />
                    <RANKING order="8" place="8" resultid="1659" />
                    <RANKING order="9" place="9" resultid="1736" />
                    <RANKING order="10" place="10" resultid="1952" />
                    <RANKING order="11" place="11" resultid="1691" />
                    <RANKING order="12" place="-1" resultid="1759" />
                    <RANKING order="13" place="-1" resultid="1719" />
                    <RANKING order="14" place="-1" resultid="1793" />
                    <RANKING order="15" place="-1" resultid="1937" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2225" daytime="16:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2226" daytime="16:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2227" daytime="16:48" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1472" daytime="16:50" gender="F" number="36" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2139" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1540" />
                    <RANKING order="2" place="2" resultid="1764" />
                    <RANKING order="3" place="3" resultid="1864" />
                    <RANKING order="4" place="4" resultid="1895" />
                    <RANKING order="5" place="5" resultid="1560" />
                    <RANKING order="6" place="6" resultid="1974" />
                    <RANKING order="7" place="7" resultid="1741" />
                    <RANKING order="8" place="-1" resultid="1642" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2228" daytime="16:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2229" daytime="16:52" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1485" daytime="16:56" gender="M" number="37" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2138" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1552" />
                    <RANKING order="2" place="2" resultid="1854" />
                    <RANKING order="3" place="3" resultid="2149" />
                    <RANKING order="4" place="4" resultid="1757" />
                    <RANKING order="5" place="5" resultid="1621" />
                    <RANKING order="6" place="6" resultid="1881" />
                    <RANKING order="7" place="7" resultid="1583" />
                    <RANKING order="8" place="8" resultid="1730" />
                    <RANKING order="9" place="9" resultid="1649" />
                    <RANKING order="10" place="10" resultid="1683" />
                    <RANKING order="11" place="-1" resultid="1712" />
                    <RANKING order="12" place="-1" resultid="1718" />
                    <RANKING order="13" place="-1" resultid="1749" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2230" daytime="16:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2231" daytime="16:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2232" daytime="17:00" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1498" daytime="17:04" gender="F" number="38" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2137" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1821" />
                    <RANKING order="2" place="2" resultid="1968" />
                    <RANKING order="3" place="3" resultid="1963" />
                    <RANKING order="4" place="4" resultid="1745" />
                    <RANKING order="5" place="5" resultid="1603" />
                    <RANKING order="6" place="-1" resultid="1824" />
                    <RANKING order="7" place="-1" resultid="1830" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2233" daytime="17:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2234" daytime="17:32" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1511" daytime="18:12" gender="M" number="39" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1512" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1917" />
                    <RANKING order="2" place="2" resultid="1609" />
                    <RANKING order="3" place="3" resultid="1697" />
                    <RANKING order="4" place="4" resultid="1787" />
                    <RANKING order="5" place="5" resultid="1990" />
                    <RANKING order="6" place="-1" resultid="1724" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2235" daytime="18:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2236" daytime="18:16" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1513" daytime="18:22" gender="F" number="40" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1514" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1914" />
                    <RANKING order="2" place="2" resultid="1606" />
                    <RANKING order="3" place="3" resultid="1785" />
                    <RANKING order="4" place="4" resultid="1987" />
                    <RANKING order="5" place="5" resultid="1694" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2237" daytime="18:22" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="13521" nation="BRA" region="PR" clubid="1788" name="Unicentro (Guarapuava)" shortname="Unicentro(Guarapuava">
          <ATHLETES>
            <ATHLETE firstname="William" lastname="Dos Lopes" birthdate="2005-12-23" gender="M" nation="BRA" license="V413313" athleteid="1789" externalid="V413313">
              <RESULTS>
                <RESULT eventid="1126" status="DSQ" swimtime="00:01:35.04" resultid="1790" heatid="2164" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" status="DNS" swimtime="00:00:00.00" resultid="1791" heatid="2206" lane="4" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="1792" heatid="2198" lane="1" />
                <RESULT eventid="1459" status="DNS" swimtime="00:00:00.00" resultid="1793" heatid="2225" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="9760" nation="BRA" region="PR" clubid="1522" name="Integrado (Campo Mourão)" shortname="Integrado (Campo M.)">
          <ATHLETES>
            <ATHLETE firstname="Henrique" lastname="Pedroso Silverio" birthdate="1994-11-21" gender="M" nation="BRA" license="115715" swrid="5603892" athleteid="1523" externalid="115715">
              <RESULTS>
                <RESULT eventid="1204" status="DNS" swimtime="00:00:00.00" resultid="1524" heatid="2181" lane="5" entrytime="00:20:45.97" entrycourse="SCM" />
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="1525" heatid="2189" lane="2" entrytime="00:05:00.79" entrycourse="SCM" />
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="1526" heatid="2213" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Franco Santos" birthdate="2002-01-03" gender="M" nation="BRA" license="290441" swrid="5546064" athleteid="1527" externalid="290441">
              <RESULTS>
                <RESULT eventid="1126" points="489" swimtime="00:01:00.18" resultid="1528" heatid="2166" lane="2" entrytime="00:00:56.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="529" swimtime="00:00:33.37" resultid="1529" heatid="2175" lane="5" />
                <RESULT eventid="1286" points="529" swimtime="00:00:26.31" resultid="1530" heatid="2201" lane="1" entrytime="00:00:25.66" entrycourse="SCM" />
                <RESULT eventid="1459" points="552" swimtime="00:00:28.22" resultid="1531" heatid="2227" lane="5" entrytime="00:00:27.76" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="12426" nation="BRA" region="PR" clubid="1698" name="Uepg (Ponta Grossa)">
          <ATHLETES>
            <ATHLETE firstname="Guinter" lastname="Sponholz Neiverth" birthdate="2003-02-18" gender="M" nation="BRA" license="V348329" athleteid="1716" externalid="V348329">
              <RESULTS>
                <RESULT eventid="1178" status="DNS" swimtime="00:00:00.00" resultid="1717" heatid="2173" lane="3" />
                <RESULT eventid="1485" status="DNS" swimtime="00:00:00.00" resultid="1718" heatid="2231" lane="1" />
                <RESULT eventid="1459" status="DNS" swimtime="00:00:00.00" resultid="1719" heatid="2226" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Mandalozzo Tebcherani" birthdate="2006-03-02" gender="M" nation="BRA" license="295181" swrid="5622289" athleteid="1713" externalid="295181">
              <RESULTS>
                <RESULT eventid="1126" status="DNS" swimtime="00:00:00.00" resultid="1714" heatid="2165" lane="2" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="1715" heatid="2198" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Gueiber" birthdate="2000-05-22" gender="M" nation="BRA" license="V121351" athleteid="1702" externalid="V121351">
              <RESULTS>
                <RESULT eventid="1126" status="DNS" swimtime="00:00:00.00" resultid="1703" heatid="2164" lane="5" />
                <RESULT eventid="1204" status="WDR" swimtime="00:00:00.00" resultid="1704" heatid="2179" lane="3" entrytime="00:20:57.58" entrycourse="SCM" />
                <RESULT eventid="1312" status="DNS" swimtime="00:00:00.00" resultid="1705" heatid="2203" lane="3" entrytime="00:02:33.62" entrycourse="SCM" />
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="1706" heatid="2201" lane="5" entrytime="00:00:25.45" entrycourse="SCM" />
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="1707" heatid="2214" lane="2" entrytime="00:10:27.98" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Carlos Cherubim" birthdate="2003-03-31" gender="M" nation="BRA" license="V295223" athleteid="1699" externalid="V295223">
              <RESULTS>
                <RESULT eventid="1100" points="198" swimtime="00:00:40.65" resultid="1700" heatid="2159" lane="5" entrytime="00:00:31.74" entrycourse="SCM" />
                <RESULT eventid="1407" status="DNS" swimtime="00:00:00.00" resultid="1701" heatid="2218" lane="5" entrytime="00:01:12.35" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Tonon" birthdate="2003-12-11" gender="M" nation="BRA" license="V387228" athleteid="1720" externalid="V387228">
              <RESULTS>
                <RESULT eventid="1286" status="DNS" swimtime="00:00:00.00" resultid="1721" heatid="2199" lane="3" entrytime="00:00:29.51" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Renato" lastname="Mandalozzo Tebcherani" birthdate="2004-03-16" gender="M" nation="BRA" license="279221" swrid="5622290" athleteid="1708" externalid="279221">
              <RESULTS>
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="1709" heatid="2155" lane="5" entrytime="00:02:32.40" entrycourse="SCM" />
                <RESULT eventid="1178" status="DNS" swimtime="00:00:00.00" resultid="1710" heatid="2174" lane="4" />
                <RESULT eventid="1260" status="DNS" swimtime="00:00:00.00" resultid="1711" heatid="2194" lane="2" entrytime="00:02:44.81" entrycourse="SCM" />
                <RESULT eventid="1485" status="DNS" swimtime="00:00:00.00" resultid="1712" heatid="2232" lane="2" entrytime="00:01:13.22" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M">
              <RESULTS>
                <RESULT eventid="1219" status="WDR" swimtime="00:00:00.00" resultid="2245" heatid="2183" lane="3" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="UEPG (PONTA GROSSA) &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1379" status="WDR" swimtime="00:00:00.00" resultid="1723" heatid="2212" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="2" reactiontime="0" />
                    <RELAYPOSITION number="3" reactiontime="0" />
                    <RELAYPOSITION number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" status="WDR" swimtime="00:00:00.00" resultid="1724" heatid="2235" lane="3" />
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="18694" nation="BRA" region="PR" clubid="1918" name="Uniguairaca (Guarapuava)" shortname="Uniguairaca (Guarapu">
          <ATHLETES>
            <ATHLETE firstname="Kevin" lastname="Roberto Carvalho" birthdate="2001-06-26" gender="M" nation="BRA" license="V374674" athleteid="1919" externalid="V374674">
              <RESULTS>
                <RESULT eventid="1204" status="DNS" swimtime="00:00:00.00" resultid="1920" heatid="2180" lane="5" />
                <RESULT eventid="1152" status="DNS" swimtime="00:00:00.00" resultid="1921" heatid="2170" lane="2" />
                <RESULT eventid="1100" points="507" swimtime="00:00:29.72" resultid="1922" heatid="2157" lane="4" />
                <RESULT eventid="1312" status="DNS" swimtime="00:00:00.00" resultid="1923" heatid="2203" lane="5" />
                <RESULT eventid="1364" points="246" swimtime="00:06:46.07" resultid="1924" heatid="2209" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                    <SPLIT distance="100" swimtime="00:01:14.19" />
                    <SPLIT distance="150" swimtime="00:02:02.62" />
                    <SPLIT distance="200" swimtime="00:02:52.43" />
                    <SPLIT distance="250" swimtime="00:03:48.39" />
                    <SPLIT distance="300" swimtime="00:04:47.09" />
                    <SPLIT distance="350" swimtime="00:05:46.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4007" nation="BRA" region="PR" clubid="1794" name="Unicesumar (Maringá)">
          <ATHLETES>
            <ATHLETE firstname="Francisco" lastname="Augusto Chiquetti" birthdate="2002-10-28" gender="M" nation="BRA" license="V318499" athleteid="1865" externalid="V318499">
              <RESULTS>
                <RESULT eventid="1204" points="206" swimtime="00:26:12.40" resultid="1866" heatid="2180" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                    <SPLIT distance="100" swimtime="00:01:21.67" />
                    <SPLIT distance="150" swimtime="00:02:05.94" />
                    <SPLIT distance="200" swimtime="00:02:53.22" />
                    <SPLIT distance="250" swimtime="00:03:42.82" />
                    <SPLIT distance="300" swimtime="00:04:33.31" />
                    <SPLIT distance="350" swimtime="00:05:26.25" />
                    <SPLIT distance="400" swimtime="00:06:19.03" />
                    <SPLIT distance="450" swimtime="00:07:15.27" />
                    <SPLIT distance="500" swimtime="00:08:08.59" />
                    <SPLIT distance="550" swimtime="00:09:02.01" />
                    <SPLIT distance="600" swimtime="00:09:56.59" />
                    <SPLIT distance="650" swimtime="00:10:51.01" />
                    <SPLIT distance="700" swimtime="00:11:46.96" />
                    <SPLIT distance="750" swimtime="00:12:41.94" />
                    <SPLIT distance="800" swimtime="00:13:36.32" />
                    <SPLIT distance="850" swimtime="00:14:30.79" />
                    <SPLIT distance="900" swimtime="00:15:26.82" />
                    <SPLIT distance="950" swimtime="00:16:21.35" />
                    <SPLIT distance="1000" swimtime="00:17:16.70" />
                    <SPLIT distance="1050" swimtime="00:18:10.76" />
                    <SPLIT distance="1100" swimtime="00:19:05.05" />
                    <SPLIT distance="1150" swimtime="00:20:00.78" />
                    <SPLIT distance="1200" swimtime="00:20:56.82" />
                    <SPLIT distance="1250" swimtime="00:21:51.66" />
                    <SPLIT distance="1300" swimtime="00:22:46.52" />
                    <SPLIT distance="1350" swimtime="00:23:39.67" />
                    <SPLIT distance="1400" swimtime="00:24:30.40" />
                    <SPLIT distance="1450" swimtime="00:25:23.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="254" swimtime="00:06:07.62" resultid="1867" heatid="2188" lane="4" entrytime="00:05:31.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                    <SPLIT distance="150" swimtime="00:01:55.28" />
                    <SPLIT distance="200" swimtime="00:02:43.13" />
                    <SPLIT distance="250" swimtime="00:03:34.70" />
                    <SPLIT distance="300" swimtime="00:04:27.11" />
                    <SPLIT distance="350" swimtime="00:05:17.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1364" points="213" swimtime="00:07:06.14" resultid="1868" heatid="2210" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                    <SPLIT distance="100" swimtime="00:01:21.87" />
                    <SPLIT distance="150" swimtime="00:02:21.43" />
                    <SPLIT distance="200" swimtime="00:03:23.07" />
                    <SPLIT distance="250" swimtime="00:04:24.19" />
                    <SPLIT distance="300" swimtime="00:05:27.94" />
                    <SPLIT distance="350" swimtime="00:06:18.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1381" points="224" swimtime="00:13:22.96" resultid="1869" heatid="2213" lane="3" entrytime="00:11:45.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:09.43" />
                    <SPLIT distance="200" swimtime="00:03:00.53" />
                    <SPLIT distance="250" swimtime="00:03:51.78" />
                    <SPLIT distance="300" swimtime="00:04:44.47" />
                    <SPLIT distance="350" swimtime="00:05:36.79" />
                    <SPLIT distance="400" swimtime="00:06:30.14" />
                    <SPLIT distance="450" swimtime="00:07:22.49" />
                    <SPLIT distance="500" swimtime="00:08:14.17" />
                    <SPLIT distance="550" swimtime="00:09:07.86" />
                    <SPLIT distance="600" swimtime="00:10:00.08" />
                    <SPLIT distance="650" swimtime="00:10:51.81" />
                    <SPLIT distance="700" swimtime="00:11:44.92" />
                    <SPLIT distance="750" swimtime="00:12:40.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carol" lastname="De Hertel" birthdate="2001-02-20" gender="F" nation="BRA" license="118424" swrid="5727648" athleteid="1822" externalid="118424">
              <RESULTS>
                <RESULT eventid="1061" status="WDR" swimtime="00:00:00.00" resultid="1823" />
                <RESULT eventid="1498" status="WDR" swimtime="00:00:00.00" resultid="1824" />
                <RESULT eventid="1420" status="WDR" swimtime="00:00:00.00" resultid="1825" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Paiz Ribeiro" birthdate="2006-02-17" gender="M" nation="BRA" license="297583" swrid="5596921" athleteid="1795" externalid="297583">
              <RESULTS>
                <RESULT eventid="1204" points="578" swimtime="00:18:35.64" resultid="1796" heatid="2180" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:09.33" />
                    <SPLIT distance="150" swimtime="00:01:46.39" />
                    <SPLIT distance="200" swimtime="00:02:23.32" />
                    <SPLIT distance="250" swimtime="00:02:59.53" />
                    <SPLIT distance="300" swimtime="00:03:36.41" />
                    <SPLIT distance="350" swimtime="00:04:13.21" />
                    <SPLIT distance="400" swimtime="00:04:49.86" />
                    <SPLIT distance="450" swimtime="00:05:26.97" />
                    <SPLIT distance="500" swimtime="00:06:03.97" />
                    <SPLIT distance="550" swimtime="00:06:40.63" />
                    <SPLIT distance="600" swimtime="00:07:17.39" />
                    <SPLIT distance="650" swimtime="00:07:55.37" />
                    <SPLIT distance="700" swimtime="00:08:33.30" />
                    <SPLIT distance="750" swimtime="00:09:11.00" />
                    <SPLIT distance="800" swimtime="00:09:48.52" />
                    <SPLIT distance="850" swimtime="00:10:26.44" />
                    <SPLIT distance="900" swimtime="00:11:04.44" />
                    <SPLIT distance="950" swimtime="00:11:42.08" />
                    <SPLIT distance="1000" swimtime="00:12:19.66" />
                    <SPLIT distance="1050" swimtime="00:12:57.85" />
                    <SPLIT distance="1100" swimtime="00:13:35.52" />
                    <SPLIT distance="1150" swimtime="00:14:13.36" />
                    <SPLIT distance="1200" swimtime="00:14:50.61" />
                    <SPLIT distance="1250" swimtime="00:15:28.42" />
                    <SPLIT distance="1300" swimtime="00:16:05.87" />
                    <SPLIT distance="1350" swimtime="00:16:43.62" />
                    <SPLIT distance="1400" swimtime="00:17:21.63" />
                    <SPLIT distance="1450" swimtime="00:17:59.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="545" swimtime="00:02:19.15" resultid="1797" heatid="2171" lane="4" entrytime="00:02:14.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.77" />
                    <SPLIT distance="100" swimtime="00:01:03.80" />
                    <SPLIT distance="150" swimtime="00:01:40.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="584" swimtime="00:02:22.20" resultid="1798" heatid="2155" lane="3" entrytime="00:02:19.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                    <SPLIT distance="100" swimtime="00:01:07.04" />
                    <SPLIT distance="150" swimtime="00:01:48.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" status="WDR" swimtime="00:00:00.00" resultid="1799" entrytime="00:04:30.38" entrycourse="SCM" />
                <RESULT eventid="1364" points="595" swimtime="00:05:02.59" resultid="1800" heatid="2210" lane="3" entrytime="00:04:52.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.98" />
                    <SPLIT distance="100" swimtime="00:01:04.85" />
                    <SPLIT distance="150" swimtime="00:01:45.47" />
                    <SPLIT distance="200" swimtime="00:02:26.36" />
                    <SPLIT distance="250" swimtime="00:03:10.24" />
                    <SPLIT distance="300" swimtime="00:03:53.77" />
                    <SPLIT distance="350" swimtime="00:04:28.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1381" status="RJC" swimtime="00:00:00.00" resultid="1801" entrytime="00:09:16.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ciro" lastname="Adriano Theiss Filho" birthdate="2003-04-01" gender="M" nation="BRA" license="V413283" athleteid="1897" externalid="V413283">
              <RESULTS>
                <RESULT eventid="1178" points="688" swimtime="00:00:30.57" resultid="2148" heatid="2175" lane="1" />
                <RESULT eventid="1485" points="704" swimtime="00:01:05.35" resultid="2149" heatid="2230" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="717" swimtime="00:02:22.48" resultid="2150" heatid="2192" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:07.71" />
                    <SPLIT distance="150" swimtime="00:01:44.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariana" lastname="Matsuda Estevam" birthdate="2004-02-06" gender="F" nation="JPN" license="336748" swrid="5687021" athleteid="1855" externalid="336748">
              <RESULTS>
                <RESULT eventid="1113" points="544" swimtime="00:00:34.15" resultid="1856" heatid="2162" lane="4" entrytime="00:00:33.53" entrycourse="SCM" />
                <RESULT eventid="1273" points="542" swimtime="00:00:30.65" resultid="1857" heatid="2197" lane="2" entrytime="00:00:29.96" entrycourse="SCM" />
                <RESULT eventid="1446" points="538" swimtime="00:00:32.13" resultid="1858" heatid="2224" lane="3" entrytime="00:00:32.01" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirian" lastname="Rose Gouveia" birthdate="1989-10-25" gender="F" nation="BRA" license="V081972" athleteid="1890" externalid="V081972">
              <RESULTS>
                <RESULT eventid="1165" points="308" swimtime="00:03:18.89" resultid="1891" heatid="2172" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                    <SPLIT distance="100" swimtime="00:01:31.86" />
                    <SPLIT distance="150" swimtime="00:02:24.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1325" points="438" swimtime="00:01:20.67" resultid="1892" heatid="2205" lane="3" entrytime="00:01:21.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1247" points="424" swimtime="00:03:20.44" resultid="1893" heatid="2190" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.00" />
                    <SPLIT distance="100" swimtime="00:01:37.90" />
                    <SPLIT distance="150" swimtime="00:02:29.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1351" status="RJC" swimtime="00:00:00.00" resultid="1894" />
                <RESULT eventid="1472" points="415" swimtime="00:01:31.91" resultid="1895" heatid="2229" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="453" swimtime="00:00:35.53" resultid="1896" heatid="2224" lane="2" entrytime="00:00:37.73" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Brotto Lemos" birthdate="2000-05-17" gender="M" nation="BRA" license="121382" swrid="5687004" athleteid="1840" externalid="121382">
              <RESULTS>
                <RESULT eventid="1100" points="616" swimtime="00:00:27.84" resultid="1841" heatid="2157" lane="2" />
                <RESULT eventid="1312" points="565" swimtime="00:02:20.30" resultid="1842" heatid="2204" lane="3" entrytime="00:02:10.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="100" swimtime="00:01:06.61" />
                    <SPLIT distance="150" swimtime="00:01:43.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1364" points="590" swimtime="00:05:03.30" resultid="1843" heatid="2209" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.60" />
                    <SPLIT distance="100" swimtime="00:01:06.00" />
                    <SPLIT distance="150" swimtime="00:01:44.19" />
                    <SPLIT distance="200" swimtime="00:02:23.26" />
                    <SPLIT distance="250" swimtime="00:03:07.29" />
                    <SPLIT distance="300" swimtime="00:03:52.53" />
                    <SPLIT distance="350" swimtime="00:04:28.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="580" swimtime="00:01:02.38" resultid="1844" heatid="2218" lane="3" entrytime="00:00:57.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yoseph" lastname="Rigoni Moraes" birthdate="2006-04-17" gender="M" nation="BRA" license="295182" swrid="5622302" athleteid="1878" externalid="295182">
              <RESULTS>
                <RESULT eventid="1260" points="417" swimtime="00:02:50.68" resultid="1879" heatid="2193" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                    <SPLIT distance="100" swimtime="00:01:18.42" />
                    <SPLIT distance="150" swimtime="00:02:04.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="467" swimtime="00:00:27.41" resultid="1880" heatid="2200" lane="4" entrytime="00:00:26.01" entrycourse="SCM" />
                <RESULT eventid="1485" points="427" swimtime="00:01:17.19" resultid="1881" heatid="2230" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Carolina Lucietto" birthdate="1996-10-21" gender="F" nation="BRA" license="110041" swrid="5687005" athleteid="1826" externalid="110041">
              <RESULTS>
                <RESULT eventid="1061" points="453" swimtime="00:11:31.39" resultid="1827" heatid="2152" lane="4" entrytime="00:11:05.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="600" swimtime="00:08:32.83" />
                    <SPLIT distance="650" swimtime="00:09:17.63" />
                    <SPLIT distance="700" swimtime="00:10:02.65" />
                    <SPLIT distance="750" swimtime="00:10:47.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1299" points="425" swimtime="00:02:53.39" resultid="1828" heatid="2202" lane="4" entrytime="00:02:46.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                    <SPLIT distance="100" swimtime="00:01:24.21" />
                    <SPLIT distance="150" swimtime="00:02:08.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1221" points="476" swimtime="00:05:24.75" resultid="1829" heatid="2186" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:15.36" />
                    <SPLIT distance="150" swimtime="00:01:56.11" />
                    <SPLIT distance="200" swimtime="00:02:37.03" />
                    <SPLIT distance="250" swimtime="00:03:18.66" />
                    <SPLIT distance="300" swimtime="00:04:00.96" />
                    <SPLIT distance="350" swimtime="00:04:44.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" status="WDR" swimtime="00:00:00.00" resultid="1830" heatid="2233" lane="3" entrytime="00:21:22.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Sossai Altoe" birthdate="2006-09-04" gender="M" nation="BRA" license="296488" swrid="5603915" athleteid="1814" externalid="296488">
              <RESULTS>
                <RESULT eventid="1126" points="652" swimtime="00:00:54.68" resultid="1815" heatid="2166" lane="3" entrytime="00:00:52.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="609" swimtime="00:00:25.10" resultid="1816" heatid="2201" lane="2" entrytime="00:00:24.53" entrycourse="SCM" />
                <RESULT eventid="1433" points="611" swimtime="00:02:03.56" resultid="1817" heatid="2223" lane="3" entrytime="00:01:55.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.44" />
                    <SPLIT distance="100" swimtime="00:00:58.07" />
                    <SPLIT distance="150" swimtime="00:01:30.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariana" lastname="Fonseca Faria" birthdate="2003-06-17" gender="F" nation="BRA" license="V250089" swrid="5600162" athleteid="1831" externalid="V250089">
              <RESULTS>
                <RESULT eventid="1087" status="WDR" swimtime="00:00:00.00" resultid="1832" heatid="2156" lane="3" entrytime="00:02:30.16" entrycourse="SCM" />
                <RESULT eventid="1299" status="WDR" swimtime="00:00:00.00" resultid="1833" heatid="2202" lane="3" entrytime="00:02:31.59" entrycourse="SCM" />
                <RESULT eventid="1394" status="WDR" swimtime="00:00:00.00" resultid="1834" heatid="2216" lane="3" entrytime="00:01:08.48" entrycourse="SCM" />
                <RESULT eventid="1420" status="WDR" swimtime="00:00:00.00" resultid="1835" heatid="2219" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isaac" lastname="Guimaraes Saraiva" birthdate="2000-02-02" gender="M" nation="BRA" license="V103705" athleteid="1882" externalid="V103705">
              <RESULTS>
                <RESULT eventid="1100" points="690" swimtime="00:00:26.81" resultid="1883" heatid="2157" lane="3" />
                <RESULT eventid="1312" points="708" swimtime="00:02:10.14" resultid="1884" heatid="2203" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.32" />
                    <SPLIT distance="100" swimtime="00:01:04.04" />
                    <SPLIT distance="150" swimtime="00:01:37.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="698" swimtime="00:00:58.65" resultid="1885" heatid="2217" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diego" lastname="Duarte Rezende" birthdate="2006-01-25" gender="M" nation="BRA" license="313013" swrid="5498173" athleteid="1870" externalid="313013">
              <RESULTS>
                <RESULT eventid="1204" points="484" swimtime="00:19:43.53" resultid="1871" heatid="2181" lane="4" entrytime="00:18:17.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                    <SPLIT distance="100" swimtime="00:01:07.45" />
                    <SPLIT distance="150" swimtime="00:01:44.07" />
                    <SPLIT distance="200" swimtime="00:02:21.02" />
                    <SPLIT distance="250" swimtime="00:02:58.60" />
                    <SPLIT distance="300" swimtime="00:03:37.21" />
                    <SPLIT distance="350" swimtime="00:04:15.69" />
                    <SPLIT distance="400" swimtime="00:04:55.18" />
                    <SPLIT distance="450" swimtime="00:05:34.48" />
                    <SPLIT distance="500" swimtime="00:06:14.74" />
                    <SPLIT distance="550" swimtime="00:06:54.61" />
                    <SPLIT distance="600" swimtime="00:07:34.86" />
                    <SPLIT distance="650" swimtime="00:08:15.46" />
                    <SPLIT distance="700" swimtime="00:08:56.54" />
                    <SPLIT distance="750" swimtime="00:09:36.61" />
                    <SPLIT distance="800" swimtime="00:10:17.03" />
                    <SPLIT distance="850" swimtime="00:10:57.47" />
                    <SPLIT distance="900" swimtime="00:11:38.68" />
                    <SPLIT distance="950" swimtime="00:12:19.85" />
                    <SPLIT distance="1000" swimtime="00:13:00.86" />
                    <SPLIT distance="1050" swimtime="00:13:42.45" />
                    <SPLIT distance="1100" swimtime="00:14:22.56" />
                    <SPLIT distance="1150" swimtime="00:15:03.38" />
                    <SPLIT distance="1200" swimtime="00:15:44.06" />
                    <SPLIT distance="1250" swimtime="00:16:25.27" />
                    <SPLIT distance="1300" swimtime="00:17:04.28" />
                    <SPLIT distance="1350" swimtime="00:17:44.21" />
                    <SPLIT distance="1400" swimtime="00:18:24.90" />
                    <SPLIT distance="1450" swimtime="00:19:05.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="537" swimtime="00:00:29.15" resultid="1872" heatid="2159" lane="3" entrytime="00:00:28.88" entrycourse="SCM" />
                <RESULT eventid="1312" points="436" swimtime="00:02:32.99" resultid="1873" heatid="2204" lane="2" entrytime="00:02:21.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:11.29" />
                    <SPLIT distance="150" swimtime="00:01:51.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="533" swimtime="00:01:04.16" resultid="1874" heatid="2218" lane="4" entrytime="00:01:02.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yohan" lastname="Rigoni Moraes" birthdate="2002-04-03" gender="M" nation="BRA" license="272187" swrid="5600245" athleteid="1851" externalid="272187">
              <RESULTS>
                <RESULT eventid="1178" points="800" swimtime="00:00:29.07" resultid="1852" heatid="2176" lane="2" entrytime="00:00:28.97" entrycourse="SCM" />
                <RESULT eventid="1260" points="601" swimtime="00:02:31.10" resultid="1853" heatid="2194" lane="4" entrytime="00:02:30.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.21" />
                    <SPLIT distance="100" swimtime="00:01:09.16" />
                    <SPLIT distance="150" swimtime="00:01:49.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1485" points="713" swimtime="00:01:05.07" resultid="1854" heatid="2232" lane="4" entrytime="00:01:04.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roberto" lastname="Iuji Nogami" birthdate="1997-09-27" gender="M" nation="BRA" license="V110021" swrid="5687016" athleteid="1848" externalid="V110021">
              <RESULTS>
                <RESULT eventid="1152" status="DNS" swimtime="00:00:00.00" resultid="1849" heatid="2171" lane="3" entrytime="00:02:13.18" entrycourse="SCM" />
                <RESULT eventid="1433" status="DNS" swimtime="00:00:00.00" resultid="1850" heatid="2223" lane="4" entrytime="00:02:01.39" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Felipe Alves" birthdate="2002-05-25" gender="M" nation="BRA" license="347979" athleteid="1886" externalid="347979">
              <RESULTS>
                <RESULT eventid="1126" points="433" swimtime="00:01:02.67" resultid="1887" heatid="2166" lane="1" entrytime="00:01:00.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="380" swimtime="00:05:21.22" resultid="1888" heatid="2188" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                    <SPLIT distance="100" swimtime="00:01:13.12" />
                    <SPLIT distance="150" swimtime="00:01:53.80" />
                    <SPLIT distance="200" swimtime="00:02:35.30" />
                    <SPLIT distance="250" swimtime="00:03:17.44" />
                    <SPLIT distance="300" swimtime="00:04:00.87" />
                    <SPLIT distance="350" swimtime="00:04:44.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="385" swimtime="00:02:24.09" resultid="1889" heatid="2221" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                    <SPLIT distance="100" swimtime="00:01:09.11" />
                    <SPLIT distance="150" swimtime="00:01:47.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Júlio" lastname="Nobuyuki Ito" birthdate="2000-09-14" gender="M" nation="BRA" license="V265311" swrid="5220012" athleteid="1836" externalid="V265311">
              <RESULTS>
                <RESULT eventid="1074" points="637" swimtime="00:02:18.18" resultid="1837" heatid="2153" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                    <SPLIT distance="150" swimtime="00:01:44.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="719" swimtime="00:00:57.35" resultid="1838" heatid="2207" lane="3" entrytime="00:00:56.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1459" points="708" swimtime="00:00:25.97" resultid="1839" heatid="2227" lane="3" entrytime="00:00:25.35" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emily" lastname="Bazan Montanari" birthdate="2003-08-10" gender="F" nation="BRA" license="253944" swrid="5687003" athleteid="1859" externalid="253944">
              <RESULTS>
                <RESULT eventid="1139" points="474" swimtime="00:01:09.80" resultid="1860" heatid="2169" lane="2" entrytime="00:01:10.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="419" swimtime="00:00:40.74" resultid="1861" heatid="2178" lane="2" entrytime="00:00:42.36" entrycourse="SCM" />
                <RESULT eventid="1247" points="406" swimtime="00:03:20.16" resultid="1862" heatid="2190" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.81" />
                    <SPLIT distance="100" swimtime="00:01:32.87" />
                    <SPLIT distance="150" swimtime="00:02:25.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="422" swimtime="00:00:33.32" resultid="1863" heatid="2196" lane="1" />
                <RESULT eventid="1472" points="409" swimtime="00:01:30.03" resultid="1864" heatid="2229" lane="4" entrytime="00:01:29.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Eduardo Rech" birthdate="2010-05-25" gender="M" nation="BRA" license="V413284" athleteid="1903" externalid="V413284">
              <RESULTS>
                <RESULT eventid="1074" status="DSQ" swimtime="00:02:14.11" resultid="1904" heatid="2154" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.32" />
                    <SPLIT distance="100" swimtime="00:01:02.38" />
                    <SPLIT distance="150" swimtime="00:01:43.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="703" swimtime="00:00:57.77" resultid="1905" heatid="2206" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="662" swimtime="00:00:24.41" resultid="1906" heatid="2199" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Pacheco" birthdate="2006-12-20" gender="M" nation="BRA" license="336850" swrid="5603854" athleteid="1875" externalid="336850">
              <RESULTS>
                <RESULT eventid="1152" points="374" swimtime="00:02:37.81" resultid="1876" heatid="2171" lane="2" entrytime="00:02:28.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                    <SPLIT distance="100" swimtime="00:01:08.19" />
                    <SPLIT distance="150" swimtime="00:01:50.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="540" swimtime="00:01:03.07" resultid="1877" heatid="2207" lane="4" entrytime="00:01:02.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Kupicki" birthdate="2004-03-02" gender="F" nation="BRA" license="311897" swrid="5624094" athleteid="1802" externalid="311897">
              <RESULTS>
                <RESULT eventid="1139" points="472" swimtime="00:01:09.88" resultid="1803" heatid="2169" lane="4" entrytime="00:01:06.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="456" swimtime="00:02:58.09" resultid="1804" heatid="2156" lane="4" entrytime="00:02:43.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.09" />
                    <SPLIT distance="150" swimtime="00:02:12.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="428" swimtime="00:00:40.46" resultid="1805" heatid="2177" lane="1" />
                <RESULT eventid="1420" points="443" swimtime="00:02:34.71" resultid="1806" heatid="2220" lane="4" entrytime="00:02:26.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                    <SPLIT distance="100" swimtime="00:01:13.19" />
                    <SPLIT distance="150" swimtime="00:01:52.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Perroni Ribeiro" birthdate="2004-11-06" gender="F" nation="BRA" license="310555" swrid="5727651" athleteid="1818" externalid="310555">
              <RESULTS>
                <RESULT eventid="1061" points="633" swimtime="00:10:18.34" resultid="1819" heatid="2151" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                    <SPLIT distance="100" swimtime="00:01:15.87" />
                    <SPLIT distance="150" swimtime="00:01:54.88" />
                    <SPLIT distance="200" swimtime="00:02:33.95" />
                    <SPLIT distance="250" swimtime="00:03:12.63" />
                    <SPLIT distance="300" swimtime="00:03:51.36" />
                    <SPLIT distance="350" swimtime="00:04:30.57" />
                    <SPLIT distance="400" swimtime="00:05:09.81" />
                    <SPLIT distance="450" swimtime="00:05:48.52" />
                    <SPLIT distance="500" swimtime="00:06:27.38" />
                    <SPLIT distance="550" swimtime="00:07:05.85" />
                    <SPLIT distance="600" swimtime="00:07:44.48" />
                    <SPLIT distance="650" swimtime="00:08:22.98" />
                    <SPLIT distance="700" swimtime="00:09:01.70" />
                    <SPLIT distance="750" swimtime="00:09:39.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1221" points="600" swimtime="00:05:00.79" resultid="1820" heatid="2186" lane="3" entrytime="00:04:47.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                    <SPLIT distance="100" swimtime="00:01:13.19" />
                    <SPLIT distance="150" swimtime="00:01:51.42" />
                    <SPLIT distance="200" swimtime="00:02:29.74" />
                    <SPLIT distance="250" swimtime="00:03:07.70" />
                    <SPLIT distance="300" swimtime="00:03:45.80" />
                    <SPLIT distance="350" swimtime="00:04:23.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="670" swimtime="00:18:58.23" resultid="1821" heatid="2234" lane="3" entrytime="00:18:09.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:14.54" />
                    <SPLIT distance="150" swimtime="00:01:53.65" />
                    <SPLIT distance="200" swimtime="00:02:32.13" />
                    <SPLIT distance="250" swimtime="00:03:11.20" />
                    <SPLIT distance="300" swimtime="00:03:49.67" />
                    <SPLIT distance="350" swimtime="00:04:27.76" />
                    <SPLIT distance="400" swimtime="00:05:05.91" />
                    <SPLIT distance="450" swimtime="00:05:43.76" />
                    <SPLIT distance="500" swimtime="00:06:21.78" />
                    <SPLIT distance="550" swimtime="00:06:59.50" />
                    <SPLIT distance="600" swimtime="00:07:37.33" />
                    <SPLIT distance="650" swimtime="00:08:15.09" />
                    <SPLIT distance="700" swimtime="00:08:53.21" />
                    <SPLIT distance="750" swimtime="00:09:31.05" />
                    <SPLIT distance="800" swimtime="00:10:08.88" />
                    <SPLIT distance="850" swimtime="00:10:46.98" />
                    <SPLIT distance="900" swimtime="00:11:24.95" />
                    <SPLIT distance="950" swimtime="00:12:02.59" />
                    <SPLIT distance="1000" swimtime="00:12:40.55" />
                    <SPLIT distance="1050" swimtime="00:13:18.73" />
                    <SPLIT distance="1100" swimtime="00:13:56.71" />
                    <SPLIT distance="1150" swimtime="00:14:34.93" />
                    <SPLIT distance="1200" swimtime="00:15:12.52" />
                    <SPLIT distance="1250" swimtime="00:15:49.87" />
                    <SPLIT distance="1300" swimtime="00:16:27.82" />
                    <SPLIT distance="1350" swimtime="00:17:05.48" />
                    <SPLIT distance="1400" swimtime="00:17:43.70" />
                    <SPLIT distance="1450" swimtime="00:18:21.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jordana" lastname="Rinaldini" birthdate="2004-09-13" gender="F" nation="BRA" license="342426" swrid="5596933" athleteid="1807" externalid="342426">
              <RESULTS>
                <RESULT eventid="1113" points="495" swimtime="00:00:35.24" resultid="1808" heatid="2160" lane="3" />
                <RESULT eventid="1191" points="469" swimtime="00:00:39.25" resultid="1809" heatid="2178" lane="3" entrytime="00:00:39.14" entrycourse="SCM" />
                <RESULT eventid="1247" points="503" swimtime="00:03:06.45" resultid="1810" heatid="2191" lane="3" entrytime="00:03:01.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.05" />
                    <SPLIT distance="100" swimtime="00:01:27.63" />
                    <SPLIT distance="150" swimtime="00:02:16.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1351" points="403" swimtime="00:06:25.63" resultid="1811" heatid="2208" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                    <SPLIT distance="150" swimtime="00:02:18.30" />
                    <SPLIT distance="200" swimtime="00:03:08.42" />
                    <SPLIT distance="250" swimtime="00:03:59.92" />
                    <SPLIT distance="300" swimtime="00:04:52.46" />
                    <SPLIT distance="350" swimtime="00:05:39.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1394" points="468" swimtime="00:01:18.04" resultid="1812" heatid="2216" lane="5" entrytime="00:01:18.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1472" status="RJC" swimtime="00:00:00.00" resultid="1813" entrytime="00:01:24.46" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nayara" lastname="Moreira Baron" birthdate="2001-05-15" gender="F" nation="BRA" license="V413285" athleteid="1907" externalid="V413285">
              <RESULTS>
                <RESULT eventid="1139" points="618" swimtime="00:01:03.89" resultid="1908" heatid="2168" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="549" swimtime="00:02:47.44" resultid="1909" heatid="2156" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.95" />
                    <SPLIT distance="100" swimtime="00:01:19.21" />
                    <SPLIT distance="150" swimtime="00:02:07.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1221" points="575" swimtime="00:05:05.05" resultid="1910" heatid="2186" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                    <SPLIT distance="150" swimtime="00:01:52.00" />
                    <SPLIT distance="200" swimtime="00:02:30.83" />
                    <SPLIT distance="250" swimtime="00:03:09.44" />
                    <SPLIT distance="300" swimtime="00:03:47.76" />
                    <SPLIT distance="350" swimtime="00:04:26.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="630" swimtime="00:00:29.15" resultid="1911" heatid="2196" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernando" lastname="Fumagalli" birthdate="1998-08-16" gender="M" nation="BRA" license="V117756" swrid="5687007" athleteid="1845" externalid="V117756">
              <RESULTS>
                <RESULT eventid="1178" points="595" swimtime="00:00:32.08" resultid="1846" heatid="2174" lane="2" />
                <RESULT eventid="1459" points="702" swimtime="00:00:26.04" resultid="1847" heatid="2227" lane="2" entrytime="00:00:25.83" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="UNICESUMAR (MARINGÃ) &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1219" swimtime="00:03:34.94" resultid="1915" heatid="2184" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.75" />
                    <SPLIT distance="100" swimtime="00:00:55.05" />
                    <SPLIT distance="150" swimtime="00:01:20.00" />
                    <SPLIT distance="200" swimtime="00:01:47.90" />
                    <SPLIT distance="250" swimtime="00:02:12.17" />
                    <SPLIT distance="300" swimtime="00:02:39.79" />
                    <SPLIT distance="350" swimtime="00:03:05.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1814" number="1" />
                    <RELAYPOSITION athleteid="1836" number="2" />
                    <RELAYPOSITION athleteid="1903" number="3" />
                    <RELAYPOSITION athleteid="1882" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1379" swimtime="00:08:27.28" resultid="1916" heatid="2212" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.37" />
                    <SPLIT distance="100" swimtime="00:00:57.66" />
                    <SPLIT distance="150" swimtime="00:01:30.25" />
                    <SPLIT distance="200" swimtime="00:02:04.15" />
                    <SPLIT distance="250" swimtime="00:02:31.42" />
                    <SPLIT distance="300" swimtime="00:03:02.52" />
                    <SPLIT distance="350" swimtime="00:03:34.66" />
                    <SPLIT distance="400" swimtime="00:04:02.56" />
                    <SPLIT distance="450" swimtime="00:04:29.35" />
                    <SPLIT distance="500" swimtime="00:05:01.18" />
                    <SPLIT distance="550" swimtime="00:05:35.28" />
                    <SPLIT distance="600" swimtime="00:06:07.32" />
                    <SPLIT distance="650" swimtime="00:06:39.54" />
                    <SPLIT distance="700" swimtime="00:07:14.69" />
                    <SPLIT distance="750" swimtime="00:07:52.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1814" number="1" />
                    <RELAYPOSITION athleteid="1903" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1897" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1840" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" swimtime="00:04:00.14" resultid="1917" heatid="2236" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.79" />
                    <SPLIT distance="100" swimtime="00:01:00.78" />
                    <SPLIT distance="150" swimtime="00:01:31.01" />
                    <SPLIT distance="200" swimtime="00:02:06.12" />
                    <SPLIT distance="250" swimtime="00:02:33.71" />
                    <SPLIT distance="300" swimtime="00:03:05.90" />
                    <SPLIT distance="350" swimtime="00:03:31.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1882" number="1" />
                    <RELAYPOSITION athleteid="1851" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1836" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1845" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="UNICESUMAR (MARINGÁ) &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1217" swimtime="00:04:30.75" resultid="1912" heatid="2182" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                    <SPLIT distance="100" swimtime="00:01:04.79" />
                    <SPLIT distance="150" swimtime="00:01:37.33" />
                    <SPLIT distance="200" swimtime="00:02:15.37" />
                    <SPLIT distance="250" swimtime="00:02:47.73" />
                    <SPLIT distance="300" swimtime="00:03:21.76" />
                    <SPLIT distance="350" swimtime="00:03:54.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1907" number="1" />
                    <RELAYPOSITION athleteid="1807" number="2" />
                    <RELAYPOSITION athleteid="1818" number="3" />
                    <RELAYPOSITION athleteid="1802" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1377" swimtime="00:10:09.48" resultid="1913" heatid="2211" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                    <SPLIT distance="100" swimtime="00:01:08.11" />
                    <SPLIT distance="150" swimtime="00:01:45.39" />
                    <SPLIT distance="200" swimtime="00:02:22.55" />
                    <SPLIT distance="250" swimtime="00:02:56.22" />
                    <SPLIT distance="300" swimtime="00:03:35.99" />
                    <SPLIT distance="350" swimtime="00:04:21.23" />
                    <SPLIT distance="400" swimtime="00:05:07.12" />
                    <SPLIT distance="450" swimtime="00:05:41.79" />
                    <SPLIT distance="500" swimtime="00:06:19.20" />
                    <SPLIT distance="550" swimtime="00:06:56.97" />
                    <SPLIT distance="600" swimtime="00:07:34.04" />
                    <SPLIT distance="650" swimtime="00:08:09.42" />
                    <SPLIT distance="700" swimtime="00:08:48.35" />
                    <SPLIT distance="750" swimtime="00:09:28.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1907" number="1" />
                    <RELAYPOSITION athleteid="1855" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1818" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1826" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1513" swimtime="00:05:06.39" resultid="1914" heatid="2237" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                    <SPLIT distance="100" swimtime="00:01:16.11" />
                    <SPLIT distance="150" swimtime="00:01:55.50" />
                    <SPLIT distance="200" swimtime="00:02:40.43" />
                    <SPLIT distance="250" swimtime="00:03:15.83" />
                    <SPLIT distance="300" swimtime="00:03:58.08" />
                    <SPLIT distance="350" swimtime="00:04:30.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1826" number="1" />
                    <RELAYPOSITION athleteid="1807" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1907" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1802" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4008" nation="BRA" region="PR" clubid="1610" name="Uem (Maringá)">
          <ATHLETES>
            <ATHLETE firstname="Juliano" lastname="Ito" birthdate="2002-11-21" gender="M" nation="BRA" license="V281999" swrid="5687015" athleteid="1611" externalid="V281999">
              <RESULTS>
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="1612" heatid="2155" lane="1" entrytime="00:02:22.70" entrycourse="SCM" />
                <RESULT eventid="1100" status="DNS" swimtime="00:00:00.00" resultid="1613" heatid="2159" lane="1" entrytime="00:00:30.02" entrycourse="SCM" />
                <RESULT eventid="1312" status="DNS" swimtime="00:00:00.00" resultid="1614" heatid="2204" lane="5" entrytime="00:02:29.58" entrycourse="SCM" />
                <RESULT eventid="1364" status="DNS" swimtime="00:00:00.00" resultid="1615" heatid="2210" lane="4" entrytime="00:05:25.12" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose" lastname="Vinicius Poletto" birthdate="2000-03-29" gender="M" nation="BRA" license="V294183" athleteid="1655" externalid="V294183">
              <RESULTS>
                <RESULT eventid="1152" points="227" swimtime="00:03:06.40" resultid="1656" heatid="2170" lane="4" entrytime="00:02:58.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:20.39" />
                    <SPLIT distance="150" swimtime="00:02:10.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="350" swimtime="00:01:12.89" resultid="1657" heatid="2207" lane="5" entrytime="00:01:10.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="338" swimtime="00:05:34.15" resultid="1658" heatid="2189" lane="3" entrytime="00:05:21.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:15.87" />
                    <SPLIT distance="150" swimtime="00:01:57.10" />
                    <SPLIT distance="200" swimtime="00:02:39.50" />
                    <SPLIT distance="250" swimtime="00:03:21.84" />
                    <SPLIT distance="300" swimtime="00:04:03.61" />
                    <SPLIT distance="350" swimtime="00:04:44.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1459" points="428" swimtime="00:00:30.71" resultid="1659" heatid="2226" lane="4" entrytime="00:00:29.88" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Gabriel Dumont Negrelli" birthdate="1999-12-29" gender="M" nation="BRA" license="V413201" athleteid="1627" externalid="V413201">
              <RESULTS>
                <RESULT eventid="1260" points="179" swimtime="00:03:45.91" resultid="1628" heatid="2192" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.64" />
                    <SPLIT distance="100" swimtime="00:01:42.80" />
                    <SPLIT distance="150" swimtime="00:02:43.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="275" swimtime="00:00:32.69" resultid="1629" heatid="2198" lane="5" />
                <RESULT eventid="1433" points="164" swimtime="00:03:11.39" resultid="1630" heatid="2222" lane="5" entrytime="00:03:06.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.05" />
                    <SPLIT distance="100" swimtime="00:01:27.75" />
                    <SPLIT distance="150" swimtime="00:02:19.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Henrique Antunes" birthdate="2003-11-23" gender="M" nation="BRA" license="V318505" athleteid="1666" externalid="V318505">
              <RESULTS>
                <RESULT eventid="1126" points="388" swimtime="00:01:05.00" resultid="1667" heatid="2165" lane="4" entrytime="00:01:03.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="445" swimtime="00:00:27.87" resultid="1668" heatid="2200" lane="5" entrytime="00:00:27.88" entrycourse="SCM" />
                <RESULT eventid="1433" points="205" swimtime="00:02:57.70" resultid="1669" heatid="2222" lane="4" entrytime="00:02:30.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                    <SPLIT distance="100" swimtime="00:01:28.69" />
                    <SPLIT distance="150" swimtime="00:02:18.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Johnny" lastname="Paulo Ito" birthdate="2005-03-31" gender="M" nation="BRA" license="282600" swrid="5687025" athleteid="1616" externalid="282600">
              <RESULTS>
                <RESULT eventid="1074" points="445" swimtime="00:02:35.65" resultid="1617" heatid="2155" lane="2" entrytime="00:02:30.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="100" swimtime="00:01:10.30" />
                    <SPLIT distance="150" swimtime="00:01:54.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="545" swimtime="00:00:33.03" resultid="1618" heatid="2175" lane="3" entrytime="00:00:35.84" entrycourse="SCM" />
                <RESULT eventid="1260" points="422" swimtime="00:02:49.95" resultid="1619" heatid="2194" lane="1" entrytime="00:02:50.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                    <SPLIT distance="100" swimtime="00:01:20.71" />
                    <SPLIT distance="150" swimtime="00:02:05.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1364" points="376" swimtime="00:05:52.41" resultid="1620" heatid="2210" lane="2" entrytime="00:05:41.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                    <SPLIT distance="100" swimtime="00:01:12.78" />
                    <SPLIT distance="150" swimtime="00:01:58.51" />
                    <SPLIT distance="200" swimtime="00:02:45.17" />
                    <SPLIT distance="250" swimtime="00:03:31.14" />
                    <SPLIT distance="300" swimtime="00:04:20.12" />
                    <SPLIT distance="350" swimtime="00:05:08.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1485" points="494" swimtime="00:01:13.54" resultid="1621" heatid="2231" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Zanetti Finotti" birthdate="1999-06-11" gender="M" nation="BRA" license="V413217" athleteid="1643" externalid="V413217">
              <RESULTS>
                <RESULT eventid="1178" points="138" swimtime="00:00:52.22" resultid="1644" heatid="2175" lane="2" entrytime="00:00:54.57" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinícius" lastname="Schuch Pimpão" birthdate="2006-12-16" gender="M" nation="BRA" license="V327807" athleteid="1670" externalid="V327807">
              <RESULTS>
                <RESULT eventid="1100" points="398" swimtime="00:00:32.21" resultid="1671" heatid="2159" lane="4" entrytime="00:00:32.84" entrycourse="SCM" />
                <RESULT eventid="1312" points="352" swimtime="00:02:44.20" resultid="1672" heatid="2203" lane="4" entrytime="00:02:44.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                    <SPLIT distance="100" swimtime="00:01:17.37" />
                    <SPLIT distance="150" swimtime="00:01:59.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="388" swimtime="00:01:11.35" resultid="1673" heatid="2217" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Marcelo Baessa Da Silva" birthdate="2005-12-03" gender="M" nation="BRA" license="V413289" athleteid="1688" externalid="V413289">
              <RESULTS>
                <RESULT eventid="1074" status="DSQ" swimtime="00:03:30.57" resultid="1689" heatid="2154" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="100" swimtime="00:01:23.70" />
                    <SPLIT distance="150" swimtime="00:02:34.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="260" swimtime="00:01:20.44" resultid="1690" heatid="2206" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1459" points="354" swimtime="00:00:32.71" resultid="1691" heatid="2225" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Padovan Otani" birthdate="2000-01-28" gender="F" nation="BRA" license="V413207" athleteid="1631" externalid="V413207">
              <RESULTS>
                <RESULT eventid="1113" points="190" swimtime="00:00:48.49" resultid="1632" heatid="2160" lane="4" />
                <RESULT eventid="1191" points="120" swimtime="00:01:01.77" resultid="1633" heatid="2177" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Lima Barbosa" birthdate="2002-07-01" gender="F" nation="BRA" license="V413208" athleteid="1634" externalid="V413208">
              <RESULTS>
                <RESULT eventid="1113" points="239" swimtime="00:00:44.88" resultid="1635" heatid="2162" lane="1" entrytime="00:00:44.18" entrycourse="SCM" />
                <RESULT eventid="1273" points="293" swimtime="00:00:37.60" resultid="1636" heatid="2195" lane="3" />
                <RESULT eventid="1394" points="215" swimtime="00:01:41.16" resultid="1637" heatid="2215" lane="3" entrytime="00:01:39.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitoria" lastname="Alice Martins" birthdate="1999-01-19" gender="F" nation="BRA" license="V383078" swrid="5687002" athleteid="1622" externalid="V383078">
              <RESULTS>
                <RESULT eventid="1113" points="307" swimtime="00:00:41.29" resultid="1623" heatid="2162" lane="2" entrytime="00:00:38.99" entrycourse="SCM" />
                <RESULT eventid="1221" points="232" swimtime="00:06:52.83" resultid="1624" heatid="2186" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.20" />
                    <SPLIT distance="100" swimtime="00:01:33.88" />
                    <SPLIT distance="150" swimtime="00:02:24.68" />
                    <SPLIT distance="200" swimtime="00:03:17.54" />
                    <SPLIT distance="250" swimtime="00:04:11.07" />
                    <SPLIT distance="300" swimtime="00:05:06.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1394" points="282" swimtime="00:01:32.44" resultid="1625" heatid="2216" lane="1" entrytime="00:01:30.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="179" swimtime="00:00:46.35" resultid="1626" heatid="2224" lane="5" entrytime="00:00:48.26" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Luisa Batista" birthdate="2001-05-30" gender="F" nation="BRA" license="V413214" athleteid="1638" externalid="V413214">
              <RESULTS>
                <RESULT eventid="1139" status="WDR" swimtime="00:00:00.00" resultid="1639" />
                <RESULT eventid="1191" status="WDR" swimtime="00:00:00.00" resultid="1640" entrytime="00:00:50.32" entrycourse="SCM" />
                <RESULT eventid="1273" status="WDR" swimtime="00:00:00.00" resultid="1641" entrytime="00:00:37.93" entrycourse="SCM" />
                <RESULT eventid="1472" status="WDR" swimtime="00:00:00.00" resultid="1642" entrytime="00:01:53.21" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Ortega" birthdate="1999-08-05" gender="M" nation="BRA" license="383118" swrid="5603852" athleteid="1674" externalid="383118">
              <RESULTS>
                <RESULT eventid="1100" points="400" swimtime="00:00:32.15" resultid="1675" heatid="2159" lane="2" entrytime="00:00:30.98" entrycourse="SCM" />
                <RESULT eventid="1312" points="396" swimtime="00:02:37.94" resultid="1676" heatid="2204" lane="1" entrytime="00:02:29.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                    <SPLIT distance="100" swimtime="00:01:16.03" />
                    <SPLIT distance="150" swimtime="00:01:58.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="345" swimtime="00:05:31.91" resultid="1677" heatid="2189" lane="1" entrytime="00:05:16.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                    <SPLIT distance="100" swimtime="00:01:15.16" />
                    <SPLIT distance="150" swimtime="00:01:56.66" />
                    <SPLIT distance="200" swimtime="00:02:38.43" />
                    <SPLIT distance="250" swimtime="00:03:21.54" />
                    <SPLIT distance="300" swimtime="00:04:04.65" />
                    <SPLIT distance="350" swimtime="00:04:47.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1407" points="388" swimtime="00:01:11.32" resultid="1678" heatid="2218" lane="2" entrytime="00:01:06.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1381" points="343" swimtime="00:11:36.57" resultid="1679" heatid="2214" lane="1" entrytime="00:11:01.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="100" swimtime="00:01:16.16" />
                    <SPLIT distance="150" swimtime="00:01:57.99" />
                    <SPLIT distance="200" swimtime="00:02:42.26" />
                    <SPLIT distance="250" swimtime="00:03:26.42" />
                    <SPLIT distance="300" swimtime="00:04:10.98" />
                    <SPLIT distance="350" swimtime="00:04:56.17" />
                    <SPLIT distance="400" swimtime="00:05:41.94" />
                    <SPLIT distance="450" swimtime="00:06:26.58" />
                    <SPLIT distance="500" swimtime="00:07:12.31" />
                    <SPLIT distance="550" swimtime="00:07:57.73" />
                    <SPLIT distance="600" swimtime="00:08:43.21" />
                    <SPLIT distance="650" swimtime="00:09:27.92" />
                    <SPLIT distance="700" swimtime="00:10:12.83" />
                    <SPLIT distance="750" swimtime="00:10:57.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Ruivo Costa" birthdate="1995-08-19" gender="M" nation="BRA" license="V110158" athleteid="1651" externalid="V110158">
              <RESULTS>
                <RESULT eventid="1126" points="461" swimtime="00:01:01.37" resultid="1652" heatid="2164" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="338" swimtime="00:01:13.69" resultid="1653" heatid="2207" lane="2" entrytime="00:01:10.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1459" points="455" swimtime="00:00:30.09" resultid="1654" heatid="2227" lane="1" entrytime="00:00:29.63" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Camila Cuenca" birthdate="2005-10-06" gender="F" nation="BRA" license="308081" swrid="5357445" athleteid="1660" externalid="308081">
              <RESULTS>
                <RESULT eventid="1139" points="578" swimtime="00:01:05.35" resultid="1661" heatid="2169" lane="3" entrytime="00:01:05.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1061" points="524" swimtime="00:10:58.85" resultid="1662" heatid="2152" lane="3" entrytime="00:10:35.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.94" />
                    <SPLIT distance="100" swimtime="00:01:15.21" />
                    <SPLIT distance="150" swimtime="00:01:55.59" />
                    <SPLIT distance="200" swimtime="00:02:36.60" />
                    <SPLIT distance="250" swimtime="00:03:17.86" />
                    <SPLIT distance="300" swimtime="00:03:59.74" />
                    <SPLIT distance="350" swimtime="00:04:41.73" />
                    <SPLIT distance="400" swimtime="00:05:24.06" />
                    <SPLIT distance="450" swimtime="00:06:06.26" />
                    <SPLIT distance="500" swimtime="00:06:48.24" />
                    <SPLIT distance="550" swimtime="00:07:30.59" />
                    <SPLIT distance="600" swimtime="00:08:12.99" />
                    <SPLIT distance="650" swimtime="00:08:54.75" />
                    <SPLIT distance="700" swimtime="00:09:36.01" />
                    <SPLIT distance="750" swimtime="00:10:18.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="625" swimtime="00:00:29.24" resultid="1663" heatid="2197" lane="3" entrytime="00:00:29.56" entrycourse="SCM" />
                <RESULT eventid="1394" points="526" swimtime="00:01:15.07" resultid="1664" heatid="2216" lane="2" entrytime="00:01:16.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1420" points="496" swimtime="00:02:29.03" resultid="1665" heatid="2220" lane="3" entrytime="00:02:22.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                    <SPLIT distance="150" swimtime="00:01:50.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Miguel Cardoso" birthdate="2004-09-23" gender="M" nation="BRA" license="V352541" athleteid="1680" externalid="V352541">
              <RESULTS>
                <RESULT eventid="1286" points="325" swimtime="00:00:30.93" resultid="1681" heatid="2198" lane="2" />
                <RESULT eventid="1407" points="159" swimtime="00:01:35.93" resultid="1682" heatid="2218" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1485" points="235" swimtime="00:01:34.18" resultid="1683" heatid="2231" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="De Lacerda Silverio" birthdate="2004-12-29" gender="M" nation="BRA" license="V413223" athleteid="1645" externalid="V413223">
              <RESULTS>
                <RESULT eventid="1126" points="440" swimtime="00:01:02.35" resultid="1646" heatid="2163" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="349" swimtime="00:00:38.31" resultid="1647" heatid="2173" lane="4" />
                <RESULT eventid="1260" points="243" swimtime="00:03:24.34" resultid="1648" heatid="2193" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.08" />
                    <SPLIT distance="100" swimtime="00:01:37.15" />
                    <SPLIT distance="150" swimtime="00:02:30.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1485" points="305" swimtime="00:01:26.33" resultid="1649" heatid="2231" lane="3" entrytime="00:01:23.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="358" swimtime="00:02:27.66" resultid="1650" heatid="2221" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                    <SPLIT distance="100" swimtime="00:01:10.50" />
                    <SPLIT distance="150" swimtime="00:01:50.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diego" lastname="Garcia Costa" birthdate="2003-05-26" gender="M" nation="BRA" license="V413288" athleteid="1684" externalid="V413288">
              <RESULTS>
                <RESULT eventid="1204" points="128" swimtime="00:30:42.71" resultid="1685" heatid="2180" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:01:28.89" />
                    <SPLIT distance="150" swimtime="00:02:20.85" />
                    <SPLIT distance="200" swimtime="00:03:17.74" />
                    <SPLIT distance="250" swimtime="00:04:16.40" />
                    <SPLIT distance="300" swimtime="00:05:14.93" />
                    <SPLIT distance="350" swimtime="00:06:17.55" />
                    <SPLIT distance="400" swimtime="00:07:20.61" />
                    <SPLIT distance="450" swimtime="00:08:21.74" />
                    <SPLIT distance="500" swimtime="00:09:24.06" />
                    <SPLIT distance="550" swimtime="00:10:27.27" />
                    <SPLIT distance="600" swimtime="00:11:31.24" />
                    <SPLIT distance="650" swimtime="00:12:34.99" />
                    <SPLIT distance="700" swimtime="00:13:39.55" />
                    <SPLIT distance="750" swimtime="00:14:43.66" />
                    <SPLIT distance="800" swimtime="00:15:47.93" />
                    <SPLIT distance="850" swimtime="00:16:52.96" />
                    <SPLIT distance="900" swimtime="00:17:58.85" />
                    <SPLIT distance="950" swimtime="00:19:05.30" />
                    <SPLIT distance="1000" swimtime="00:20:11.26" />
                    <SPLIT distance="1050" swimtime="00:21:17.97" />
                    <SPLIT distance="1100" swimtime="00:22:23.62" />
                    <SPLIT distance="1150" swimtime="00:23:29.35" />
                    <SPLIT distance="1200" swimtime="00:24:33.23" />
                    <SPLIT distance="1250" swimtime="00:25:36.43" />
                    <SPLIT distance="1300" swimtime="00:26:38.89" />
                    <SPLIT distance="1350" swimtime="00:27:39.03" />
                    <SPLIT distance="1400" swimtime="00:28:41.75" />
                    <SPLIT distance="1450" swimtime="00:29:44.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="147" swimtime="00:07:20.29" resultid="1686" heatid="2188" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:01:26.72" />
                    <SPLIT distance="150" swimtime="00:02:23.04" />
                    <SPLIT distance="200" swimtime="00:03:21.91" />
                    <SPLIT distance="250" swimtime="00:04:22.26" />
                    <SPLIT distance="300" swimtime="00:05:21.51" />
                    <SPLIT distance="350" swimtime="00:06:22.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1381" points="151" swimtime="00:15:15.15" resultid="1687" heatid="2213" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.58" />
                    <SPLIT distance="100" swimtime="00:01:33.96" />
                    <SPLIT distance="150" swimtime="00:02:27.58" />
                    <SPLIT distance="200" swimtime="00:03:23.54" />
                    <SPLIT distance="250" swimtime="00:04:20.96" />
                    <SPLIT distance="300" swimtime="00:05:19.88" />
                    <SPLIT distance="350" swimtime="00:06:18.89" />
                    <SPLIT distance="400" swimtime="00:07:18.40" />
                    <SPLIT distance="450" swimtime="00:08:18.90" />
                    <SPLIT distance="500" swimtime="00:09:18.30" />
                    <SPLIT distance="550" swimtime="00:10:18.93" />
                    <SPLIT distance="600" swimtime="00:11:19.25" />
                    <SPLIT distance="650" swimtime="00:12:19.65" />
                    <SPLIT distance="700" swimtime="00:13:19.77" />
                    <SPLIT distance="750" swimtime="00:14:19.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="UEM (MARINGÃ) &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1219" swimtime="00:04:08.05" resultid="1695" heatid="2184" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.31" />
                    <SPLIT distance="100" swimtime="00:00:59.27" />
                    <SPLIT distance="150" swimtime="00:01:28.14" />
                    <SPLIT distance="200" swimtime="00:02:01.32" />
                    <SPLIT distance="250" swimtime="00:02:30.49" />
                    <SPLIT distance="300" swimtime="00:03:05.78" />
                    <SPLIT distance="350" swimtime="00:03:34.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1616" number="1" />
                    <RELAYPOSITION athleteid="1651" number="2" />
                    <RELAYPOSITION athleteid="1674" number="3" />
                    <RELAYPOSITION athleteid="1645" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1379" swimtime="00:09:44.72" resultid="1696" heatid="2212" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:07.19" />
                    <SPLIT distance="150" swimtime="00:01:44.45" />
                    <SPLIT distance="200" swimtime="00:02:23.17" />
                    <SPLIT distance="250" swimtime="00:02:55.52" />
                    <SPLIT distance="300" swimtime="00:03:32.11" />
                    <SPLIT distance="350" swimtime="00:04:10.74" />
                    <SPLIT distance="400" swimtime="00:04:47.55" />
                    <SPLIT distance="450" swimtime="00:05:20.82" />
                    <SPLIT distance="500" swimtime="00:06:00.02" />
                    <SPLIT distance="550" swimtime="00:06:41.43" />
                    <SPLIT distance="600" swimtime="00:07:25.58" />
                    <SPLIT distance="650" swimtime="00:07:54.37" />
                    <SPLIT distance="700" swimtime="00:08:28.44" />
                    <SPLIT distance="750" swimtime="00:09:05.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1645" number="1" />
                    <RELAYPOSITION athleteid="1655" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1666" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1616" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" swimtime="00:04:42.09" resultid="1697" heatid="2236" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                    <SPLIT distance="150" swimtime="00:01:44.58" />
                    <SPLIT distance="200" swimtime="00:02:28.79" />
                    <SPLIT distance="250" swimtime="00:03:01.28" />
                    <SPLIT distance="300" swimtime="00:03:39.79" />
                    <SPLIT distance="350" swimtime="00:04:08.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1670" number="1" />
                    <RELAYPOSITION athleteid="1666" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1655" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1674" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="UEM (MARINGÁ) &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1217" swimtime="00:05:30.85" resultid="1692" heatid="2182" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                    <SPLIT distance="100" swimtime="00:01:05.67" />
                    <SPLIT distance="150" swimtime="00:01:45.08" />
                    <SPLIT distance="200" swimtime="00:02:28.37" />
                    <SPLIT distance="250" swimtime="00:03:09.89" />
                    <SPLIT distance="300" swimtime="00:04:03.09" />
                    <SPLIT distance="350" swimtime="00:04:43.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1660" number="1" />
                    <RELAYPOSITION athleteid="1622" number="2" />
                    <RELAYPOSITION athleteid="1631" number="3" />
                    <RELAYPOSITION athleteid="1634" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1377" status="WDR" swimtime="00:00:00.00" resultid="1693" heatid="2211" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="2" reactiontime="0" />
                    <RELAYPOSITION number="3" reactiontime="0" />
                    <RELAYPOSITION number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1513" swimtime="00:06:35.45" resultid="1694" heatid="2237" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.54" />
                    <SPLIT distance="100" swimtime="00:01:40.44" />
                    <SPLIT distance="150" swimtime="00:02:34.21" />
                    <SPLIT distance="200" swimtime="00:03:36.67" />
                    <SPLIT distance="250" swimtime="00:04:17.89" />
                    <SPLIT distance="300" swimtime="00:05:05.12" />
                    <SPLIT distance="350" swimtime="00:05:46.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1634" number="1" />
                    <RELAYPOSITION athleteid="1622" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1660" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1631" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6608" nation="BRA" region="PR" clubid="1532" name="Pucpr (Curitiba)">
          <ATHLETES>
            <ATHLETE firstname="Pedro" lastname="Henrique Araujo" birthdate="2003-11-09" gender="M" nation="BRA" license="307551" athleteid="1561" externalid="307551">
              <RESULTS>
                <RESULT eventid="1126" points="661" swimtime="00:00:54.44" resultid="1562" heatid="2165" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="508" swimtime="00:01:04.37" resultid="1563" heatid="2207" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="567" swimtime="00:02:06.67" resultid="1564" heatid="2222" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="100" swimtime="00:01:01.42" />
                    <SPLIT distance="150" swimtime="00:01:33.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Victor Araujo" birthdate="2001-12-29" gender="M" nation="BRA" license="281163" athleteid="1549" externalid="281163">
              <RESULTS>
                <RESULT eventid="1178" points="823" swimtime="00:00:28.79" resultid="1550" heatid="2176" lane="4" entrytime="00:00:28.92" entrycourse="SCM" />
                <RESULT eventid="1260" points="680" swimtime="00:02:25.02" resultid="1551" heatid="2194" lane="3" entrytime="00:02:26.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="100" swimtime="00:01:09.03" />
                    <SPLIT distance="150" swimtime="00:01:45.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1485" points="756" swimtime="00:01:03.80" resultid="1552" heatid="2232" lane="3" entrytime="00:01:02.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Campesi" birthdate="2004-10-30" gender="M" nation="BRA" license="V383112" athleteid="1577" externalid="V383112">
              <RESULTS>
                <RESULT eventid="1126" points="527" swimtime="00:00:58.71" resultid="1578" heatid="2166" lane="5" entrytime="00:00:58.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="550" swimtime="00:00:25.96" resultid="1579" heatid="2200" lane="3" entrytime="00:00:25.90" entrycourse="SCM" />
                <RESULT eventid="1459" points="433" swimtime="00:00:30.60" resultid="1580" heatid="2226" lane="2" entrytime="00:00:30.92" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="David" lastname="Nycholas Fernandes" birthdate="2000-07-02" gender="M" nation="BRA" license="V312500" athleteid="1565" externalid="V312500">
              <RESULTS>
                <RESULT eventid="1204" points="254" swimtime="00:24:26.11" resultid="1566" heatid="2180" lane="3" entrytime="00:22:27.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                    <SPLIT distance="100" swimtime="00:01:11.66" />
                    <SPLIT distance="150" swimtime="00:01:51.22" />
                    <SPLIT distance="200" swimtime="00:02:32.59" />
                    <SPLIT distance="250" swimtime="00:03:16.23" />
                    <SPLIT distance="300" swimtime="00:04:01.40" />
                    <SPLIT distance="350" swimtime="00:04:48.20" />
                    <SPLIT distance="400" swimtime="00:05:37.82" />
                    <SPLIT distance="450" swimtime="00:06:28.72" />
                    <SPLIT distance="500" swimtime="00:07:18.48" />
                    <SPLIT distance="550" swimtime="00:08:07.11" />
                    <SPLIT distance="600" swimtime="00:08:58.54" />
                    <SPLIT distance="650" swimtime="00:09:49.33" />
                    <SPLIT distance="700" swimtime="00:10:41.04" />
                    <SPLIT distance="750" swimtime="00:11:31.27" />
                    <SPLIT distance="800" swimtime="00:12:23.02" />
                    <SPLIT distance="850" swimtime="00:13:13.69" />
                    <SPLIT distance="900" swimtime="00:14:05.10" />
                    <SPLIT distance="950" swimtime="00:14:57.11" />
                    <SPLIT distance="1000" swimtime="00:15:48.76" />
                    <SPLIT distance="1050" swimtime="00:16:41.50" />
                    <SPLIT distance="1100" swimtime="00:17:34.30" />
                    <SPLIT distance="1150" swimtime="00:18:26.47" />
                    <SPLIT distance="1200" swimtime="00:19:20.18" />
                    <SPLIT distance="1250" swimtime="00:20:12.51" />
                    <SPLIT distance="1300" swimtime="00:21:03.15" />
                    <SPLIT distance="1350" swimtime="00:21:54.86" />
                    <SPLIT distance="1400" swimtime="00:22:47.55" />
                    <SPLIT distance="1450" swimtime="00:23:38.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="327" swimtime="00:05:37.71" resultid="1567" heatid="2188" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:01:17.98" />
                    <SPLIT distance="150" swimtime="00:01:56.91" />
                    <SPLIT distance="200" swimtime="00:02:37.06" />
                    <SPLIT distance="250" swimtime="00:03:20.14" />
                    <SPLIT distance="300" swimtime="00:04:03.93" />
                    <SPLIT distance="350" swimtime="00:04:51.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1381" points="317" swimtime="00:11:55.35" resultid="1568" heatid="2213" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                    <SPLIT distance="100" swimtime="00:01:15.37" />
                    <SPLIT distance="150" swimtime="00:01:57.05" />
                    <SPLIT distance="200" swimtime="00:02:39.73" />
                    <SPLIT distance="250" swimtime="00:03:23.97" />
                    <SPLIT distance="300" swimtime="00:04:10.12" />
                    <SPLIT distance="350" swimtime="00:04:55.67" />
                    <SPLIT distance="400" swimtime="00:05:42.06" />
                    <SPLIT distance="450" swimtime="00:06:28.57" />
                    <SPLIT distance="500" swimtime="00:07:15.50" />
                    <SPLIT distance="550" swimtime="00:08:03.16" />
                    <SPLIT distance="600" swimtime="00:08:51.40" />
                    <SPLIT distance="650" swimtime="00:09:41.03" />
                    <SPLIT distance="700" swimtime="00:10:28.13" />
                    <SPLIT distance="750" swimtime="00:11:14.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Luiza Sacramento" birthdate="2004-06-27" gender="F" nation="BRA" license="V413249" athleteid="1593" externalid="V413249">
              <RESULTS>
                <RESULT eventid="1113" points="205" swimtime="00:00:47.21" resultid="1594" heatid="2161" lane="2" />
                <RESULT eventid="1273" points="316" swimtime="00:00:36.70" resultid="1595" heatid="2195" lane="2" />
                <RESULT eventid="1394" points="184" swimtime="00:01:46.43" resultid="1596" heatid="2215" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luan" lastname="Schwarzbach Paula" birthdate="2005-07-29" gender="M" nation="BRA" license="358250" swrid="5622305" athleteid="1581" externalid="358250">
              <RESULTS>
                <RESULT eventid="1260" points="396" swimtime="00:02:53.69" resultid="1582" heatid="2194" lane="5" entrytime="00:02:47.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                    <SPLIT distance="100" swimtime="00:01:20.93" />
                    <SPLIT distance="150" swimtime="00:02:06.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1485" points="407" swimtime="00:01:18.45" resultid="1583" heatid="2232" lane="5" entrytime="00:01:18.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="419" swimtime="00:02:20.15" resultid="1584" heatid="2223" lane="2" entrytime="00:02:14.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                    <SPLIT distance="100" swimtime="00:01:07.48" />
                    <SPLIT distance="150" swimtime="00:01:43.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrielly" lastname="Rebbeka Silva" birthdate="2002-08-30" gender="F" nation="BRA" license="V413251" athleteid="1601" externalid="V413251">
              <RESULTS>
                <RESULT eventid="1113" points="301" swimtime="00:00:41.60" resultid="1602" heatid="2160" lane="2" />
                <RESULT eventid="1498" points="199" swimtime="00:28:23.96" resultid="1603" heatid="2234" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.41" />
                    <SPLIT distance="100" swimtime="00:01:35.34" />
                    <SPLIT distance="150" swimtime="00:02:27.86" />
                    <SPLIT distance="200" swimtime="00:03:23.35" />
                    <SPLIT distance="250" swimtime="00:04:18.78" />
                    <SPLIT distance="300" swimtime="00:05:15.43" />
                    <SPLIT distance="350" swimtime="00:06:12.52" />
                    <SPLIT distance="400" swimtime="00:07:10.15" />
                    <SPLIT distance="450" swimtime="00:08:07.38" />
                    <SPLIT distance="500" swimtime="00:09:05.30" />
                    <SPLIT distance="550" swimtime="00:10:03.82" />
                    <SPLIT distance="600" swimtime="00:11:03.75" />
                    <SPLIT distance="650" swimtime="00:12:04.56" />
                    <SPLIT distance="700" swimtime="00:13:00.01" />
                    <SPLIT distance="750" swimtime="00:13:56.37" />
                    <SPLIT distance="800" swimtime="00:14:52.32" />
                    <SPLIT distance="850" swimtime="00:15:49.98" />
                    <SPLIT distance="900" swimtime="00:16:48.90" />
                    <SPLIT distance="950" swimtime="00:17:47.73" />
                    <SPLIT distance="1000" swimtime="00:18:48.37" />
                    <SPLIT distance="1050" swimtime="00:19:46.70" />
                    <SPLIT distance="1100" swimtime="00:20:45.99" />
                    <SPLIT distance="1150" swimtime="00:21:44.29" />
                    <SPLIT distance="1200" swimtime="00:22:45.55" />
                    <SPLIT distance="1250" swimtime="00:23:45.17" />
                    <SPLIT distance="1300" swimtime="00:24:42.48" />
                    <SPLIT distance="1350" swimtime="00:25:39.98" />
                    <SPLIT distance="1400" swimtime="00:26:37.93" />
                    <SPLIT distance="1450" swimtime="00:27:35.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcos" lastname="Vinicius Bontorin" birthdate="2002-10-13" gender="M" nation="BRA" license="280586" athleteid="1533" externalid="280586">
              <RESULTS>
                <RESULT eventid="1152" points="276" swimtime="00:02:54.52" resultid="1534" heatid="2170" lane="3" entrytime="00:02:39.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                    <SPLIT distance="100" swimtime="00:01:16.05" />
                    <SPLIT distance="150" swimtime="00:02:04.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="373" swimtime="00:02:45.13" resultid="1535" heatid="2155" lane="4" entrytime="00:02:39.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                    <SPLIT distance="100" swimtime="00:01:14.49" />
                    <SPLIT distance="150" swimtime="00:02:02.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="394" swimtime="00:01:10.05" resultid="1536" heatid="2206" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Boff Da Silva" birthdate="2006-09-23" gender="F" nation="BRA" license="V413250" athleteid="1597" externalid="V413250">
              <RESULTS>
                <RESULT eventid="1139" points="412" swimtime="00:01:13.13" resultid="1598" heatid="2168" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="294" swimtime="00:00:45.83" resultid="1599" heatid="2177" lane="4" />
                <RESULT eventid="1299" points="288" swimtime="00:03:17.30" resultid="1600" heatid="2202" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                    <SPLIT distance="100" swimtime="00:01:31.91" />
                    <SPLIT distance="150" swimtime="00:02:25.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Schlickmann Assis" birthdate="2003-07-24" gender="F" nation="BRA" license="303874" swrid="5600257" athleteid="1537" externalid="303874">
              <RESULTS>
                <RESULT eventid="1087" points="651" swimtime="00:02:38.27" resultid="1538" heatid="2156" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:15.88" />
                    <SPLIT distance="150" swimtime="00:01:58.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="604" swimtime="00:00:29.56" resultid="1539" heatid="2197" lane="4" entrytime="00:00:29.69" entrycourse="SCM" />
                <RESULT eventid="1472" points="611" swimtime="00:01:18.74" resultid="1540" heatid="2229" lane="3" entrytime="00:01:15.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Kuwaki" birthdate="1990-07-02" gender="M" nation="BRA" license="267975" athleteid="1553" externalid="267975">
              <RESULTS>
                <RESULT eventid="1178" points="783" swimtime="00:00:28.98" resultid="1554" heatid="2176" lane="3" entrytime="00:00:28.88" entrycourse="SCM" />
                <RESULT eventid="1286" points="814" swimtime="00:00:23.05" resultid="1555" heatid="2201" lane="4" entrytime="00:00:23.82" entrycourse="SCM" />
                <RESULT eventid="1459" points="741" swimtime="00:00:25.27" resultid="1556" heatid="2227" lane="4" entrytime="00:00:25.41" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rodrigo" lastname="Rieping" birthdate="1989-11-03" gender="M" nation="BRA" license="V413222" athleteid="1541" externalid="V413222">
              <RESULTS>
                <RESULT eventid="1204" points="445" swimtime="00:20:32.66" resultid="1542" heatid="2181" lane="2" entrytime="00:19:26.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="100" swimtime="00:01:04.35" />
                    <SPLIT distance="150" swimtime="00:01:39.24" />
                    <SPLIT distance="200" swimtime="00:02:16.54" />
                    <SPLIT distance="250" swimtime="00:02:55.44" />
                    <SPLIT distance="300" swimtime="00:03:34.72" />
                    <SPLIT distance="350" swimtime="00:04:15.41" />
                    <SPLIT distance="400" swimtime="00:04:55.13" />
                    <SPLIT distance="450" swimtime="00:05:35.95" />
                    <SPLIT distance="500" swimtime="00:06:18.12" />
                    <SPLIT distance="550" swimtime="00:07:00.07" />
                    <SPLIT distance="600" swimtime="00:07:43.95" />
                    <SPLIT distance="650" swimtime="00:08:29.21" />
                    <SPLIT distance="700" swimtime="00:09:13.17" />
                    <SPLIT distance="750" swimtime="00:09:56.35" />
                    <SPLIT distance="800" swimtime="00:10:39.66" />
                    <SPLIT distance="850" swimtime="00:11:23.11" />
                    <SPLIT distance="900" swimtime="00:12:06.46" />
                    <SPLIT distance="950" swimtime="00:12:49.11" />
                    <SPLIT distance="1000" swimtime="00:13:32.74" />
                    <SPLIT distance="1050" swimtime="00:14:15.09" />
                    <SPLIT distance="1100" swimtime="00:14:57.48" />
                    <SPLIT distance="1150" swimtime="00:15:39.69" />
                    <SPLIT distance="1200" swimtime="00:16:22.47" />
                    <SPLIT distance="1250" swimtime="00:17:05.21" />
                    <SPLIT distance="1300" swimtime="00:17:47.86" />
                    <SPLIT distance="1350" swimtime="00:18:29.88" />
                    <SPLIT distance="1400" swimtime="00:19:12.07" />
                    <SPLIT distance="1450" swimtime="00:19:52.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="588" swimtime="00:04:43.66" resultid="1543" heatid="2189" lane="4" entrytime="00:04:48.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="100" swimtime="00:01:07.82" />
                    <SPLIT distance="150" swimtime="00:01:43.18" />
                    <SPLIT distance="200" swimtime="00:02:19.42" />
                    <SPLIT distance="250" swimtime="00:02:56.06" />
                    <SPLIT distance="300" swimtime="00:03:33.38" />
                    <SPLIT distance="350" swimtime="00:04:09.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1381" points="523" swimtime="00:10:15.63" resultid="1544" heatid="2214" lane="4" entrytime="00:10:07.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:10.01" />
                    <SPLIT distance="150" swimtime="00:01:46.74" />
                    <SPLIT distance="200" swimtime="00:02:24.47" />
                    <SPLIT distance="250" swimtime="00:03:02.71" />
                    <SPLIT distance="300" swimtime="00:03:41.48" />
                    <SPLIT distance="350" swimtime="00:04:20.68" />
                    <SPLIT distance="400" swimtime="00:04:59.81" />
                    <SPLIT distance="450" swimtime="00:05:39.01" />
                    <SPLIT distance="500" swimtime="00:06:19.22" />
                    <SPLIT distance="550" swimtime="00:06:59.28" />
                    <SPLIT distance="600" swimtime="00:07:39.38" />
                    <SPLIT distance="650" swimtime="00:08:19.96" />
                    <SPLIT distance="700" swimtime="00:08:59.90" />
                    <SPLIT distance="750" swimtime="00:09:39.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marilia" lastname="Cato Oliveira" birthdate="2002-10-30" gender="F" nation="BRA" license="V383072" athleteid="1569" externalid="V383072">
              <RESULTS>
                <RESULT eventid="1113" points="645" swimtime="00:00:32.26" resultid="1570" heatid="2162" lane="3" entrytime="00:00:32.60" entrycourse="SCM" />
                <RESULT eventid="1394" points="614" swimtime="00:01:11.33" resultid="1571" heatid="2216" lane="4" entrytime="00:01:12.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1446" points="554" swimtime="00:00:31.81" resultid="1572" heatid="2224" lane="4" entrytime="00:00:32.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Carvalho Rodrigues" birthdate="2004-01-17" gender="F" nation="BRA" license="V249307" athleteid="1557" externalid="V249307">
              <RESULTS>
                <RESULT eventid="1191" points="399" swimtime="00:00:41.42" resultid="1558" heatid="2178" lane="4" entrytime="00:00:41.47" entrycourse="SCM" />
                <RESULT eventid="1247" points="372" swimtime="00:03:26.19" resultid="1559" heatid="2191" lane="4" entrytime="00:03:21.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.80" />
                    <SPLIT distance="100" swimtime="00:01:36.81" />
                    <SPLIT distance="150" swimtime="00:02:31.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1472" points="362" swimtime="00:01:33.74" resultid="1560" heatid="2229" lane="2" entrytime="00:01:33.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Brassac Kniggendorf" birthdate="2002-09-18" gender="F" nation="BRA" license="282706" athleteid="1585" externalid="282706">
              <RESULTS>
                <RESULT eventid="1139" points="414" swimtime="00:01:13.01" resultid="1586" heatid="2169" lane="5" entrytime="00:01:13.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1325" points="268" swimtime="00:01:30.02" resultid="1587" heatid="2205" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="484" swimtime="00:00:31.84" resultid="1588" heatid="2197" lane="5" entrytime="00:00:32.23" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andryws" lastname="Farinhuka" birthdate="2004-03-10" gender="M" nation="BRA" license="V285246" athleteid="1573" externalid="V285246">
              <RESULTS>
                <RESULT eventid="1074" points="359" swimtime="00:02:47.27" resultid="1574" heatid="2153" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="100" swimtime="00:01:16.57" />
                    <SPLIT distance="150" swimtime="00:02:07.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="378" swimtime="00:05:21.79" resultid="1575" heatid="2188" lane="2" entrytime="00:05:31.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                    <SPLIT distance="100" swimtime="00:01:14.11" />
                    <SPLIT distance="150" swimtime="00:01:54.51" />
                    <SPLIT distance="200" swimtime="00:02:36.79" />
                    <SPLIT distance="250" swimtime="00:03:20.84" />
                    <SPLIT distance="300" swimtime="00:04:04.91" />
                    <SPLIT distance="350" swimtime="00:04:47.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="377" swimtime="00:02:25.19" resultid="1576" heatid="2222" lane="3" entrytime="00:02:29.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.74" />
                    <SPLIT distance="100" swimtime="00:01:04.51" />
                    <SPLIT distance="150" swimtime="00:01:44.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Fagundes" birthdate="2002-06-02" gender="M" nation="BRA" license="331902" athleteid="1589" externalid="331902">
              <RESULTS>
                <RESULT eventid="1100" status="WDR" swimtime="00:00:00.00" resultid="1590" />
                <RESULT eventid="1312" status="WDR" swimtime="00:00:00.00" resultid="1591" />
                <RESULT eventid="1407" status="WDR" swimtime="00:00:00.00" resultid="1592" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Letícia" lastname="Ramos Souza" birthdate="2002-01-03" gender="F" nation="BRA" license="266069" athleteid="1545" externalid="266069">
              <RESULTS>
                <RESULT eventid="1061" points="311" swimtime="00:13:03.40" resultid="1546" heatid="2151" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                    <SPLIT distance="100" swimtime="00:01:18.97" />
                    <SPLIT distance="150" swimtime="00:02:04.06" />
                    <SPLIT distance="200" swimtime="00:02:50.19" />
                    <SPLIT distance="250" swimtime="00:03:38.67" />
                    <SPLIT distance="300" swimtime="00:04:29.70" />
                    <SPLIT distance="350" swimtime="00:05:20.18" />
                    <SPLIT distance="400" swimtime="00:06:11.01" />
                    <SPLIT distance="450" swimtime="00:07:02.41" />
                    <SPLIT distance="500" swimtime="00:07:52.21" />
                    <SPLIT distance="550" swimtime="00:08:43.98" />
                    <SPLIT distance="600" swimtime="00:09:35.70" />
                    <SPLIT distance="650" swimtime="00:10:28.06" />
                    <SPLIT distance="700" swimtime="00:11:20.15" />
                    <SPLIT distance="750" swimtime="00:12:11.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1221" points="327" swimtime="00:06:08.22" resultid="1547" heatid="2185" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:21.63" />
                    <SPLIT distance="150" swimtime="00:02:06.41" />
                    <SPLIT distance="200" swimtime="00:02:53.31" />
                    <SPLIT distance="250" swimtime="00:03:41.38" />
                    <SPLIT distance="300" swimtime="00:04:30.06" />
                    <SPLIT distance="350" swimtime="00:05:20.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1394" points="348" swimtime="00:01:26.17" resultid="1548" heatid="2215" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="PUCPR (CURITIBA) &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1219" swimtime="00:03:38.66" resultid="1607" heatid="2184" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.81" />
                    <SPLIT distance="100" swimtime="00:00:59.40" />
                    <SPLIT distance="150" swimtime="00:01:24.47" />
                    <SPLIT distance="200" swimtime="00:01:53.49" />
                    <SPLIT distance="250" swimtime="00:02:18.64" />
                    <SPLIT distance="300" swimtime="00:02:46.25" />
                    <SPLIT distance="350" swimtime="00:03:09.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1577" number="1" />
                    <RELAYPOSITION athleteid="1561" number="2" />
                    <RELAYPOSITION athleteid="1549" number="3" />
                    <RELAYPOSITION athleteid="1553" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1379" swimtime="00:09:02.62" resultid="1608" heatid="2212" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.55" />
                    <SPLIT distance="100" swimtime="00:01:01.58" />
                    <SPLIT distance="150" swimtime="00:01:35.36" />
                    <SPLIT distance="200" swimtime="00:02:10.68" />
                    <SPLIT distance="250" swimtime="00:02:42.78" />
                    <SPLIT distance="300" swimtime="00:03:19.35" />
                    <SPLIT distance="350" swimtime="00:03:56.52" />
                    <SPLIT distance="400" swimtime="00:04:31.53" />
                    <SPLIT distance="450" swimtime="00:05:03.42" />
                    <SPLIT distance="500" swimtime="00:05:39.07" />
                    <SPLIT distance="550" swimtime="00:06:15.88" />
                    <SPLIT distance="600" swimtime="00:06:52.02" />
                    <SPLIT distance="650" swimtime="00:07:21.00" />
                    <SPLIT distance="700" swimtime="00:07:54.14" />
                    <SPLIT distance="750" swimtime="00:08:27.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1541" number="1" />
                    <RELAYPOSITION athleteid="1549" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1581" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1561" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" swimtime="00:04:17.98" resultid="1609" heatid="2236" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                    <SPLIT distance="100" swimtime="00:01:03.51" />
                    <SPLIT distance="150" swimtime="00:01:35.34" />
                    <SPLIT distance="200" swimtime="00:02:11.13" />
                    <SPLIT distance="250" swimtime="00:02:40.47" />
                    <SPLIT distance="300" swimtime="00:03:16.34" />
                    <SPLIT distance="350" swimtime="00:03:44.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1549" number="1" />
                    <RELAYPOSITION athleteid="1553" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1561" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1573" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="PUCPR (CURITIBA) &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1217" swimtime="00:04:34.89" resultid="1604" heatid="2182" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                    <SPLIT distance="100" swimtime="00:01:12.11" />
                    <SPLIT distance="150" swimtime="00:01:46.32" />
                    <SPLIT distance="200" swimtime="00:02:26.24" />
                    <SPLIT distance="250" swimtime="00:02:56.84" />
                    <SPLIT distance="300" swimtime="00:03:31.36" />
                    <SPLIT distance="350" swimtime="00:04:01.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1545" number="1" />
                    <RELAYPOSITION athleteid="1557" number="2" />
                    <RELAYPOSITION athleteid="1569" number="3" />
                    <RELAYPOSITION athleteid="1537" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1377" swimtime="00:10:56.58" resultid="1605" heatid="2211" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:18.33" />
                    <SPLIT distance="150" swimtime="00:02:04.22" />
                    <SPLIT distance="200" swimtime="00:02:53.14" />
                    <SPLIT distance="250" swimtime="00:03:32.21" />
                    <SPLIT distance="300" swimtime="00:04:15.92" />
                    <SPLIT distance="350" swimtime="00:05:02.47" />
                    <SPLIT distance="400" swimtime="00:05:47.96" />
                    <SPLIT distance="450" swimtime="00:06:22.60" />
                    <SPLIT distance="500" swimtime="00:07:01.00" />
                    <SPLIT distance="550" swimtime="00:07:41.44" />
                    <SPLIT distance="600" swimtime="00:08:22.93" />
                    <SPLIT distance="650" swimtime="00:08:58.93" />
                    <SPLIT distance="700" swimtime="00:09:38.73" />
                    <SPLIT distance="750" swimtime="00:10:17.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1545" number="1" />
                    <RELAYPOSITION athleteid="1557" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1569" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1537" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1513" swimtime="00:05:15.87" resultid="1606" heatid="2237" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="100" swimtime="00:01:27.55" />
                    <SPLIT distance="150" swimtime="00:02:03.80" />
                    <SPLIT distance="200" swimtime="00:02:45.27" />
                    <SPLIT distance="250" swimtime="00:03:19.81" />
                    <SPLIT distance="300" swimtime="00:04:03.92" />
                    <SPLIT distance="350" swimtime="00:04:36.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1545" number="1" />
                    <RELAYPOSITION athleteid="1537" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1569" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1585" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="16614" nation="BRA" region="PR" clubid="1516" name="Fag (Cascavel)">
          <ATHLETES>
            <ATHLETE firstname="Gustavo" lastname="Henrique Wiebbeling" birthdate="2003-08-06" gender="M" nation="BRA" license="290420" swrid="4471225" athleteid="1517" externalid="290420">
              <RESULTS>
                <RESULT eventid="1204" points="638" swimtime="00:17:59.71" resultid="1518" heatid="2181" lane="3" entrytime="00:17:34.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                    <SPLIT distance="100" swimtime="00:01:03.76" />
                    <SPLIT distance="150" swimtime="00:01:37.70" />
                    <SPLIT distance="200" swimtime="00:02:12.37" />
                    <SPLIT distance="250" swimtime="00:02:47.51" />
                    <SPLIT distance="300" swimtime="00:03:22.74" />
                    <SPLIT distance="350" swimtime="00:03:58.55" />
                    <SPLIT distance="400" swimtime="00:04:34.66" />
                    <SPLIT distance="450" swimtime="00:05:10.81" />
                    <SPLIT distance="500" swimtime="00:05:47.18" />
                    <SPLIT distance="550" swimtime="00:06:23.94" />
                    <SPLIT distance="600" swimtime="00:07:00.17" />
                    <SPLIT distance="650" swimtime="00:07:36.68" />
                    <SPLIT distance="700" swimtime="00:08:13.03" />
                    <SPLIT distance="750" swimtime="00:08:49.69" />
                    <SPLIT distance="800" swimtime="00:09:26.57" />
                    <SPLIT distance="850" swimtime="00:10:03.52" />
                    <SPLIT distance="900" swimtime="00:10:40.31" />
                    <SPLIT distance="950" swimtime="00:11:16.87" />
                    <SPLIT distance="1000" swimtime="00:11:53.94" />
                    <SPLIT distance="1050" swimtime="00:12:30.73" />
                    <SPLIT distance="1100" swimtime="00:13:07.83" />
                    <SPLIT distance="1150" swimtime="00:13:44.58" />
                    <SPLIT distance="1200" swimtime="00:14:20.96" />
                    <SPLIT distance="1250" swimtime="00:14:57.90" />
                    <SPLIT distance="1300" swimtime="00:15:34.49" />
                    <SPLIT distance="1350" swimtime="00:16:11.50" />
                    <SPLIT distance="1400" swimtime="00:16:48.70" />
                    <SPLIT distance="1450" swimtime="00:17:25.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" status="DNS" swimtime="00:00:00.00" resultid="1519" heatid="2204" lane="4" entrytime="00:02:17.43" entrycourse="SCM" />
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="1520" heatid="2187" lane="2" entrytime="00:04:21.56" entrycourse="SCM" />
                <RESULT eventid="1381" status="DNS" swimtime="00:00:00.00" resultid="1521" heatid="2214" lane="3" entrytime="00:09:03.49" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6489" nation="BRA" region="PR" clubid="1725" name="Ufpr (Curitiba)">
          <ATHLETES>
            <ATHLETE firstname="Isabella" lastname="Coelho Gentil" birthdate="2003-08-14" gender="F" nation="BRA" license="250061" athleteid="1750" externalid="250061">
              <RESULTS>
                <RESULT eventid="1299" points="461" swimtime="00:02:48.72" resultid="1751" heatid="2202" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.02" />
                    <SPLIT distance="100" swimtime="00:01:21.97" />
                    <SPLIT distance="150" swimtime="00:02:05.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1221" points="409" swimtime="00:05:41.72" resultid="1752" heatid="2185" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:14.00" />
                    <SPLIT distance="150" swimtime="00:01:54.32" />
                    <SPLIT distance="200" swimtime="00:02:36.78" />
                    <SPLIT distance="250" swimtime="00:03:21.97" />
                    <SPLIT distance="300" swimtime="00:04:07.58" />
                    <SPLIT distance="350" swimtime="00:04:54.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1394" points="488" swimtime="00:01:16.97" resultid="1753" heatid="2215" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Jose Ferrarini" birthdate="1999-01-31" gender="M" nation="BRA" license="151451" athleteid="1779" externalid="151451">
              <RESULTS>
                <RESULT eventid="1126" points="317" swimtime="00:01:09.51" resultid="1780" heatid="2164" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="297" swimtime="00:00:35.49" resultid="1781" heatid="2158" lane="2" />
                <RESULT eventid="1407" points="308" swimtime="00:01:17.02" resultid="1782" heatid="2217" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Adelaide" lastname="Ely Tigrinho" birthdate="2004-05-17" gender="F" nation="BRA" license="315043" athleteid="1737" externalid="315043">
              <RESULTS>
                <RESULT eventid="1139" points="352" swimtime="00:01:17.08" resultid="1738" heatid="2168" lane="3" entrytime="00:01:20.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="402" swimtime="00:00:41.30" resultid="1739" heatid="2178" lane="5" entrytime="00:00:43.47" entrycourse="SCM" />
                <RESULT eventid="1273" points="397" swimtime="00:00:34.00" resultid="1740" heatid="2196" lane="3" entrytime="00:00:33.88" entrycourse="SCM" />
                <RESULT eventid="1472" points="313" swimtime="00:01:38.33" resultid="1741" heatid="2228" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Friedrich Jakobi" birthdate="2004-02-10" gender="M" nation="BRA" license="V413275" athleteid="1768" externalid="V413275">
              <RESULTS>
                <RESULT eventid="1126" points="417" swimtime="00:01:03.47" resultid="1769" heatid="2165" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1338" points="386" swimtime="00:01:10.52" resultid="1770" heatid="2206" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="459" swimtime="00:00:27.58" resultid="1771" heatid="2198" lane="3" />
                <RESULT eventid="1459" points="459" swimtime="00:00:30.01" resultid="1772" heatid="2225" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kathierry" lastname="Lazarin Wolff" birthdate="2005-03-18" gender="F" nation="BRA" license="V307778" athleteid="1773" externalid="V307778">
              <RESULTS>
                <RESULT eventid="1139" points="174" swimtime="00:01:37.42" resultid="1774" heatid="2168" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="187" swimtime="00:00:48.72" resultid="1775" heatid="2161" lane="5" />
                <RESULT eventid="1191" points="210" swimtime="00:00:51.29" resultid="1776" heatid="2177" lane="5" />
                <RESULT eventid="1247" status="DSQ" swimtime="00:04:19.61" resultid="1777" heatid="2190" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.48" />
                    <SPLIT distance="100" swimtime="00:01:56.46" />
                    <SPLIT distance="150" swimtime="00:03:08.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="211" swimtime="00:00:41.97" resultid="1778" heatid="2196" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natan" lastname="Romão Freire" birthdate="2000-07-13" gender="M" nation="BRA" license="273578" athleteid="1754" externalid="273578">
              <RESULTS>
                <RESULT eventid="1178" points="572" swimtime="00:00:32.51" resultid="1755" heatid="2173" lane="2" />
                <RESULT eventid="1286" points="527" swimtime="00:00:26.34" resultid="1756" heatid="2199" lane="2" />
                <RESULT eventid="1485" points="512" swimtime="00:01:12.65" resultid="1757" heatid="2230" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Maria Ramos" birthdate="2002-03-09" gender="F" nation="BRA" license="V413200" athleteid="1742" externalid="V413200">
              <RESULTS>
                <RESULT eventid="1165" points="186" swimtime="00:03:46.98" resultid="1743" heatid="2172" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.81" />
                    <SPLIT distance="100" swimtime="00:01:45.75" />
                    <SPLIT distance="150" swimtime="00:02:45.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1061" points="254" swimtime="00:13:58.23" resultid="1744" heatid="2151" lane="3" entrytime="00:14:07.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.63" />
                    <SPLIT distance="100" swimtime="00:01:36.12" />
                    <SPLIT distance="150" swimtime="00:02:27.83" />
                    <SPLIT distance="200" swimtime="00:03:20.80" />
                    <SPLIT distance="250" swimtime="00:04:13.57" />
                    <SPLIT distance="300" swimtime="00:05:07.00" />
                    <SPLIT distance="350" swimtime="00:06:00.52" />
                    <SPLIT distance="400" swimtime="00:06:54.40" />
                    <SPLIT distance="450" swimtime="00:07:47.89" />
                    <SPLIT distance="500" swimtime="00:08:42.03" />
                    <SPLIT distance="550" swimtime="00:09:36.06" />
                    <SPLIT distance="600" swimtime="00:10:29.74" />
                    <SPLIT distance="650" swimtime="00:11:23.42" />
                    <SPLIT distance="700" swimtime="00:12:17.50" />
                    <SPLIT distance="750" swimtime="00:13:09.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1498" points="235" swimtime="00:26:52.45" resultid="1745" heatid="2234" lane="1" entrytime="00:27:12.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.85" />
                    <SPLIT distance="100" swimtime="00:01:33.09" />
                    <SPLIT distance="150" swimtime="00:02:24.73" />
                    <SPLIT distance="200" swimtime="00:03:17.12" />
                    <SPLIT distance="250" swimtime="00:04:10.51" />
                    <SPLIT distance="300" swimtime="00:05:04.43" />
                    <SPLIT distance="350" swimtime="00:05:58.43" />
                    <SPLIT distance="400" swimtime="00:06:52.65" />
                    <SPLIT distance="450" swimtime="00:07:46.89" />
                    <SPLIT distance="500" swimtime="00:08:40.69" />
                    <SPLIT distance="550" swimtime="00:09:35.03" />
                    <SPLIT distance="600" swimtime="00:10:29.40" />
                    <SPLIT distance="650" swimtime="00:11:24.21" />
                    <SPLIT distance="700" swimtime="00:12:18.34" />
                    <SPLIT distance="750" swimtime="00:13:12.29" />
                    <SPLIT distance="800" swimtime="00:14:06.89" />
                    <SPLIT distance="850" swimtime="00:15:01.29" />
                    <SPLIT distance="900" swimtime="00:15:56.44" />
                    <SPLIT distance="950" swimtime="00:16:50.76" />
                    <SPLIT distance="1000" swimtime="00:17:45.77" />
                    <SPLIT distance="1050" swimtime="00:18:41.08" />
                    <SPLIT distance="1100" swimtime="00:19:36.32" />
                    <SPLIT distance="1150" swimtime="00:20:30.89" />
                    <SPLIT distance="1200" swimtime="00:21:25.13" />
                    <SPLIT distance="1250" swimtime="00:22:20.50" />
                    <SPLIT distance="1300" swimtime="00:23:15.53" />
                    <SPLIT distance="1350" swimtime="00:24:10.91" />
                    <SPLIT distance="1400" swimtime="00:25:05.51" />
                    <SPLIT distance="1450" swimtime="00:26:00.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="André" lastname="Cherbaty Filho" birthdate="2006-01-01" gender="M" nation="BRA" license="V285322" athleteid="1758" externalid="V285322">
              <RESULTS>
                <RESULT eventid="1459" status="DSQ" swimtime="00:00:33.26" resultid="1759" heatid="2225" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Caroleski" birthdate="2005-08-10" gender="M" nation="BRA" license="366980" swrid="5622266" athleteid="1732" externalid="366980">
              <RESULTS>
                <RESULT eventid="1126" points="417" swimtime="00:01:03.45" resultid="1733" heatid="2165" lane="3" entrytime="00:01:01.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="286" swimtime="00:00:35.93" resultid="1734" heatid="2158" lane="3" entrytime="00:00:33.24" entrycourse="SCM" />
                <RESULT eventid="1286" points="424" swimtime="00:00:28.32" resultid="1735" heatid="2200" lane="2" entrytime="00:00:27.57" entrycourse="SCM" />
                <RESULT eventid="1459" points="376" swimtime="00:00:32.05" resultid="1736" heatid="2226" lane="3" entrytime="00:00:29.68" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karolyne" lastname="Magario Hayashi" birthdate="2001-03-19" gender="F" nation="BRA" license="V413272" athleteid="1760" externalid="V413272">
              <RESULTS>
                <RESULT eventid="1191" points="461" swimtime="00:00:39.46" resultid="1761" heatid="2177" lane="2" />
                <RESULT eventid="1247" points="475" swimtime="00:03:10.05" resultid="1762" heatid="2191" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.12" />
                    <SPLIT distance="100" swimtime="00:01:29.86" />
                    <SPLIT distance="150" swimtime="00:02:18.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="501" swimtime="00:00:31.46" resultid="1763" heatid="2195" lane="4" />
                <RESULT eventid="1472" points="453" swimtime="00:01:27.00" resultid="1764" heatid="2228" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Pivetta Caldana" birthdate="2005-04-16" gender="F" nation="BRA" license="V413273" athleteid="1765" externalid="V413273">
              <RESULTS>
                <RESULT eventid="1139" status="WDR" swimtime="00:00:00.00" resultid="1766" heatid="2167" lane="2" />
                <RESULT eventid="1113" status="WDR" swimtime="00:00:00.00" resultid="1767" heatid="2161" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Barros Zagonel" birthdate="2006-06-01" gender="M" nation="BRA" license="347856" swrid="5622261" athleteid="1726" externalid="347856">
              <RESULTS>
                <RESULT eventid="1074" points="369" swimtime="00:02:45.78" resultid="1727" heatid="2154" lane="3" entrytime="00:02:51.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                    <SPLIT distance="100" swimtime="00:01:19.30" />
                    <SPLIT distance="150" swimtime="00:02:09.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="406" swimtime="00:00:36.43" resultid="1728" heatid="2176" lane="1" entrytime="00:00:35.13" entrycourse="SCM" />
                <RESULT eventid="1260" points="326" swimtime="00:03:05.31" resultid="1729" heatid="2193" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                    <SPLIT distance="100" swimtime="00:01:27.86" />
                    <SPLIT distance="150" swimtime="00:02:17.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1485" points="338" swimtime="00:01:23.43" resultid="1730" heatid="2232" lane="1" entrytime="00:01:20.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1433" points="373" swimtime="00:02:25.71" resultid="1731" heatid="2221" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:09.89" />
                    <SPLIT distance="150" swimtime="00:01:49.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Erick" lastname="Eduardo Taner" birthdate="1999-05-31" gender="M" nation="BRA" license="V413212" athleteid="1746" externalid="V413212">
              <RESULTS>
                <RESULT eventid="1178" status="DNS" swimtime="00:00:00.00" resultid="1747" heatid="2175" lane="4" entrytime="00:00:41.19" entrycourse="SCM" />
                <RESULT eventid="1260" status="WDR" swimtime="00:00:00.00" resultid="1748" heatid="2192" lane="2" />
                <RESULT eventid="1485" status="WDR" swimtime="00:00:00.00" resultid="1749" heatid="2231" lane="4" entrytime="00:01:28.49" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="UFPR (CURITIBA) &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1219" swimtime="00:04:17.21" resultid="1786" heatid="2184" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                    <SPLIT distance="100" swimtime="00:01:04.50" />
                    <SPLIT distance="150" swimtime="00:01:35.06" />
                    <SPLIT distance="200" swimtime="00:02:13.72" />
                    <SPLIT distance="250" swimtime="00:02:44.22" />
                    <SPLIT distance="300" swimtime="00:03:19.06" />
                    <SPLIT distance="350" swimtime="00:03:46.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1732" number="1" />
                    <RELAYPOSITION athleteid="1758" number="2" />
                    <RELAYPOSITION athleteid="1726" number="3" />
                    <RELAYPOSITION athleteid="1754" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" swimtime="00:04:47.02" resultid="1787" heatid="2236" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.43" />
                    <SPLIT distance="100" swimtime="00:01:21.04" />
                    <SPLIT distance="150" swimtime="00:01:55.23" />
                    <SPLIT distance="200" swimtime="00:02:33.97" />
                    <SPLIT distance="250" swimtime="00:03:04.49" />
                    <SPLIT distance="300" swimtime="00:03:42.76" />
                    <SPLIT distance="350" swimtime="00:04:12.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1732" number="1" />
                    <RELAYPOSITION athleteid="1754" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1768" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1726" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="UFPR (CURITIBA) &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1217" swimtime="00:05:22.65" resultid="1783" heatid="2182" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                    <SPLIT distance="150" swimtime="00:01:49.40" />
                    <SPLIT distance="200" swimtime="00:02:32.43" />
                    <SPLIT distance="250" swimtime="00:03:11.83" />
                    <SPLIT distance="300" swimtime="00:04:07.38" />
                    <SPLIT distance="350" swimtime="00:04:42.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1760" number="1" />
                    <RELAYPOSITION athleteid="1737" number="2" />
                    <RELAYPOSITION athleteid="1773" number="3" />
                    <RELAYPOSITION athleteid="1750" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1377" swimtime="00:12:03.79" resultid="1784" heatid="2211" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="100" swimtime="00:01:25.91" />
                    <SPLIT distance="150" swimtime="00:02:15.82" />
                    <SPLIT distance="200" swimtime="00:03:07.04" />
                    <SPLIT distance="250" swimtime="00:03:49.18" />
                    <SPLIT distance="300" swimtime="00:04:35.85" />
                    <SPLIT distance="350" swimtime="00:05:24.89" />
                    <SPLIT distance="400" swimtime="00:06:11.38" />
                    <SPLIT distance="450" swimtime="00:06:50.88" />
                    <SPLIT distance="500" swimtime="00:07:35.73" />
                    <SPLIT distance="550" swimtime="00:08:20.39" />
                    <SPLIT distance="600" swimtime="00:09:04.67" />
                    <SPLIT distance="650" swimtime="00:09:46.17" />
                    <SPLIT distance="700" swimtime="00:10:31.66" />
                    <SPLIT distance="750" swimtime="00:11:17.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1737" number="1" />
                    <RELAYPOSITION athleteid="1742" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1760" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1750" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1513" swimtime="00:05:52.33" resultid="1785" heatid="2237" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                    <SPLIT distance="100" swimtime="00:01:20.23" />
                    <SPLIT distance="150" swimtime="00:02:01.54" />
                    <SPLIT distance="200" swimtime="00:02:50.15" />
                    <SPLIT distance="250" swimtime="00:03:39.74" />
                    <SPLIT distance="300" swimtime="00:04:36.58" />
                    <SPLIT distance="350" swimtime="00:05:11.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1750" number="1" />
                    <RELAYPOSITION athleteid="1760" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1742" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1737" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="10898" nation="BRA" region="PR" clubid="1925" name="Unioeste (Cascavel)">
          <ATHLETES>
            <ATHLETE firstname="Enzo" lastname="Valiente Rizzi" birthdate="2001-05-24" gender="M" nation="BRA" license="V304700" athleteid="1930" externalid="V304700">
              <RESULTS>
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="1931" heatid="2187" lane="3" />
                <RESULT eventid="1433" status="DNS" swimtime="00:00:00.00" resultid="1932" heatid="2221" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julio" lastname="Heck" birthdate="1998-02-15" gender="M" nation="BRA" license="185880" swrid="5596906" athleteid="1933" externalid="185880">
              <RESULTS>
                <RESULT eventid="1126" points="676" swimtime="00:00:54.03" resultid="1934" heatid="2166" lane="4" entrytime="00:00:52.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="440" swimtime="00:00:35.46" resultid="1935" heatid="2176" lane="5" entrytime="00:00:33.58" entrycourse="SCM" />
                <RESULT eventid="1286" points="690" swimtime="00:00:24.08" resultid="1936" heatid="2201" lane="3" entrytime="00:00:23.75" entrycourse="SCM" />
                <RESULT eventid="1459" status="DNS" swimtime="00:00:00.00" resultid="1937" heatid="2225" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="Mayumi  Novais" birthdate="2002-11-23" gender="F" nation="BRA" license="V134816" athleteid="1938" externalid="V134816">
              <RESULTS>
                <RESULT eventid="1139" points="206" swimtime="00:01:32.09" resultid="1939" heatid="2167" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="305" swimtime="00:00:41.40" resultid="1940" heatid="2161" lane="4" />
                <RESULT eventid="1273" status="DNS" swimtime="00:00:00.00" resultid="1941" heatid="2195" lane="1" />
                <RESULT eventid="1394" status="DNS" swimtime="00:00:00.00" resultid="1942" heatid="2215" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Andrade" birthdate="1999-10-06" gender="M" nation="BRA" license="V109962" athleteid="1926" externalid="V109962">
              <RESULTS>
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="1927" heatid="2154" lane="4" entrytime="00:02:57.51" entrycourse="SCM" />
                <RESULT eventid="1234" status="DNS" swimtime="00:00:00.00" resultid="1928" heatid="2187" lane="4" />
                <RESULT eventid="1433" status="DNS" swimtime="00:00:00.00" resultid="1929" heatid="2222" lane="2" entrytime="00:02:34.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6510" nation="BRA" region="PR" clubid="1943" name="Utfpr (Curitiba)">
          <ATHLETES>
            <ATHLETE firstname="Isabelle" lastname="Haygert" birthdate="2004-07-02" gender="F" nation="BRA" license="V325677" athleteid="1970" externalid="V325677">
              <RESULTS>
                <RESULT eventid="1139" points="361" swimtime="00:01:16.44" resultid="1971" heatid="2167" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="327" swimtime="00:00:44.27" resultid="1972" heatid="2178" lane="1" />
                <RESULT eventid="1221" points="293" swimtime="00:06:21.67" resultid="1973" heatid="2185" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:01:19.94" />
                    <SPLIT distance="150" swimtime="00:02:08.32" />
                    <SPLIT distance="200" swimtime="00:02:58.30" />
                    <SPLIT distance="250" swimtime="00:03:50.03" />
                    <SPLIT distance="300" swimtime="00:04:42.14" />
                    <SPLIT distance="350" swimtime="00:05:33.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1472" points="345" swimtime="00:01:35.24" resultid="1974" heatid="2228" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1420" points="297" swimtime="00:02:56.75" resultid="1975" heatid="2220" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                    <SPLIT distance="100" swimtime="00:01:23.45" />
                    <SPLIT distance="150" swimtime="00:02:11.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Paulo Ferreira" birthdate="2005-12-16" gender="M" nation="BRA" license="400266" swrid="5653300" athleteid="1981" externalid="400266">
              <RESULTS>
                <RESULT eventid="1126" points="246" swimtime="00:01:15.64" resultid="1982" heatid="2163" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="188" swimtime="00:03:27.31" resultid="1983" heatid="2153" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.26" />
                    <SPLIT distance="100" swimtime="00:01:32.99" />
                    <SPLIT distance="150" swimtime="00:02:31.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1178" points="225" swimtime="00:00:44.36" resultid="1984" heatid="2174" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Loane" lastname="Ady Chiareto Tigrinho" birthdate="2002-03-11" gender="F" nation="BRA" license="306752" athleteid="1959" externalid="306752">
              <RESULTS>
                <RESULT eventid="1061" points="363" swimtime="00:12:24.58" resultid="1960" heatid="2152" lane="5" entrytime="00:11:51.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                    <SPLIT distance="100" swimtime="00:01:21.45" />
                    <SPLIT distance="150" swimtime="00:02:06.44" />
                    <SPLIT distance="200" swimtime="00:02:52.26" />
                    <SPLIT distance="250" swimtime="00:03:39.76" />
                    <SPLIT distance="300" swimtime="00:04:27.09" />
                    <SPLIT distance="350" swimtime="00:05:14.85" />
                    <SPLIT distance="400" swimtime="00:06:02.70" />
                    <SPLIT distance="450" swimtime="00:06:50.78" />
                    <SPLIT distance="500" swimtime="00:07:38.13" />
                    <SPLIT distance="550" swimtime="00:08:26.23" />
                    <SPLIT distance="600" swimtime="00:09:14.61" />
                    <SPLIT distance="650" swimtime="00:10:02.69" />
                    <SPLIT distance="700" swimtime="00:10:50.82" />
                    <SPLIT distance="750" swimtime="00:11:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1221" points="360" swimtime="00:05:56.52" resultid="1961" heatid="2185" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                    <SPLIT distance="100" swimtime="00:01:21.11" />
                    <SPLIT distance="150" swimtime="00:02:05.48" />
                    <SPLIT distance="200" swimtime="00:02:51.57" />
                    <SPLIT distance="250" swimtime="00:03:38.07" />
                    <SPLIT distance="300" swimtime="00:04:24.29" />
                    <SPLIT distance="350" swimtime="00:05:10.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="358" swimtime="00:00:35.20" resultid="1962" heatid="2195" lane="5" />
                <RESULT eventid="1498" points="371" swimtime="00:23:05.26" resultid="1963" heatid="2234" lane="4" entrytime="00:23:06.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.58" />
                    <SPLIT distance="100" swimtime="00:01:24.04" />
                    <SPLIT distance="150" swimtime="00:02:08.49" />
                    <SPLIT distance="200" swimtime="00:02:54.20" />
                    <SPLIT distance="250" swimtime="00:03:40.22" />
                    <SPLIT distance="300" swimtime="00:04:26.70" />
                    <SPLIT distance="350" swimtime="00:05:13.52" />
                    <SPLIT distance="400" swimtime="00:05:59.94" />
                    <SPLIT distance="450" swimtime="00:06:46.68" />
                    <SPLIT distance="500" swimtime="00:07:33.14" />
                    <SPLIT distance="550" swimtime="00:08:20.46" />
                    <SPLIT distance="600" swimtime="00:09:07.10" />
                    <SPLIT distance="650" swimtime="00:09:54.03" />
                    <SPLIT distance="700" swimtime="00:10:41.00" />
                    <SPLIT distance="750" swimtime="00:11:27.87" />
                    <SPLIT distance="800" swimtime="00:12:14.74" />
                    <SPLIT distance="850" swimtime="00:13:01.50" />
                    <SPLIT distance="900" swimtime="00:13:48.15" />
                    <SPLIT distance="950" swimtime="00:14:35.42" />
                    <SPLIT distance="1000" swimtime="00:15:22.26" />
                    <SPLIT distance="1050" swimtime="00:16:09.06" />
                    <SPLIT distance="1100" swimtime="00:16:55.72" />
                    <SPLIT distance="1150" swimtime="00:17:42.28" />
                    <SPLIT distance="1200" swimtime="00:18:29.06" />
                    <SPLIT distance="1250" swimtime="00:19:16.51" />
                    <SPLIT distance="1300" swimtime="00:20:03.44" />
                    <SPLIT distance="1350" swimtime="00:20:49.77" />
                    <SPLIT distance="1400" swimtime="00:21:35.22" />
                    <SPLIT distance="1450" swimtime="00:22:20.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Gonçalves" birthdate="2000-04-17" gender="M" nation="BRA" license="V123198" athleteid="1944" externalid="V123198">
              <RESULTS>
                <RESULT eventid="1364" points="382" swimtime="00:05:50.73" resultid="1945" heatid="2209" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                    <SPLIT distance="100" swimtime="00:01:14.02" />
                    <SPLIT distance="150" swimtime="00:01:58.39" />
                    <SPLIT distance="200" swimtime="00:02:40.90" />
                    <SPLIT distance="250" swimtime="00:03:30.67" />
                    <SPLIT distance="300" swimtime="00:04:24.40" />
                    <SPLIT distance="350" swimtime="00:05:09.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="552" swimtime="00:00:25.93" resultid="1946" heatid="2199" lane="5" />
                <RESULT eventid="1433" points="482" swimtime="00:02:13.79" resultid="1947" heatid="2223" lane="5" entrytime="00:02:18.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:03.99" />
                    <SPLIT distance="150" swimtime="00:01:38.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="455" swimtime="00:00:30.81" resultid="2238" heatid="2158" lane="5" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Sant&apos; Anna" birthdate="2006-06-13" gender="M" nation="BRA" license="377059" swrid="5622303" athleteid="1948" externalid="377059">
              <RESULTS>
                <RESULT eventid="1126" points="370" swimtime="00:01:06.05" resultid="1949" heatid="2163" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="340" swimtime="00:00:33.93" resultid="1950" heatid="2158" lane="4" entrytime="00:00:33.35" entrycourse="SCM" />
                <RESULT eventid="1286" points="426" swimtime="00:00:28.27" resultid="1951" heatid="2200" lane="1" entrytime="00:00:28.13" entrycourse="SCM" />
                <RESULT eventid="1459" points="355" swimtime="00:00:32.69" resultid="1952" heatid="2226" lane="5" entrytime="00:00:32.16" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Fernanda Pinto" birthdate="2004-09-17" gender="F" nation="BRA" license="391144" swrid="5600157" athleteid="1976" externalid="391144">
              <RESULTS>
                <RESULT eventid="1139" points="390" swimtime="00:01:14.51" resultid="1977" heatid="2169" lane="1" entrytime="00:01:16.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1113" points="313" swimtime="00:00:41.06" resultid="1978" heatid="2162" lane="5" entrytime="00:00:42.10" entrycourse="SCM" />
                <RESULT eventid="1273" points="445" swimtime="00:00:32.73" resultid="1979" heatid="2197" lane="1" entrytime="00:00:33.80" entrycourse="SCM" />
                <RESULT eventid="1420" points="331" swimtime="00:02:50.42" resultid="1980" heatid="2220" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.97" />
                    <SPLIT distance="100" swimtime="00:01:23.10" />
                    <SPLIT distance="150" swimtime="00:02:07.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karine" lastname="Correa" birthdate="2002-08-01" gender="F" nation="BRA" license="385191" swrid="5600141" athleteid="1964" externalid="385191">
              <RESULTS>
                <RESULT eventid="1061" points="432" swimtime="00:11:42.46" resultid="1965" heatid="2152" lane="2" entrytime="00:11:19.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                    <SPLIT distance="100" swimtime="00:01:19.74" />
                    <SPLIT distance="150" swimtime="00:02:01.30" />
                    <SPLIT distance="200" swimtime="00:02:43.51" />
                    <SPLIT distance="250" swimtime="00:03:26.33" />
                    <SPLIT distance="300" swimtime="00:04:10.78" />
                    <SPLIT distance="350" swimtime="00:04:53.51" />
                    <SPLIT distance="400" swimtime="00:05:37.98" />
                    <SPLIT distance="450" swimtime="00:06:23.27" />
                    <SPLIT distance="500" swimtime="00:07:08.59" />
                    <SPLIT distance="550" swimtime="00:07:54.45" />
                    <SPLIT distance="600" swimtime="00:08:40.91" />
                    <SPLIT distance="650" swimtime="00:09:26.81" />
                    <SPLIT distance="700" swimtime="00:10:13.43" />
                    <SPLIT distance="750" swimtime="00:10:59.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1221" points="475" swimtime="00:05:25.04" resultid="1966" heatid="2186" lane="4" entrytime="00:05:35.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                    <SPLIT distance="100" swimtime="00:01:15.44" />
                    <SPLIT distance="150" swimtime="00:01:55.97" />
                    <SPLIT distance="200" swimtime="00:02:36.99" />
                    <SPLIT distance="250" swimtime="00:03:18.97" />
                    <SPLIT distance="300" swimtime="00:04:01.52" />
                    <SPLIT distance="350" swimtime="00:04:44.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1273" points="410" swimtime="00:00:33.64" resultid="1967" heatid="2196" lane="2" />
                <RESULT eventid="1498" points="402" swimtime="00:22:29.09" resultid="1968" heatid="2234" lane="2" entrytime="00:21:54.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.00" />
                    <SPLIT distance="100" swimtime="00:01:20.91" />
                    <SPLIT distance="200" swimtime="00:02:48.18" />
                    <SPLIT distance="250" swimtime="00:03:33.29" />
                    <SPLIT distance="300" swimtime="00:04:18.41" />
                    <SPLIT distance="350" swimtime="00:05:02.62" />
                    <SPLIT distance="400" swimtime="00:05:47.16" />
                    <SPLIT distance="450" swimtime="00:06:32.52" />
                    <SPLIT distance="500" swimtime="00:07:18.20" />
                    <SPLIT distance="550" swimtime="00:08:02.76" />
                    <SPLIT distance="600" swimtime="00:08:48.23" />
                    <SPLIT distance="650" swimtime="00:09:34.00" />
                    <SPLIT distance="700" swimtime="00:10:20.00" />
                    <SPLIT distance="750" swimtime="00:11:06.05" />
                    <SPLIT distance="800" swimtime="00:11:52.26" />
                    <SPLIT distance="850" swimtime="00:12:38.04" />
                    <SPLIT distance="900" swimtime="00:13:24.21" />
                    <SPLIT distance="950" swimtime="00:14:09.47" />
                    <SPLIT distance="1000" swimtime="00:14:55.48" />
                    <SPLIT distance="1050" swimtime="00:15:40.72" />
                    <SPLIT distance="1100" swimtime="00:16:27.13" />
                    <SPLIT distance="1150" swimtime="00:17:13.79" />
                    <SPLIT distance="1200" swimtime="00:18:00.17" />
                    <SPLIT distance="1250" swimtime="00:18:46.25" />
                    <SPLIT distance="1300" swimtime="00:19:32.06" />
                    <SPLIT distance="1350" swimtime="00:20:17.65" />
                    <SPLIT distance="1400" swimtime="00:21:02.93" />
                    <SPLIT distance="1450" swimtime="00:21:47.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1420" points="433" swimtime="00:02:35.85" resultid="1969" heatid="2220" lane="2" entrytime="00:02:39.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                    <SPLIT distance="100" swimtime="00:01:15.50" />
                    <SPLIT distance="150" swimtime="00:01:55.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Teodoro" lastname="Valenca Wacholski" birthdate="2002-10-23" gender="M" nation="BRA" license="V413180" athleteid="1953" externalid="V413180">
              <RESULTS>
                <RESULT eventid="1204" points="417" swimtime="00:20:43.57" resultid="1954" heatid="2181" lane="1" entrytime="00:21:03.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:11.91" />
                    <SPLIT distance="150" swimtime="00:01:51.54" />
                    <SPLIT distance="200" swimtime="00:02:31.75" />
                    <SPLIT distance="250" swimtime="00:03:12.06" />
                    <SPLIT distance="300" swimtime="00:03:53.16" />
                    <SPLIT distance="350" swimtime="00:04:34.42" />
                    <SPLIT distance="400" swimtime="00:05:17.78" />
                    <SPLIT distance="450" swimtime="00:06:01.27" />
                    <SPLIT distance="500" swimtime="00:06:44.44" />
                    <SPLIT distance="550" swimtime="00:07:27.45" />
                    <SPLIT distance="600" swimtime="00:08:09.65" />
                    <SPLIT distance="650" swimtime="00:08:52.96" />
                    <SPLIT distance="700" swimtime="00:09:37.99" />
                    <SPLIT distance="750" swimtime="00:10:21.93" />
                    <SPLIT distance="800" swimtime="00:11:04.90" />
                    <SPLIT distance="850" swimtime="00:11:47.11" />
                    <SPLIT distance="900" swimtime="00:12:29.69" />
                    <SPLIT distance="950" swimtime="00:13:12.49" />
                    <SPLIT distance="1000" swimtime="00:13:55.55" />
                    <SPLIT distance="1050" swimtime="00:14:38.40" />
                    <SPLIT distance="1100" swimtime="00:15:20.43" />
                    <SPLIT distance="1150" swimtime="00:16:02.87" />
                    <SPLIT distance="1200" swimtime="00:16:45.23" />
                    <SPLIT distance="1250" swimtime="00:17:27.18" />
                    <SPLIT distance="1300" swimtime="00:18:09.27" />
                    <SPLIT distance="1350" swimtime="00:18:50.44" />
                    <SPLIT distance="1400" swimtime="00:19:30.90" />
                    <SPLIT distance="1450" swimtime="00:20:08.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1234" points="485" swimtime="00:04:56.33" resultid="1955" heatid="2189" lane="5" entrytime="00:05:03.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:12.93" />
                    <SPLIT distance="150" swimtime="00:01:50.74" />
                    <SPLIT distance="200" swimtime="00:02:28.64" />
                    <SPLIT distance="250" swimtime="00:03:06.53" />
                    <SPLIT distance="300" swimtime="00:03:44.59" />
                    <SPLIT distance="350" swimtime="00:04:21.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1286" points="501" swimtime="00:00:26.78" resultid="1956" heatid="2199" lane="4" />
                <RESULT eventid="1433" points="473" swimtime="00:02:14.63" resultid="1957" heatid="2223" lane="1" entrytime="00:02:25.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                    <SPLIT distance="100" swimtime="00:01:06.44" />
                    <SPLIT distance="150" swimtime="00:01:41.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1381" points="442" swimtime="00:10:40.21" resultid="1958" heatid="2214" lane="5" entrytime="00:10:50.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                    <SPLIT distance="100" swimtime="00:01:10.83" />
                    <SPLIT distance="150" swimtime="00:01:49.01" />
                    <SPLIT distance="200" swimtime="00:02:29.12" />
                    <SPLIT distance="250" swimtime="00:03:09.42" />
                    <SPLIT distance="300" swimtime="00:03:50.06" />
                    <SPLIT distance="350" swimtime="00:04:30.79" />
                    <SPLIT distance="400" swimtime="00:05:12.70" />
                    <SPLIT distance="450" swimtime="00:05:54.93" />
                    <SPLIT distance="500" swimtime="00:06:37.07" />
                    <SPLIT distance="550" swimtime="00:07:20.02" />
                    <SPLIT distance="600" swimtime="00:08:02.17" />
                    <SPLIT distance="650" swimtime="00:08:44.12" />
                    <SPLIT distance="700" swimtime="00:09:26.14" />
                    <SPLIT distance="750" swimtime="00:10:05.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="UTFPR (CURITIBA) &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1219" swimtime="00:04:19.83" resultid="1988" heatid="2184" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                    <SPLIT distance="100" swimtime="00:01:01.22" />
                    <SPLIT distance="150" swimtime="00:01:31.07" />
                    <SPLIT distance="200" swimtime="00:02:04.50" />
                    <SPLIT distance="250" swimtime="00:02:33.18" />
                    <SPLIT distance="300" swimtime="00:03:02.83" />
                    <SPLIT distance="350" swimtime="00:03:36.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1953" number="1" />
                    <RELAYPOSITION athleteid="1948" number="2" />
                    <RELAYPOSITION athleteid="1944" number="3" />
                    <RELAYPOSITION athleteid="1981" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1379" swimtime="00:10:29.67" resultid="1989" heatid="2212" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.92" />
                    <SPLIT distance="100" swimtime="00:01:10.14" />
                    <SPLIT distance="150" swimtime="00:01:47.07" />
                    <SPLIT distance="200" swimtime="00:02:21.55" />
                    <SPLIT distance="250" swimtime="00:02:56.58" />
                    <SPLIT distance="300" swimtime="00:03:34.02" />
                    <SPLIT distance="350" swimtime="00:04:11.18" />
                    <SPLIT distance="400" swimtime="00:04:45.58" />
                    <SPLIT distance="450" swimtime="00:05:25.82" />
                    <SPLIT distance="500" swimtime="00:06:10.94" />
                    <SPLIT distance="550" swimtime="00:06:59.58" />
                    <SPLIT distance="600" swimtime="00:07:48.83" />
                    <SPLIT distance="650" swimtime="00:08:24.46" />
                    <SPLIT distance="700" swimtime="00:09:05.48" />
                    <SPLIT distance="750" swimtime="00:09:47.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1953" number="1" />
                    <RELAYPOSITION athleteid="1944" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1981" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1948" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1511" swimtime="00:05:03.47" resultid="1990" heatid="2236" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="100" swimtime="00:01:16.57" />
                    <SPLIT distance="150" swimtime="00:01:54.13" />
                    <SPLIT distance="200" swimtime="00:02:37.40" />
                    <SPLIT distance="250" swimtime="00:03:09.64" />
                    <SPLIT distance="300" swimtime="00:03:47.30" />
                    <SPLIT distance="350" swimtime="00:04:19.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1948" number="1" />
                    <RELAYPOSITION athleteid="1953" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1944" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1981" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="UTFPR (CURITIBA) &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1217" swimtime="00:05:02.64" resultid="1985" heatid="2182" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:17.99" />
                    <SPLIT distance="150" swimtime="00:01:54.84" />
                    <SPLIT distance="200" swimtime="00:02:36.28" />
                    <SPLIT distance="250" swimtime="00:03:12.99" />
                    <SPLIT distance="300" swimtime="00:03:50.88" />
                    <SPLIT distance="350" swimtime="00:04:24.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1959" number="1" />
                    <RELAYPOSITION athleteid="1970" number="2" />
                    <RELAYPOSITION athleteid="1976" number="3" />
                    <RELAYPOSITION athleteid="1964" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1377" swimtime="00:11:12.53" resultid="1986" heatid="2211" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.21" />
                    <SPLIT distance="100" swimtime="00:01:19.45" />
                    <SPLIT distance="150" swimtime="00:02:03.13" />
                    <SPLIT distance="200" swimtime="00:02:47.59" />
                    <SPLIT distance="250" swimtime="00:03:24.15" />
                    <SPLIT distance="300" swimtime="00:04:07.39" />
                    <SPLIT distance="350" swimtime="00:04:57.99" />
                    <SPLIT distance="400" swimtime="00:05:45.05" />
                    <SPLIT distance="450" swimtime="00:06:23.62" />
                    <SPLIT distance="500" swimtime="00:07:06.86" />
                    <SPLIT distance="550" swimtime="00:07:51.41" />
                    <SPLIT distance="600" swimtime="00:08:34.22" />
                    <SPLIT distance="650" swimtime="00:09:09.50" />
                    <SPLIT distance="700" swimtime="00:09:48.56" />
                    <SPLIT distance="750" swimtime="00:10:29.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1959" number="1" />
                    <RELAYPOSITION athleteid="1970" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1976" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1964" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1513" swimtime="00:05:57.19" resultid="1987" heatid="2237" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                    <SPLIT distance="100" swimtime="00:01:31.88" />
                    <SPLIT distance="150" swimtime="00:02:17.51" />
                    <SPLIT distance="200" swimtime="00:03:10.13" />
                    <SPLIT distance="250" swimtime="00:03:50.93" />
                    <SPLIT distance="300" swimtime="00:04:39.52" />
                    <SPLIT distance="350" swimtime="00:05:14.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1976" number="1" />
                    <RELAYPOSITION athleteid="1970" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1964" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1959" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="UNATTACHED">
          <OFFICIALS>
            <OFFICIAL officialid="2246" gender="M" />
          </OFFICIALS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
