<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.79413">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Curitiba" name="Troféu Luciano Cabrine (Infantil/Sênior) 2024" course="LCM" deadline="2024-04-07" entrystartdate="2024-03-31" entrytype="INVITATION" hostclub="Clube Curitibano" hostclub.url="https://clubecuritibano.com.br/" number="38307" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/evento/natacao/" startmethod="1" timing="AUTOMATIC" masters="F" withdrawuntil="2024-04-09" state="PR" nation="BRA">
      <AGEDATE value="2024-04-12" type="YEAR" />
      <POOL name="Parque Aquático do Clube Curitibano" lanemax="9" />
      <FACILITY city="Curitiba" name="Parque Aquático do Clube Curitibano" nation="BRA" state="PR" street="Avenida Presidente Getúlio Vargas, 2857" street2="Água Verde" zip="80240-040" />
      <POINTTABLE pointtableid="3017" name="FINA Point Scoring" version="2024" />
      <QUALIFY from="2023-04-12" until="2024-04-11" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-04-12" daytime="08:45" endtime="13:41" number="1" officialmeeting="08:00" teamleadermeeting="08:30" warmupfrom="07:30" warmupuntil="08:30">
          <EVENTS>
            <EVENT eventid="1064" daytime="08:46" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1065" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2824" />
                    <RANKING order="2" place="2" resultid="2806" />
                    <RANKING order="3" place="3" resultid="2870" />
                    <RANKING order="4" place="4" resultid="1538" />
                    <RANKING order="5" place="5" resultid="2946" />
                    <RANKING order="6" place="6" resultid="2326" />
                    <RANKING order="7" place="7" resultid="2002" />
                    <RANKING order="8" place="-1" resultid="2398" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2272" />
                    <RANKING order="2" place="2" resultid="1428" />
                    <RANKING order="3" place="3" resultid="2671" />
                    <RANKING order="4" place="4" resultid="3807" />
                    <RANKING order="5" place="5" resultid="1678" />
                    <RANKING order="6" place="6" resultid="1434" />
                    <RANKING order="7" place="7" resultid="2689" />
                    <RANKING order="8" place="8" resultid="1767" />
                    <RANKING order="9" place="9" resultid="2993" />
                    <RANKING order="10" place="10" resultid="2713" />
                    <RANKING order="11" place="11" resultid="3324" />
                    <RANKING order="12" place="12" resultid="3723" />
                    <RANKING order="13" place="13" resultid="3717" />
                    <RANKING order="14" place="14" resultid="2416" />
                    <RANKING order="15" place="15" resultid="3384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1870" />
                    <RANKING order="2" place="2" resultid="1476" />
                    <RANKING order="3" place="3" resultid="2626" />
                    <RANKING order="4" place="4" resultid="1610" />
                    <RANKING order="5" place="5" resultid="2278" />
                    <RANKING order="6" place="6" resultid="1492" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2964" />
                    <RANKING order="2" place="2" resultid="2266" />
                    <RANKING order="3" place="3" resultid="2044" />
                    <RANKING order="4" place="4" resultid="3262" />
                    <RANKING order="5" place="5" resultid="1416" />
                    <RANKING order="6" place="6" resultid="3396" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3488" />
                    <RANKING order="2" place="2" resultid="1486" />
                    <RANKING order="3" place="3" resultid="1972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2069" />
                    <RANKING order="2" place="2" resultid="1735" />
                    <RANKING order="3" place="3" resultid="3795" />
                    <RANKING order="4" place="4" resultid="3307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4266" daytime="08:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4267" daytime="08:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4268" daytime="08:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4269" daytime="09:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4270" daytime="09:06" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4271" daytime="09:10" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1072" daytime="09:14" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1073" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2858" />
                    <RANKING order="2" place="2" resultid="2302" />
                    <RANKING order="3" place="3" resultid="2308" />
                    <RANKING order="4" place="4" resultid="3577" />
                    <RANKING order="5" place="5" resultid="2770" />
                    <RANKING order="6" place="6" resultid="2392" />
                    <RANKING order="7" place="7" resultid="3172" />
                    <RANKING order="8" place="8" resultid="3124" />
                    <RANKING order="9" place="9" resultid="3226" />
                    <RANKING order="10" place="-1" resultid="3190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2284" />
                    <RANKING order="2" place="2" resultid="2929" />
                    <RANKING order="3" place="3" resultid="2141" />
                    <RANKING order="4" place="4" resultid="2701" />
                    <RANKING order="5" place="5" resultid="2153" />
                    <RANKING order="6" place="6" resultid="2665" />
                    <RANKING order="7" place="7" resultid="2380" />
                    <RANKING order="8" place="8" resultid="1642" />
                    <RANKING order="9" place="9" resultid="1955" />
                    <RANKING order="10" place="10" resultid="3677" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1875" />
                    <RANKING order="2" place="2" resultid="3007" />
                    <RANKING order="3" place="3" resultid="2636" />
                    <RANKING order="4" place="4" resultid="3178" />
                    <RANKING order="5" place="5" resultid="2117" />
                    <RANKING order="6" place="6" resultid="2601" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1076" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2642" />
                    <RANKING order="2" place="2" resultid="2474" />
                    <RANKING order="3" place="3" resultid="2576" />
                    <RANKING order="4" place="4" resultid="2571" />
                    <RANKING order="5" place="5" resultid="3784" />
                    <RANKING order="6" place="6" resultid="2597" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1077" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2988" />
                    <RANKING order="2" place="2" resultid="3405" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2466" />
                    <RANKING order="2" place="2" resultid="2469" />
                    <RANKING order="3" place="3" resultid="3559" />
                    <RANKING order="4" place="4" resultid="2081" />
                    <RANKING order="5" place="5" resultid="2093" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2835" />
                    <RANKING order="2" place="2" resultid="2075" />
                    <RANKING order="3" place="3" resultid="2422" />
                    <RANKING order="4" place="4" resultid="1885" />
                    <RANKING order="5" place="5" resultid="2087" />
                    <RANKING order="6" place="6" resultid="3130" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4272" daytime="09:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4273" daytime="09:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4274" daytime="09:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4275" daytime="09:28" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4276" daytime="09:32" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4277" daytime="09:38" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1080" daytime="09:42" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1081" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2882" />
                    <RANKING order="2" place="2" resultid="2776" />
                    <RANKING order="3" place="3" resultid="2800" />
                    <RANKING order="4" place="4" resultid="2368" />
                    <RANKING order="5" place="5" resultid="2952" />
                    <RANKING order="6" place="6" resultid="3822" />
                    <RANKING order="7" place="7" resultid="3641" />
                    <RANKING order="8" place="8" resultid="3166" />
                    <RANKING order="9" place="9" resultid="3571" />
                    <RANKING order="10" place="10" resultid="2788" />
                    <RANKING order="11" place="11" resultid="1708" />
                    <RANKING order="12" place="12" resultid="3689" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3653" />
                    <RANKING order="2" place="2" resultid="2374" />
                    <RANKING order="3" place="3" resultid="2527" />
                    <RANKING order="4" place="4" resultid="3289" />
                    <RANKING order="5" place="5" resultid="2917" />
                    <RANKING order="6" place="6" resultid="3659" />
                    <RANKING order="7" place="7" resultid="3136" />
                    <RANKING order="8" place="8" resultid="2864" />
                    <RANKING order="9" place="9" resultid="2147" />
                    <RANKING order="10" place="10" resultid="1532" />
                    <RANKING order="11" place="-1" resultid="3813" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2611" />
                    <RANKING order="2" place="2" resultid="1943" />
                    <RANKING order="3" place="3" resultid="2616" />
                    <RANKING order="4" place="4" resultid="3100" />
                    <RANKING order="5" place="-1" resultid="2532" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2446" />
                    <RANKING order="2" place="2" resultid="2876" />
                    <RANKING order="3" place="3" resultid="2314" />
                    <RANKING order="4" place="4" resultid="1752" />
                    <RANKING order="5" place="5" resultid="3512" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2499" />
                    <RANKING order="2" place="2" resultid="1966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2979" />
                    <RANKING order="2" place="2" resultid="3087" />
                    <RANKING order="3" place="-1" resultid="1470" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3060" />
                    <RANKING order="2" place="2" resultid="2254" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4278" daytime="09:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4279" daytime="09:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4280" daytime="09:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4281" daytime="09:56" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4282" daytime="10:00" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1088" daytime="10:04" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1089" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2320" />
                    <RANKING order="2" place="2" resultid="1654" />
                    <RANKING order="3" place="3" resultid="2764" />
                    <RANKING order="4" place="4" resultid="2812" />
                    <RANKING order="5" place="5" resultid="2338" />
                    <RANKING order="6" place="6" resultid="2897" />
                    <RANKING order="7" place="7" resultid="1593" />
                    <RANKING order="8" place="8" resultid="3593" />
                    <RANKING order="9" place="9" resultid="2362" />
                    <RANKING order="10" place="10" resultid="2404" />
                    <RANKING order="11" place="11" resultid="1842" />
                    <RANKING order="12" place="12" resultid="3647" />
                    <RANKING order="13" place="13" resultid="2782" />
                    <RANKING order="14" place="-1" resultid="2830" />
                    <RANKING order="15" place="-1" resultid="1859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3160" />
                    <RANKING order="2" place="2" resultid="2719" />
                    <RANKING order="3" place="3" resultid="2659" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1460" />
                    <RANKING order="2" place="2" resultid="3671" />
                    <RANKING order="3" place="3" resultid="3295" />
                    <RANKING order="4" place="4" resultid="2621" />
                    <RANKING order="5" place="5" resultid="1914" />
                    <RANKING order="6" place="6" resultid="1581" />
                    <RANKING order="7" place="7" resultid="2344" />
                    <RANKING order="8" place="8" resultid="1672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1092" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2479" />
                    <RANKING order="2" place="2" resultid="2495" />
                    <RANKING order="3" place="3" resultid="1620" />
                    <RANKING order="4" place="4" resultid="2892" />
                    <RANKING order="5" place="5" resultid="2099" />
                    <RANKING order="6" place="6" resultid="2356" />
                    <RANKING order="7" place="7" resultid="1587" />
                    <RANKING order="8" place="8" resultid="2903" />
                    <RANKING order="9" place="9" resultid="3142" />
                    <RANKING order="10" place="10" resultid="2129" />
                    <RANKING order="11" place="11" resultid="2213" />
                    <RANKING order="12" place="-1" resultid="3318" />
                    <RANKING order="13" place="-1" resultid="2587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2554" />
                    <RANKING order="2" place="2" resultid="1405" />
                    <RANKING order="3" place="3" resultid="2296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2514" />
                    <RANKING order="2" place="2" resultid="1599" />
                    <RANKING order="3" place="3" resultid="2230" />
                    <RANKING order="4" place="4" resultid="3801" />
                    <RANKING order="5" place="5" resultid="3253" />
                    <RANKING order="6" place="-1" resultid="3617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2560" />
                    <RANKING order="2" place="2" resultid="2999" />
                    <RANKING order="3" place="3" resultid="1559" />
                    <RANKING order="4" place="4" resultid="1466" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4283" daytime="10:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4284" daytime="10:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4285" daytime="10:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4286" daytime="10:18" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4287" daytime="10:22" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4288" daytime="10:26" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4289" daytime="10:30" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1096" daytime="10:34" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1097" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1696" />
                    <RANKING order="2" place="2" resultid="1660" />
                    <RANKING order="3" place="3" resultid="2410" />
                    <RANKING order="4" place="4" resultid="3817" />
                    <RANKING order="5" place="5" resultid="1666" />
                    <RANKING order="6" place="6" resultid="3572" />
                    <RANKING order="7" place="7" resultid="1709" />
                    <RANKING order="8" place="8" resultid="1783" />
                    <RANKING order="9" place="9" resultid="3642" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3611" />
                    <RANKING order="2" place="2" resultid="1684" />
                    <RANKING order="3" place="3" resultid="3705" />
                    <RANKING order="4" place="4" resultid="3808" />
                    <RANKING order="5" place="5" resultid="3390" />
                    <RANKING order="6" place="6" resultid="1814" />
                    <RANKING order="7" place="7" resultid="3385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3482" />
                    <RANKING order="2" place="2" resultid="2461" />
                    <RANKING order="3" place="3" resultid="3635" />
                    <RANKING order="4" place="4" resultid="1615" />
                    <RANKING order="5" place="5" resultid="1949" />
                    <RANKING order="6" place="6" resultid="3565" />
                    <RANKING order="7" place="7" resultid="3417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2455" />
                    <RANKING order="2" place="2" resultid="1746" />
                    <RANKING order="3" place="3" resultid="1631" />
                    <RANKING order="4" place="4" resultid="1992" />
                    <RANKING order="5" place="5" resultid="1778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2057" />
                    <RANKING order="2" place="2" resultid="1973" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3500" />
                    <RANKING order="2" place="2" resultid="3313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2236" />
                    <RANKING order="2" place="2" resultid="3789" />
                    <RANKING order="3" place="3" resultid="3061" />
                    <RANKING order="4" place="4" resultid="3379" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4290" daytime="10:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4291" daytime="10:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4292" daytime="10:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4293" daytime="10:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4294" daytime="10:42" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1104" daytime="10:44" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1105" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1648" />
                    <RANKING order="2" place="2" resultid="2303" />
                    <RANKING order="3" place="3" resultid="3629" />
                    <RANKING order="4" place="4" resultid="3683" />
                    <RANKING order="5" place="5" resultid="3184" />
                    <RANKING order="6" place="6" resultid="1853" />
                    <RANKING order="7" place="7" resultid="1594" />
                    <RANKING order="8" place="8" resultid="1920" />
                    <RANKING order="9" place="9" resultid="2223" />
                    <RANKING order="10" place="10" resultid="1521" />
                    <RANKING order="11" place="11" resultid="3402" />
                    <RANKING order="12" place="-1" resultid="1690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1569" />
                    <RANKING order="2" place="2" resultid="3583" />
                    <RANKING order="3" place="3" resultid="3605" />
                    <RANKING order="4" place="4" resultid="3666" />
                    <RANKING order="5" place="5" resultid="1956" />
                    <RANKING order="6" place="6" resultid="3440" />
                    <RANKING order="7" place="7" resultid="1714" />
                    <RANKING order="8" place="8" resultid="2014" />
                    <RANKING order="9" place="9" resultid="2020" />
                    <RANKING order="10" place="10" resultid="2026" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1107" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1563" />
                    <RANKING order="2" place="2" resultid="3518" />
                    <RANKING order="3" place="3" resultid="2970" />
                    <RANKING order="4" place="4" resultid="1626" />
                    <RANKING order="5" place="5" resultid="1498" />
                    <RANKING order="6" place="6" resultid="2606" />
                    <RANKING order="7" place="7" resultid="3424" />
                    <RANKING order="8" place="8" resultid="3711" />
                    <RANKING order="9" place="9" resultid="1978" />
                    <RANKING order="10" place="10" resultid="3065" />
                    <RANKING order="11" place="11" resultid="2632" />
                    <RANKING order="12" place="12" resultid="1931" />
                    <RANKING order="13" place="13" resultid="3449" />
                    <RANKING order="14" place="-1" resultid="2648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1108" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2582" />
                    <RANKING order="2" place="2" resultid="2490" />
                    <RANKING order="3" place="3" resultid="3148" />
                    <RANKING order="4" place="4" resultid="2941" />
                    <RANKING order="5" place="5" resultid="3785" />
                    <RANKING order="6" place="6" resultid="2386" />
                    <RANKING order="7" place="7" resultid="3506" />
                    <RANKING order="8" place="8" resultid="3536" />
                    <RANKING order="9" place="9" resultid="1575" />
                    <RANKING order="10" place="10" resultid="2912" />
                    <RANKING order="11" place="11" resultid="1702" />
                    <RANKING order="12" place="12" resultid="3094" />
                    <RANKING order="13" place="13" resultid="1762" />
                    <RANKING order="14" place="14" resultid="1987" />
                    <RANKING order="15" place="15" resultid="1996" />
                    <RANKING order="16" place="16" resultid="3458" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2548" />
                    <RANKING order="2" place="2" resultid="3268" />
                    <RANKING order="3" place="3" resultid="2508" />
                    <RANKING order="4" place="4" resultid="3738" />
                    <RANKING order="5" place="5" resultid="3429" />
                    <RANKING order="6" place="6" resultid="3453" />
                    <RANKING order="7" place="7" resultid="3360" />
                    <RANKING order="8" place="8" resultid="3202" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1110" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3012" />
                    <RANKING order="2" place="2" resultid="2747" />
                    <RANKING order="3" place="3" resultid="1554" />
                    <RANKING order="4" place="4" resultid="3623" />
                    <RANKING order="5" place="5" resultid="3330" />
                    <RANKING order="6" place="6" resultid="1509" />
                    <RANKING order="7" place="7" resultid="2350" />
                    <RANKING order="8" place="8" resultid="3618" />
                    <RANKING order="9" place="9" resultid="1604" />
                    <RANKING order="10" place="10" resultid="1848" />
                    <RANKING order="11" place="11" resultid="1637" />
                    <RANKING order="12" place="12" resultid="3091" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1820" />
                    <RANKING order="2" place="2" resultid="3744" />
                    <RANKING order="3" place="3" resultid="2923" />
                    <RANKING order="4" place="4" resultid="1411" />
                    <RANKING order="5" place="5" resultid="1826" />
                    <RANKING order="6" place="6" resultid="1890" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4295" daytime="10:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4296" daytime="10:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4297" daytime="10:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4298" daytime="10:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4299" daytime="10:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4300" daytime="10:52" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4301" daytime="10:54" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4302" daytime="10:56" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4303" daytime="10:56" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4304" daytime="10:58" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1112" daytime="11:00" gender="X" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1113" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3043" />
                    <RANKING order="2" place="2" resultid="3056" />
                    <RANKING order="3" place="3" resultid="1729" />
                    <RANKING order="4" place="4" resultid="2425" />
                    <RANKING order="5" place="5" resultid="3776" />
                    <RANKING order="6" place="6" resultid="3249" />
                    <RANKING order="7" place="7" resultid="1732" />
                    <RANKING order="8" place="-1" resultid="2440" />
                    <RANKING order="9" place="-1" resultid="3763" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4305" daytime="11:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4306" daytime="11:08" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1114" daytime="11:14" gender="X" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1115" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3044" />
                    <RANKING order="2" place="2" resultid="1730" />
                    <RANKING order="3" place="3" resultid="3057" />
                    <RANKING order="4" place="4" resultid="2441" />
                    <RANKING order="5" place="5" resultid="3764" />
                    <RANKING order="6" place="6" resultid="3250" />
                    <RANKING order="7" place="-1" resultid="3777" />
                    <RANKING order="8" place="-1" resultid="2183" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4307" daytime="11:14" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1116" daytime="11:22" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1117" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2327" />
                    <RANKING order="2" place="2" resultid="2332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2135" />
                    <RANKING order="2" place="2" resultid="2683" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2521" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1831" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1422" />
                    <RANKING order="2" place="2" resultid="2242" />
                    <RANKING order="3" place="3" resultid="3214" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2888" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2935" />
                    <RANKING order="2" place="2" resultid="2975" />
                    <RANKING order="3" place="3" resultid="3347" />
                    <RANKING order="4" place="-1" resultid="3003" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4308" daytime="11:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4309" daytime="11:46" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1124" daytime="12:10" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1125" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2752" />
                    <RANKING order="2" place="2" resultid="2771" />
                    <RANKING order="3" place="3" resultid="2758" />
                    <RANKING order="4" place="4" resultid="2339" />
                    <RANKING order="5" place="5" resultid="2907" />
                    <RANKING order="6" place="6" resultid="2405" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2695" />
                    <RANKING order="2" place="2" resultid="2846" />
                    <RANKING order="3" place="3" resultid="2707" />
                    <RANKING order="4" place="4" resultid="2741" />
                    <RANKING order="5" place="5" resultid="3665" />
                    <RANKING order="6" place="6" resultid="2290" />
                    <RANKING order="7" place="-1" resultid="2381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2260" />
                    <RANKING order="2" place="2" resultid="3274" />
                    <RANKING order="3" place="3" resultid="2637" />
                    <RANKING order="4" place="4" resultid="2537" />
                    <RANKING order="5" place="5" resultid="1503" />
                    <RANKING order="6" place="6" resultid="2602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2248" />
                    <RANKING order="2" place="2" resultid="2852" />
                    <RANKING order="3" place="3" resultid="2357" />
                    <RANKING order="4" place="4" resultid="2591" />
                    <RANKING order="5" place="5" resultid="2123" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3494" />
                    <RANKING order="2" place="2" resultid="2105" />
                    <RANKING order="3" place="3" resultid="3729" />
                    <RANKING order="4" place="4" resultid="3359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3258" />
                    <RANKING order="2" place="2" resultid="2565" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3335" />
                    <RANKING order="2" place="2" resultid="1900" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4310" daytime="12:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4311" daytime="12:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4312" daytime="12:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4313" daytime="12:46" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-04-12" daytime="16:15" endtime="20:10" number="2" officialmeeting="16:30" warmupfrom="15:00" warmupuntil="16:00">
          <EVENTS>
            <EVENT eventid="1132" daytime="16:16" gender="F" number="11" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1133" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2328" />
                    <RANKING order="2" place="2" resultid="2412" />
                    <RANKING order="3" place="3" resultid="2369" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1134" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2273" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2450" />
                    <RANKING order="2" place="2" resultid="2279" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2045" />
                    <RANKING order="2" place="2" resultid="2316" />
                    <RANKING order="3" place="3" resultid="3263" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1137" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2244" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1139" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2936" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4314" daytime="16:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4315" daytime="16:22" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1140" daytime="16:32" gender="M" number="12" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1141" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2321" />
                    <RANKING order="2" place="2" resultid="2309" />
                    <RANKING order="3" place="3" resultid="2393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2285" />
                    <RANKING order="2" place="2" resultid="1925" />
                    <RANKING order="3" place="-1" resultid="3606" />
                    <RANKING order="4" place="-1" resultid="2731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1143" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1876" />
                    <RANKING order="2" place="2" resultid="1462" />
                    <RANKING order="3" place="3" resultid="3275" />
                    <RANKING order="4" place="4" resultid="2538" />
                    <RANKING order="5" place="5" resultid="2345" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1144" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2250" />
                    <RANKING order="2" place="2" resultid="2480" />
                    <RANKING order="3" place="3" resultid="2100" />
                    <RANKING order="4" place="-1" resultid="2475" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2470" />
                    <RANKING order="2" place="2" resultid="1605" />
                    <RANKING order="3" place="-1" resultid="2351" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2088" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4316" daytime="16:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4317" daytime="16:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4318" daytime="16:46" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1148" daytime="16:52" gender="F" number="13" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1149" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2825" />
                    <RANKING order="2" place="2" resultid="2807" />
                    <RANKING order="3" place="3" resultid="2801" />
                    <RANKING order="4" place="4" resultid="1539" />
                    <RANKING order="5" place="5" resultid="3823" />
                    <RANKING order="6" place="6" resultid="2777" />
                    <RANKING order="7" place="7" resultid="1697" />
                    <RANKING order="8" place="8" resultid="2871" />
                    <RANKING order="9" place="9" resultid="2199" />
                    <RANKING order="10" place="10" resultid="3167" />
                    <RANKING order="11" place="11" resultid="2947" />
                    <RANKING order="12" place="12" resultid="3208" />
                    <RANKING order="13" place="13" resultid="2789" />
                    <RANKING order="14" place="14" resultid="1661" />
                    <RANKING order="15" place="15" resultid="3301" />
                    <RANKING order="16" place="16" resultid="1667" />
                    <RANKING order="17" place="17" resultid="2003" />
                    <RANKING order="18" place="18" resultid="1808" />
                    <RANKING order="19" place="19" resultid="1789" />
                    <RANKING order="20" place="20" resultid="3700" />
                    <RANKING order="21" place="21" resultid="2159" />
                    <RANKING order="22" place="22" resultid="1785" />
                    <RANKING order="23" place="23" resultid="3690" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2677" />
                    <RANKING order="2" place="2" resultid="1435" />
                    <RANKING order="3" place="3" resultid="2684" />
                    <RANKING order="4" place="4" resultid="1429" />
                    <RANKING order="5" place="5" resultid="2528" />
                    <RANKING order="6" place="6" resultid="3706" />
                    <RANKING order="7" place="7" resultid="1768" />
                    <RANKING order="8" place="8" resultid="1685" />
                    <RANKING order="9" place="9" resultid="2690" />
                    <RANKING order="10" place="10" resultid="2918" />
                    <RANKING order="11" place="11" resultid="2714" />
                    <RANKING order="12" place="12" resultid="3654" />
                    <RANKING order="13" place="13" resultid="2148" />
                    <RANKING order="14" place="14" resultid="2672" />
                    <RANKING order="15" place="15" resultid="2136" />
                    <RANKING order="16" place="16" resultid="3660" />
                    <RANKING order="17" place="17" resultid="2417" />
                    <RANKING order="18" place="18" resultid="2840" />
                    <RANKING order="19" place="19" resultid="1815" />
                    <RANKING order="20" place="20" resultid="1741" />
                    <RANKING order="21" place="21" resultid="2865" />
                    <RANKING order="22" place="22" resultid="3718" />
                    <RANKING order="23" place="23" resultid="3724" />
                    <RANKING order="24" place="24" resultid="3391" />
                    <RANKING order="25" place="25" resultid="1533" />
                    <RANKING order="26" place="26" resultid="3238" />
                    <RANKING order="27" place="27" resultid="3386" />
                    <RANKING order="28" place="28" resultid="1799" />
                    <RANKING order="29" place="29" resultid="3115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1151" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2462" />
                    <RANKING order="2" place="2" resultid="2522" />
                    <RANKING order="3" place="3" resultid="3636" />
                    <RANKING order="4" place="4" resultid="1477" />
                    <RANKING order="5" place="5" resultid="3154" />
                    <RANKING order="6" place="6" resultid="3530" />
                    <RANKING order="7" place="7" resultid="2627" />
                    <RANKING order="8" place="8" resultid="1871" />
                    <RANKING order="9" place="9" resultid="1950" />
                    <RANKING order="10" place="10" resultid="3542" />
                    <RANKING order="11" place="11" resultid="3566" />
                    <RANKING order="12" place="12" resultid="2111" />
                    <RANKING order="13" place="13" resultid="3418" />
                    <RANKING order="14" place="14" resultid="1616" />
                    <RANKING order="15" place="15" resultid="3101" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1152" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3411" />
                    <RANKING order="2" place="2" resultid="1747" />
                    <RANKING order="3" place="3" resultid="2267" />
                    <RANKING order="4" place="4" resultid="2877" />
                    <RANKING order="5" place="5" resultid="2965" />
                    <RANKING order="6" place="6" resultid="3353" />
                    <RANKING order="7" place="7" resultid="3513" />
                    <RANKING order="8" place="8" resultid="1417" />
                    <RANKING order="9" place="9" resultid="1832" />
                    <RANKING order="10" place="10" resultid="1632" />
                    <RANKING order="11" place="11" resultid="1779" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2543" />
                    <RANKING order="2" place="2" resultid="1423" />
                    <RANKING order="3" place="3" resultid="2058" />
                    <RANKING order="4" place="4" resultid="1487" />
                    <RANKING order="5" place="5" resultid="1974" />
                    <RANKING order="6" place="6" resultid="1967" />
                    <RANKING order="7" place="-1" resultid="1482" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1736" />
                    <RANKING order="2" place="2" resultid="2070" />
                    <RANKING order="3" place="3" resultid="3501" />
                    <RANKING order="4" place="4" resultid="3796" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3554" />
                    <RANKING order="2" place="2" resultid="2237" />
                    <RANKING order="3" place="3" resultid="3380" />
                    <RANKING order="4" place="4" resultid="3348" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4319" daytime="16:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4320" daytime="16:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4321" daytime="16:58" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4322" daytime="17:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4323" daytime="17:02" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4324" daytime="17:04" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4325" daytime="17:08" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4326" daytime="17:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4327" daytime="17:12" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4328" daytime="17:14" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4329" daytime="17:16" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4330" daytime="17:18" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1156" daytime="17:20" gender="M" number="14" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1157" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2859" />
                    <RANKING order="2" place="2" resultid="1649" />
                    <RANKING order="3" place="3" resultid="2813" />
                    <RANKING order="4" place="4" resultid="1794" />
                    <RANKING order="5" place="5" resultid="2765" />
                    <RANKING order="6" place="6" resultid="2171" />
                    <RANKING order="7" place="7" resultid="2753" />
                    <RANKING order="8" place="8" resultid="3630" />
                    <RANKING order="9" place="9" resultid="3599" />
                    <RANKING order="10" place="10" resultid="1526" />
                    <RANKING order="11" place="11" resultid="2204" />
                    <RANKING order="12" place="12" resultid="3191" />
                    <RANKING order="13" place="13" resultid="3173" />
                    <RANKING order="14" place="14" resultid="3684" />
                    <RANKING order="15" place="15" resultid="2818" />
                    <RANKING order="16" place="16" resultid="1854" />
                    <RANKING order="17" place="17" resultid="3365" />
                    <RANKING order="18" place="18" resultid="2908" />
                    <RANKING order="19" place="19" resultid="3125" />
                    <RANKING order="20" place="20" resultid="3071" />
                    <RANKING order="21" place="21" resultid="1961" />
                    <RANKING order="22" place="22" resultid="3435" />
                    <RANKING order="23" place="23" resultid="1522" />
                    <RANKING order="24" place="24" resultid="3589" />
                    <RANKING order="25" place="25" resultid="1691" />
                    <RANKING order="26" place="26" resultid="1921" />
                    <RANKING order="27" place="27" resultid="1860" />
                    <RANKING order="28" place="28" resultid="1803" />
                    <RANKING order="29" place="29" resultid="2224" />
                    <RANKING order="30" place="30" resultid="3227" />
                    <RANKING order="31" place="31" resultid="3232" />
                    <RANKING order="32" place="32" resultid="1843" />
                    <RANKING order="33" place="33" resultid="2165" />
                    <RANKING order="34" place="34" resultid="3695" />
                    <RANKING order="35" place="35" resultid="3403" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1570" />
                    <RANKING order="2" place="2" resultid="2847" />
                    <RANKING order="3" place="3" resultid="2930" />
                    <RANKING order="4" place="4" resultid="2696" />
                    <RANKING order="5" place="5" resultid="2660" />
                    <RANKING order="6" place="6" resultid="2702" />
                    <RANKING order="7" place="7" resultid="2720" />
                    <RANKING order="8" place="8" resultid="2742" />
                    <RANKING order="9" place="9" resultid="2708" />
                    <RANKING order="10" place="10" resultid="2142" />
                    <RANKING order="11" place="11" resultid="2154" />
                    <RANKING order="12" place="12" resultid="2730" />
                    <RANKING order="13" place="13" resultid="2666" />
                    <RANKING order="14" place="14" resultid="1715" />
                    <RANKING order="15" place="15" resultid="1957" />
                    <RANKING order="16" place="16" resultid="2015" />
                    <RANKING order="17" place="17" resultid="2027" />
                    <RANKING order="18" place="18" resultid="3678" />
                    <RANKING order="19" place="19" resultid="3220" />
                    <RANKING order="20" place="20" resultid="2021" />
                    <RANKING order="21" place="21" resultid="2210" />
                    <RANKING order="22" place="22" resultid="3111" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1454" />
                    <RANKING order="2" place="2" resultid="1564" />
                    <RANKING order="3" place="3" resultid="2485" />
                    <RANKING order="4" place="4" resultid="3008" />
                    <RANKING order="5" place="5" resultid="1937" />
                    <RANKING order="6" place="6" resultid="3524" />
                    <RANKING order="7" place="7" resultid="2607" />
                    <RANKING order="8" place="8" resultid="3519" />
                    <RANKING order="9" place="9" resultid="1499" />
                    <RANKING order="10" place="10" resultid="3548" />
                    <RANKING order="11" place="11" resultid="1915" />
                    <RANKING order="12" place="12" resultid="1504" />
                    <RANKING order="13" place="13" resultid="2638" />
                    <RANKING order="14" place="14" resultid="3672" />
                    <RANKING order="15" place="15" resultid="3179" />
                    <RANKING order="16" place="16" resultid="1979" />
                    <RANKING order="17" place="17" resultid="3066" />
                    <RANKING order="18" place="18" resultid="3712" />
                    <RANKING order="19" place="19" resultid="2118" />
                    <RANKING order="20" place="20" resultid="3341" />
                    <RANKING order="21" place="21" resultid="2633" />
                    <RANKING order="22" place="22" resultid="3075" />
                    <RANKING order="23" place="23" resultid="1932" />
                    <RANKING order="24" place="24" resultid="2008" />
                    <RANKING order="25" place="25" resultid="2219" />
                    <RANKING order="26" place="26" resultid="3450" />
                    <RANKING order="27" place="-1" resultid="3079" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1160" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2958" />
                    <RANKING order="2" place="2" resultid="2853" />
                    <RANKING order="3" place="3" resultid="2913" />
                    <RANKING order="4" place="4" resultid="3537" />
                    <RANKING order="5" place="5" resultid="2583" />
                    <RANKING order="6" place="6" resultid="1576" />
                    <RANKING order="7" place="7" resultid="2643" />
                    <RANKING order="8" place="8" resultid="2592" />
                    <RANKING order="9" place="9" resultid="1837" />
                    <RANKING order="10" place="10" resultid="2063" />
                    <RANKING order="11" place="11" resultid="3507" />
                    <RANKING order="12" place="12" resultid="2942" />
                    <RANKING order="13" place="13" resultid="2577" />
                    <RANKING order="14" place="14" resultid="3095" />
                    <RANKING order="15" place="15" resultid="1763" />
                    <RANKING order="16" place="16" resultid="2130" />
                    <RANKING order="17" place="17" resultid="1997" />
                    <RANKING order="18" place="18" resultid="2124" />
                    <RANKING order="19" place="19" resultid="1703" />
                    <RANKING order="20" place="20" resultid="3143" />
                    <RANKING order="21" place="21" resultid="2214" />
                    <RANKING order="22" place="22" resultid="1773" />
                    <RANKING order="23" place="-1" resultid="1988" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1161" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2549" />
                    <RANKING order="2" place="2" resultid="3495" />
                    <RANKING order="3" place="3" resultid="2989" />
                    <RANKING order="4" place="4" resultid="3406" />
                    <RANKING order="5" place="5" resultid="3269" />
                    <RANKING order="6" place="6" resultid="3739" />
                    <RANKING order="7" place="7" resultid="3196" />
                    <RANKING order="8" place="8" resultid="3730" />
                    <RANKING order="9" place="9" resultid="3454" />
                    <RANKING order="10" place="10" resultid="3430" />
                    <RANKING order="11" place="11" resultid="3203" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1162" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2504" />
                    <RANKING order="2" place="2" resultid="2983" />
                    <RANKING order="3" place="3" resultid="1555" />
                    <RANKING order="4" place="4" resultid="3560" />
                    <RANKING order="5" place="5" resultid="3013" />
                    <RANKING order="6" place="6" resultid="3331" />
                    <RANKING order="7" place="7" resultid="2094" />
                    <RANKING order="8" place="8" resultid="1895" />
                    <RANKING order="9" place="9" resultid="1638" />
                    <RANKING order="10" place="10" resultid="2195" />
                    <RANKING order="11" place="11" resultid="3374" />
                    <RANKING order="12" place="12" resultid="2566" />
                    <RANKING order="13" place="13" resultid="1544" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1163" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2836" />
                    <RANKING order="2" place="2" resultid="2653" />
                    <RANKING order="3" place="3" resultid="1827" />
                    <RANKING order="4" place="4" resultid="2924" />
                    <RANKING order="5" place="5" resultid="1821" />
                    <RANKING order="6" place="6" resultid="1412" />
                    <RANKING order="7" place="7" resultid="1891" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4331" daytime="17:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4332" daytime="17:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4333" daytime="17:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4334" daytime="17:28" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4335" daytime="17:32" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4336" daytime="17:34" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4337" daytime="17:36" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4338" daytime="17:38" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4339" daytime="17:40" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4340" daytime="17:42" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4341" daytime="17:44" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4342" daytime="17:46" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="4343" daytime="17:48" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="4344" daytime="17:50" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="4345" daytime="17:52" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="4346" daytime="17:54" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="4347" daytime="17:56" number="17" order="17" status="OFFICIAL" />
                <HEAT heatid="4348" daytime="17:58" number="18" order="18" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1164" daytime="18:02" gender="F" number="15" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1165" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2883" />
                    <RANKING order="2" place="2" resultid="2333" />
                    <RANKING order="3" place="3" resultid="2411" />
                    <RANKING order="4" place="4" resultid="3818" />
                    <RANKING order="5" place="5" resultid="1784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2724" />
                    <RANKING order="2" place="2" resultid="3612" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2456" />
                    <RANKING order="2" place="2" resultid="2315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1446" />
                    <RANKING order="2" place="2" resultid="2243" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1171" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4349" daytime="18:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4350" daytime="18:06" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1172" daytime="18:10" gender="M" number="16" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1173" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2304" />
                    <RANKING order="2" place="2" resultid="2340" />
                    <RANKING order="3" place="3" resultid="2794" />
                    <RANKING order="4" place="4" resultid="2759" />
                    <RANKING order="5" place="5" resultid="3578" />
                    <RANKING order="6" place="6" resultid="2898" />
                    <RANKING order="7" place="7" resultid="3185" />
                    <RANKING order="8" place="8" resultid="3648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3584" />
                    <RANKING order="2" place="2" resultid="2291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2261" />
                    <RANKING order="2" place="2" resultid="1461" />
                    <RANKING order="3" place="3" resultid="2971" />
                    <RANKING order="4" place="4" resultid="1627" />
                    <RANKING order="5" place="5" resultid="1933" />
                    <RANKING order="6" place="-1" resultid="2649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1176" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2249" />
                    <RANKING order="2" place="2" resultid="2387" />
                    <RANKING order="3" place="3" resultid="2491" />
                    <RANKING order="4" place="4" resultid="3149" />
                    <RANKING order="5" place="5" resultid="3459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1177" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2509" />
                    <RANKING order="2" place="2" resultid="1406" />
                    <RANKING order="3" place="3" resultid="3270" />
                    <RANKING order="4" place="4" resultid="2106" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2748" />
                    <RANKING order="2" place="2" resultid="2082" />
                    <RANKING order="3" place="3" resultid="2231" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1909" />
                    <RANKING order="2" place="2" resultid="3336" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4351" daytime="18:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4352" daytime="18:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4353" daytime="18:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4354" daytime="18:24" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1180" daytime="18:28" gender="F" number="17" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1181" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3824" />
                    <RANKING order="2" place="2" resultid="2790" />
                    <RANKING order="3" place="3" resultid="1710" />
                    <RANKING order="4" place="4" resultid="3573" />
                    <RANKING order="5" place="5" resultid="3106" />
                    <RANKING order="6" place="6" resultid="2200" />
                    <RANKING order="7" place="7" resultid="2160" />
                    <RANKING order="8" place="8" resultid="1790" />
                    <RANKING order="9" place="9" resultid="3691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2919" />
                    <RANKING order="2" place="2" resultid="3290" />
                    <RANKING order="3" place="3" resultid="1679" />
                    <RANKING order="4" place="4" resultid="2375" />
                    <RANKING order="5" place="5" resultid="3137" />
                    <RANKING order="6" place="6" resultid="3239" />
                    <RANKING order="7" place="7" resultid="3814" />
                    <RANKING order="8" place="8" resultid="1534" />
                    <RANKING order="9" place="9" resultid="1515" />
                    <RANKING order="10" place="10" resultid="1742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1183" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2612" />
                    <RANKING order="2" place="2" resultid="1944" />
                    <RANKING order="3" place="3" resultid="2617" />
                    <RANKING order="4" place="4" resultid="1493" />
                    <RANKING order="5" place="5" resultid="3531" />
                    <RANKING order="6" place="-1" resultid="2533" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1184" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2878" />
                    <RANKING order="2" place="2" resultid="3412" />
                    <RANKING order="3" place="3" resultid="1753" />
                    <RANKING order="4" place="4" resultid="3514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2500" />
                    <RANKING order="2" place="2" resultid="1447" />
                    <RANKING order="3" place="3" resultid="3489" />
                    <RANKING order="4" place="4" resultid="1757" />
                    <RANKING order="5" place="5" resultid="1968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2980" />
                    <RANKING order="2" place="2" resultid="1471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3555" />
                    <RANKING order="2" place="2" resultid="2255" />
                    <RANKING order="3" place="3" resultid="2238" />
                    <RANKING order="4" place="4" resultid="3790" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4355" daytime="18:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4356" daytime="18:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4357" daytime="18:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4358" daytime="18:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4359" daytime="18:34" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1188" daytime="18:38" gender="M" number="18" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1189" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1655" />
                    <RANKING order="2" place="2" resultid="2766" />
                    <RANKING order="3" place="3" resultid="1527" />
                    <RANKING order="4" place="4" resultid="2172" />
                    <RANKING order="5" place="5" resultid="1595" />
                    <RANKING order="6" place="6" resultid="2363" />
                    <RANKING order="7" place="7" resultid="3594" />
                    <RANKING order="8" place="8" resultid="1962" />
                    <RANKING order="9" place="9" resultid="3436" />
                    <RANKING order="10" place="10" resultid="3366" />
                    <RANKING order="11" place="11" resultid="3072" />
                    <RANKING order="12" place="12" resultid="3233" />
                    <RANKING order="13" place="13" resultid="3228" />
                    <RANKING order="14" place="14" resultid="3590" />
                    <RANKING order="15" place="15" resultid="1523" />
                    <RANKING order="16" place="16" resultid="2225" />
                    <RANKING order="17" place="17" resultid="1804" />
                    <RANKING order="18" place="18" resultid="3696" />
                    <RANKING order="19" place="19" resultid="2166" />
                    <RANKING order="20" place="-1" resultid="2406" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3161" />
                    <RANKING order="2" place="2" resultid="1643" />
                    <RANKING order="3" place="3" resultid="2022" />
                    <RANKING order="4" place="4" resultid="3280" />
                    <RANKING order="5" place="5" resultid="3285" />
                    <RANKING order="6" place="6" resultid="3441" />
                    <RANKING order="7" place="7" resultid="3112" />
                    <RANKING order="8" place="8" resultid="2211" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3296" />
                    <RANKING order="2" place="2" resultid="2622" />
                    <RANKING order="3" place="3" resultid="1938" />
                    <RANKING order="4" place="4" resultid="3549" />
                    <RANKING order="5" place="5" resultid="3673" />
                    <RANKING order="6" place="6" resultid="1582" />
                    <RANKING order="7" place="7" resultid="1673" />
                    <RANKING order="8" place="8" resultid="3342" />
                    <RANKING order="9" place="-1" resultid="3451" />
                    <RANKING order="10" place="-1" resultid="3076" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2959" />
                    <RANKING order="2" place="2" resultid="1621" />
                    <RANKING order="3" place="3" resultid="2496" />
                    <RANKING order="4" place="4" resultid="2893" />
                    <RANKING order="5" place="5" resultid="1588" />
                    <RANKING order="6" place="6" resultid="2904" />
                    <RANKING order="7" place="7" resultid="1838" />
                    <RANKING order="8" place="8" resultid="2588" />
                    <RANKING order="9" place="9" resultid="3083" />
                    <RANKING order="10" place="10" resultid="3319" />
                    <RANKING order="11" place="11" resultid="1704" />
                    <RANKING order="12" place="12" resultid="3144" />
                    <RANKING order="13" place="13" resultid="2215" />
                    <RANKING order="14" place="14" resultid="3120" />
                    <RANKING order="15" place="15" resultid="1774" />
                    <RANKING order="16" place="16" resultid="3096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2555" />
                    <RANKING order="2" place="2" resultid="2297" />
                    <RANKING order="3" place="3" resultid="3197" />
                    <RANKING order="4" place="4" resultid="3361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2515" />
                    <RANKING order="2" place="2" resultid="1880" />
                    <RANKING order="3" place="3" resultid="1600" />
                    <RANKING order="4" place="4" resultid="3802" />
                    <RANKING order="5" place="5" resultid="1510" />
                    <RANKING order="6" place="6" resultid="3619" />
                    <RANKING order="7" place="7" resultid="1849" />
                    <RANKING order="8" place="8" resultid="3624" />
                    <RANKING order="9" place="9" resultid="3254" />
                    <RANKING order="10" place="10" resultid="1545" />
                    <RANKING order="11" place="11" resultid="3375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2561" />
                    <RANKING order="2" place="2" resultid="1467" />
                    <RANKING order="3" place="3" resultid="1560" />
                    <RANKING order="4" place="4" resultid="3000" />
                    <RANKING order="5" place="5" resultid="2654" />
                    <RANKING order="6" place="6" resultid="1905" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4360" daytime="18:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4361" daytime="18:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4362" daytime="18:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4363" daytime="18:44" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4364" daytime="18:46" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4365" daytime="18:46" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4366" daytime="18:48" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4367" daytime="18:50" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4368" daytime="18:52" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4369" daytime="18:54" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1196" daytime="18:56" gender="F" number="19" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1197" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3017" />
                    <RANKING order="2" place="2" resultid="3766" />
                    <RANKING order="3" place="3" resultid="2426" />
                    <RANKING order="4" place="4" resultid="3463" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4370" daytime="18:56" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1198" daytime="19:06" gender="F" number="20" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1199" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3019" />
                    <RANKING order="2" place="2" resultid="3747" />
                    <RANKING order="3" place="3" resultid="3464" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4371" daytime="19:06" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1200" daytime="19:18" gender="F" number="21" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1201" agemax="19" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3018" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4372" daytime="19:18" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1202" daytime="19:28" gender="F" number="22" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1203" agemax="-1" agemin="20" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1204" daytime="19:28" gender="M" number="23" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1205" agemax="14" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3030" />
                    <RANKING order="2" place="2" resultid="2431" />
                    <RANKING order="3" place="3" resultid="3771" />
                    <RANKING order="4" place="4" resultid="3244" />
                    <RANKING order="5" place="5" resultid="3470" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4373" daytime="19:28" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1206" daytime="19:38" gender="M" number="24" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1207" agemax="16" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3032" />
                    <RANKING order="2" place="2" resultid="2432" />
                    <RANKING order="3" place="3" resultid="3753" />
                    <RANKING order="4" place="4" resultid="3472" />
                    <RANKING order="5" place="5" resultid="2176" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4374" daytime="19:38" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1208" daytime="19:48" gender="M" number="25" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1209" agemax="19" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3031" />
                    <RANKING order="2" place="2" resultid="3752" />
                    <RANKING order="3" place="3" resultid="3471" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4375" daytime="19:48" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1210" daytime="20:00" gender="M" number="26" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1211" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2033" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4376" daytime="20:00" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-04-13" daytime="08:45" endtime="12:46" number="3" officialmeeting="08:00" warmupfrom="07:30" warmupuntil="08:30">
          <EVENTS>
            <EVENT eventid="1212" daytime="08:46" gender="F" number="27" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1213" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2953" />
                    <RANKING order="2" place="2" resultid="2778" />
                    <RANKING order="3" place="3" resultid="3826" />
                    <RANKING order="4" place="4" resultid="2803" />
                    <RANKING order="5" place="5" resultid="2370" />
                    <RANKING order="6" place="6" resultid="3168" />
                    <RANKING order="7" place="7" resultid="2872" />
                    <RANKING order="8" place="8" resultid="3643" />
                    <RANKING order="9" place="9" resultid="3575" />
                    <RANKING order="10" place="10" resultid="1711" />
                    <RANKING order="11" place="11" resultid="2791" />
                    <RANKING order="12" place="12" resultid="3210" />
                    <RANKING order="13" place="13" resultid="3107" />
                    <RANKING order="14" place="14" resultid="1792" />
                    <RANKING order="15" place="15" resultid="3693" />
                    <RANKING order="16" place="16" resultid="1441" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3291" />
                    <RANKING order="2" place="2" resultid="2529" />
                    <RANKING order="3" place="3" resultid="2920" />
                    <RANKING order="4" place="4" resultid="2995" />
                    <RANKING order="5" place="5" resultid="2376" />
                    <RANKING order="6" place="6" resultid="3661" />
                    <RANKING order="7" place="7" resultid="3138" />
                    <RANKING order="8" place="8" resultid="2867" />
                    <RANKING order="9" place="9" resultid="3815" />
                    <RANKING order="10" place="10" resultid="2418" />
                    <RANKING order="11" place="11" resultid="1517" />
                    <RANKING order="12" place="12" resultid="1536" />
                    <RANKING order="13" place="13" resultid="3447" />
                    <RANKING order="14" place="14" resultid="3116" />
                    <RANKING order="15" place="-1" resultid="3656" />
                    <RANKING order="16" place="-1" resultid="1743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2613" />
                    <RANKING order="2" place="2" resultid="1945" />
                    <RANKING order="3" place="3" resultid="2618" />
                    <RANKING order="4" place="4" resultid="3156" />
                    <RANKING order="5" place="5" resultid="2280" />
                    <RANKING order="6" place="6" resultid="1494" />
                    <RANKING order="7" place="7" resultid="3102" />
                    <RANKING order="8" place="-1" resultid="2534" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1216" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2447" />
                    <RANKING order="2" place="2" resultid="2880" />
                    <RANKING order="3" place="3" resultid="1755" />
                    <RANKING order="4" place="4" resultid="3516" />
                    <RANKING order="5" place="5" resultid="1418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2501" />
                    <RANKING order="2" place="2" resultid="3215" />
                    <RANKING order="3" place="3" resultid="1759" />
                    <RANKING order="4" place="4" resultid="1969" />
                    <RANKING order="5" place="-1" resultid="1448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2981" />
                    <RANKING order="2" place="2" resultid="1472" />
                    <RANKING order="3" place="3" resultid="3308" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3557" />
                    <RANKING order="2" place="2" resultid="3063" />
                    <RANKING order="3" place="3" resultid="2256" />
                    <RANKING order="4" place="4" resultid="3736" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4377" daytime="08:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4378" daytime="08:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4379" daytime="08:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4380" daytime="08:54" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4381" daytime="08:58" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4382" daytime="09:00" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4383" daytime="09:02" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4384" daytime="09:04" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4912" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1220" daytime="09:08" gender="M" number="28" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1221" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2322" />
                    <RANKING order="2" place="2" resultid="2767" />
                    <RANKING order="3" place="3" resultid="1656" />
                    <RANKING order="4" place="4" resultid="2814" />
                    <RANKING order="5" place="5" resultid="2899" />
                    <RANKING order="6" place="6" resultid="2831" />
                    <RANKING order="7" place="7" resultid="2310" />
                    <RANKING order="8" place="8" resultid="1596" />
                    <RANKING order="9" place="9" resultid="1528" />
                    <RANKING order="10" place="10" resultid="2407" />
                    <RANKING order="11" place="11" resultid="3595" />
                    <RANKING order="12" place="12" resultid="2364" />
                    <RANKING order="13" place="13" resultid="3600" />
                    <RANKING order="14" place="14" resultid="3186" />
                    <RANKING order="15" place="15" resultid="2205" />
                    <RANKING order="16" place="16" resultid="3437" />
                    <RANKING order="17" place="17" resultid="1844" />
                    <RANKING order="18" place="18" resultid="2783" />
                    <RANKING order="19" place="19" resultid="3649" />
                    <RANKING order="20" place="20" resultid="1861" />
                    <RANKING order="21" place="21" resultid="2226" />
                    <RANKING order="22" place="22" resultid="3234" />
                    <RANKING order="23" place="23" resultid="3697" />
                    <RANKING order="24" place="-1" resultid="1963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1222" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3162" />
                    <RANKING order="2" place="2" resultid="1926" />
                    <RANKING order="3" place="3" resultid="2721" />
                    <RANKING order="4" place="4" resultid="2661" />
                    <RANKING order="5" place="5" resultid="1644" />
                    <RANKING order="6" place="6" resultid="2023" />
                    <RANKING order="7" place="7" resultid="3281" />
                    <RANKING order="8" place="8" resultid="3442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1223" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1463" />
                    <RANKING order="2" place="2" resultid="3297" />
                    <RANKING order="3" place="3" resultid="2623" />
                    <RANKING order="4" place="4" resultid="3674" />
                    <RANKING order="5" place="5" resultid="1916" />
                    <RANKING order="6" place="6" resultid="2608" />
                    <RANKING order="7" place="7" resultid="3550" />
                    <RANKING order="8" place="8" resultid="2346" />
                    <RANKING order="9" place="9" resultid="1674" />
                    <RANKING order="10" place="10" resultid="3343" />
                    <RANKING order="11" place="11" resultid="3425" />
                    <RANKING order="12" place="-1" resultid="1583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1622" />
                    <RANKING order="2" place="2" resultid="2497" />
                    <RANKING order="3" place="3" resultid="2481" />
                    <RANKING order="4" place="4" resultid="2960" />
                    <RANKING order="5" place="5" resultid="2894" />
                    <RANKING order="6" place="6" resultid="2101" />
                    <RANKING order="7" place="7" resultid="2905" />
                    <RANKING order="8" place="8" resultid="1589" />
                    <RANKING order="9" place="9" resultid="3145" />
                    <RANKING order="10" place="10" resultid="3320" />
                    <RANKING order="11" place="11" resultid="2589" />
                    <RANKING order="12" place="12" resultid="3084" />
                    <RANKING order="13" place="13" resultid="1705" />
                    <RANKING order="14" place="14" resultid="2131" />
                    <RANKING order="15" place="15" resultid="2216" />
                    <RANKING order="16" place="16" resultid="1775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1225" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2556" />
                    <RANKING order="2" place="2" resultid="1407" />
                    <RANKING order="3" place="3" resultid="2510" />
                    <RANKING order="4" place="4" resultid="2299" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1226" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2516" />
                    <RANKING order="2" place="2" resultid="1601" />
                    <RANKING order="3" place="3" resultid="1881" />
                    <RANKING order="4" place="4" resultid="1850" />
                    <RANKING order="5" place="5" resultid="3803" />
                    <RANKING order="6" place="6" resultid="2232" />
                    <RANKING order="7" place="7" resultid="3255" />
                    <RANKING order="8" place="8" resultid="2196" />
                    <RANKING order="9" place="9" resultid="1546" />
                    <RANKING order="10" place="-1" resultid="3620" />
                    <RANKING order="11" place="-1" resultid="2471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1227" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2562" />
                    <RANKING order="2" place="2" resultid="1561" />
                    <RANKING order="3" place="3" resultid="1468" />
                    <RANKING order="4" place="4" resultid="2655" />
                    <RANKING order="5" place="5" resultid="1886" />
                    <RANKING order="6" place="6" resultid="1906" />
                    <RANKING order="7" place="-1" resultid="3001" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4385" daytime="09:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4386" daytime="09:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4387" daytime="09:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4388" daytime="09:16" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4389" daytime="09:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4390" daytime="09:22" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4391" daytime="09:24" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4392" daytime="09:26" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4393" daytime="09:28" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4394" daytime="09:32" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4395" daytime="09:34" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1228" daytime="09:36" gender="F" number="29" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1229" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2808" />
                    <RANKING order="2" place="2" resultid="1540" />
                    <RANKING order="3" place="3" resultid="1698" />
                    <RANKING order="4" place="4" resultid="3209" />
                    <RANKING order="5" place="5" resultid="2802" />
                    <RANKING order="6" place="6" resultid="3825" />
                    <RANKING order="7" place="7" resultid="2201" />
                    <RANKING order="8" place="8" resultid="3574" />
                    <RANKING order="9" place="9" resultid="1662" />
                    <RANKING order="10" place="10" resultid="3302" />
                    <RANKING order="11" place="11" resultid="1668" />
                    <RANKING order="12" place="12" resultid="1809" />
                    <RANKING order="13" place="13" resultid="2004" />
                    <RANKING order="14" place="14" resultid="2161" />
                    <RANKING order="15" place="15" resultid="1791" />
                    <RANKING order="16" place="16" resultid="3701" />
                    <RANKING order="17" place="17" resultid="1786" />
                    <RANKING order="18" place="18" resultid="1440" />
                    <RANKING order="19" place="19" resultid="3692" />
                    <RANKING order="20" place="-1" resultid="3422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2678" />
                    <RANKING order="2" place="2" resultid="1436" />
                    <RANKING order="3" place="3" resultid="1769" />
                    <RANKING order="4" place="4" resultid="1430" />
                    <RANKING order="5" place="5" resultid="1686" />
                    <RANKING order="6" place="6" resultid="3707" />
                    <RANKING order="7" place="7" resultid="2994" />
                    <RANKING order="8" place="8" resultid="2149" />
                    <RANKING order="9" place="9" resultid="2673" />
                    <RANKING order="10" place="10" resultid="1680" />
                    <RANKING order="11" place="11" resultid="3809" />
                    <RANKING order="12" place="12" resultid="3655" />
                    <RANKING order="13" place="13" resultid="2841" />
                    <RANKING order="14" place="14" resultid="1816" />
                    <RANKING order="15" place="15" resultid="2866" />
                    <RANKING order="16" place="16" resultid="3719" />
                    <RANKING order="17" place="17" resultid="3392" />
                    <RANKING order="18" place="18" resultid="3240" />
                    <RANKING order="19" place="19" resultid="1535" />
                    <RANKING order="20" place="20" resultid="3446" />
                    <RANKING order="21" place="21" resultid="1800" />
                    <RANKING order="22" place="22" resultid="1516" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2463" />
                    <RANKING order="2" place="2" resultid="3484" />
                    <RANKING order="3" place="3" resultid="3637" />
                    <RANKING order="4" place="4" resultid="1478" />
                    <RANKING order="5" place="5" resultid="1951" />
                    <RANKING order="6" place="6" resultid="3532" />
                    <RANKING order="7" place="7" resultid="3543" />
                    <RANKING order="8" place="8" resultid="3155" />
                    <RANKING order="9" place="9" resultid="2112" />
                    <RANKING order="10" place="10" resultid="1617" />
                    <RANKING order="11" place="11" resultid="2191" />
                    <RANKING order="12" place="12" resultid="3567" />
                    <RANKING order="13" place="13" resultid="3419" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1232" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3413" />
                    <RANKING order="2" place="2" resultid="1748" />
                    <RANKING order="3" place="3" resultid="2268" />
                    <RANKING order="4" place="4" resultid="2879" />
                    <RANKING order="5" place="5" resultid="3515" />
                    <RANKING order="6" place="6" resultid="1754" />
                    <RANKING order="7" place="7" resultid="1633" />
                    <RANKING order="8" place="8" resultid="3397" />
                    <RANKING order="9" place="9" resultid="3118" />
                    <RANKING order="10" place="10" resultid="1780" />
                    <RANKING order="11" place="-1" resultid="1993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3490" />
                    <RANKING order="2" place="2" resultid="1488" />
                    <RANKING order="3" place="3" resultid="1483" />
                    <RANKING order="4" place="4" resultid="1758" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1737" />
                    <RANKING order="2" place="2" resultid="2071" />
                    <RANKING order="3" place="3" resultid="2050" />
                    <RANKING order="4" place="4" resultid="3797" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1235" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3062" />
                    <RANKING order="2" place="2" resultid="3556" />
                    <RANKING order="3" place="3" resultid="3735" />
                    <RANKING order="4" place="4" resultid="3791" />
                    <RANKING order="5" place="5" resultid="2239" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4396" daytime="09:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4397" daytime="09:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4398" daytime="09:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4399" daytime="09:42" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4400" daytime="09:44" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4401" daytime="09:44" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4402" daytime="09:46" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4403" daytime="09:48" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4404" daytime="09:50" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4405" daytime="09:50" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1236" daytime="09:52" gender="M" number="30" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1237" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1650" />
                    <RANKING order="2" place="2" resultid="2860" />
                    <RANKING order="3" place="3" resultid="1795" />
                    <RANKING order="4" place="4" resultid="3192" />
                    <RANKING order="5" place="5" resultid="2815" />
                    <RANKING order="6" place="6" resultid="1529" />
                    <RANKING order="7" place="7" resultid="2173" />
                    <RANKING order="8" place="8" resultid="3631" />
                    <RANKING order="9" place="9" resultid="3579" />
                    <RANKING order="10" place="10" resultid="3601" />
                    <RANKING order="11" place="11" resultid="2394" />
                    <RANKING order="12" place="12" resultid="2206" />
                    <RANKING order="13" place="13" resultid="3685" />
                    <RANKING order="14" place="14" resultid="3174" />
                    <RANKING order="15" place="15" resultid="1855" />
                    <RANKING order="16" place="16" resultid="2909" />
                    <RANKING order="17" place="17" resultid="1657" />
                    <RANKING order="18" place="18" resultid="1964" />
                    <RANKING order="19" place="19" resultid="2819" />
                    <RANKING order="20" place="20" resultid="3073" />
                    <RANKING order="21" place="21" resultid="1805" />
                    <RANKING order="22" place="22" resultid="1524" />
                    <RANKING order="23" place="23" resultid="2784" />
                    <RANKING order="24" place="24" resultid="1692" />
                    <RANKING order="25" place="25" resultid="1922" />
                    <RANKING order="26" place="26" resultid="3591" />
                    <RANKING order="27" place="27" resultid="3235" />
                    <RANKING order="28" place="28" resultid="1845" />
                    <RANKING order="29" place="29" resultid="2227" />
                    <RANKING order="30" place="30" resultid="2167" />
                    <RANKING order="31" place="31" resultid="3698" />
                    <RANKING order="32" place="-1" resultid="3368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1238" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1571" />
                    <RANKING order="2" place="2" resultid="2931" />
                    <RANKING order="3" place="3" resultid="2848" />
                    <RANKING order="4" place="4" resultid="2662" />
                    <RANKING order="5" place="5" resultid="2155" />
                    <RANKING order="6" place="6" resultid="2703" />
                    <RANKING order="7" place="7" resultid="2143" />
                    <RANKING order="8" place="8" resultid="3585" />
                    <RANKING order="9" place="9" resultid="2732" />
                    <RANKING order="10" place="10" resultid="1716" />
                    <RANKING order="11" place="11" resultid="2028" />
                    <RANKING order="12" place="12" resultid="3679" />
                    <RANKING order="13" place="13" resultid="3221" />
                    <RANKING order="14" place="14" resultid="1984" />
                    <RANKING order="15" place="15" resultid="2016" />
                    <RANKING order="16" place="15" resultid="2024" />
                    <RANKING order="17" place="17" resultid="3443" />
                    <RANKING order="18" place="18" resultid="3113" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1239" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2486" />
                    <RANKING order="2" place="2" resultid="1455" />
                    <RANKING order="3" place="3" resultid="1939" />
                    <RANKING order="4" place="4" resultid="1565" />
                    <RANKING order="5" place="5" resultid="2972" />
                    <RANKING order="6" place="6" resultid="2539" />
                    <RANKING order="7" place="7" resultid="3526" />
                    <RANKING order="8" place="8" resultid="3520" />
                    <RANKING order="9" place="9" resultid="1500" />
                    <RANKING order="10" place="10" resultid="3551" />
                    <RANKING order="11" place="11" resultid="1980" />
                    <RANKING order="12" place="12" resultid="1628" />
                    <RANKING order="13" place="13" resultid="1917" />
                    <RANKING order="14" place="14" resultid="1506" />
                    <RANKING order="15" place="15" resultid="3713" />
                    <RANKING order="16" place="16" resultid="3067" />
                    <RANKING order="17" place="17" resultid="3344" />
                    <RANKING order="18" place="18" resultid="3077" />
                    <RANKING order="19" place="19" resultid="3080" />
                    <RANKING order="20" place="20" resultid="2009" />
                    <RANKING order="21" place="21" resultid="2603" />
                    <RANKING order="22" place="22" resultid="1675" />
                    <RANKING order="23" place="23" resultid="2220" />
                    <RANKING order="24" place="-1" resultid="2650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1240" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2961" />
                    <RANKING order="2" place="2" resultid="2584" />
                    <RANKING order="3" place="3" resultid="2914" />
                    <RANKING order="4" place="4" resultid="3538" />
                    <RANKING order="5" place="5" resultid="1577" />
                    <RANKING order="6" place="6" resultid="2064" />
                    <RANKING order="7" place="7" resultid="1839" />
                    <RANKING order="8" place="8" resultid="3508" />
                    <RANKING order="9" place="9" resultid="2943" />
                    <RANKING order="10" place="10" resultid="2593" />
                    <RANKING order="11" place="11" resultid="2388" />
                    <RANKING order="12" place="12" resultid="1866" />
                    <RANKING order="13" place="13" resultid="2578" />
                    <RANKING order="14" place="14" resultid="2644" />
                    <RANKING order="15" place="15" resultid="3097" />
                    <RANKING order="16" place="16" resultid="2572" />
                    <RANKING order="17" place="17" resultid="1998" />
                    <RANKING order="18" place="18" resultid="3150" />
                    <RANKING order="19" place="19" resultid="1989" />
                    <RANKING order="20" place="20" resultid="1764" />
                    <RANKING order="21" place="21" resultid="3460" />
                    <RANKING order="22" place="22" resultid="2217" />
                    <RANKING order="23" place="23" resultid="3121" />
                    <RANKING order="24" place="24" resultid="3085" />
                    <RANKING order="25" place="25" resultid="1706" />
                    <RANKING order="26" place="26" resultid="1776" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2550" />
                    <RANKING order="2" place="2" resultid="3496" />
                    <RANKING order="3" place="3" resultid="3407" />
                    <RANKING order="4" place="4" resultid="3271" />
                    <RANKING order="5" place="5" resultid="3740" />
                    <RANKING order="6" place="6" resultid="3198" />
                    <RANKING order="7" place="7" resultid="3204" />
                    <RANKING order="8" place="8" resultid="3431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2984" />
                    <RANKING order="2" place="2" resultid="3014" />
                    <RANKING order="3" place="3" resultid="3625" />
                    <RANKING order="4" place="4" resultid="1556" />
                    <RANKING order="5" place="5" resultid="1882" />
                    <RANKING order="6" place="6" resultid="3332" />
                    <RANKING order="7" place="7" resultid="2083" />
                    <RANKING order="8" place="8" resultid="1511" />
                    <RANKING order="9" place="9" resultid="3621" />
                    <RANKING order="10" place="10" resultid="1639" />
                    <RANKING order="11" place="11" resultid="1606" />
                    <RANKING order="12" place="12" resultid="1896" />
                    <RANKING order="13" place="13" resultid="2188" />
                    <RANKING order="14" place="14" resultid="3804" />
                    <RANKING order="15" place="15" resultid="2352" />
                    <RANKING order="16" place="16" resultid="3092" />
                    <RANKING order="17" place="17" resultid="2567" />
                    <RANKING order="18" place="-1" resultid="1547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1243" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2656" />
                    <RANKING order="2" place="2" resultid="2054" />
                    <RANKING order="3" place="3" resultid="1828" />
                    <RANKING order="4" place="4" resultid="2925" />
                    <RANKING order="5" place="5" resultid="1413" />
                    <RANKING order="6" place="6" resultid="3745" />
                    <RANKING order="7" place="7" resultid="2076" />
                    <RANKING order="8" place="8" resultid="1910" />
                    <RANKING order="9" place="9" resultid="3131" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4406" daytime="09:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4407" daytime="09:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4408" daytime="09:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4409" daytime="09:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4410" daytime="10:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4411" daytime="10:02" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4412" daytime="10:04" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4413" daytime="10:04" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4414" daytime="10:06" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4415" daytime="10:08" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4416" daytime="10:10" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4417" daytime="10:10" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="4418" daytime="10:12" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="4419" daytime="10:14" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="4420" daytime="10:16" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="4421" daytime="10:16" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="4422" daytime="10:18" number="17" order="17" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1244" daytime="10:20" gender="X" number="31" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1245" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3047" />
                    <RANKING order="2" place="2" resultid="2041" />
                    <RANKING order="3" place="3" resultid="3765" />
                    <RANKING order="4" place="4" resultid="1551" />
                    <RANKING order="5" place="5" resultid="1731" />
                    <RANKING order="6" place="6" resultid="3760" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4423" daytime="10:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1246" daytime="10:26" gender="X" number="32" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1247" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3046" />
                    <RANKING order="2" place="2" resultid="2443" />
                    <RANKING order="3" place="3" resultid="2185" />
                    <RANKING order="4" place="4" resultid="3479" />
                    <RANKING order="5" place="5" resultid="3759" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4424" daytime="10:26" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1248" daytime="10:34" gender="X" number="33" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1249" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3045" />
                    <RANKING order="2" place="2" resultid="1451" />
                    <RANKING order="3" place="3" resultid="2184" />
                    <RANKING order="4" place="4" resultid="3758" />
                    <RANKING order="5" place="5" resultid="1550" />
                    <RANKING order="6" place="6" resultid="2442" />
                    <RANKING order="7" place="7" resultid="3478" />
                    <RANKING order="8" place="8" resultid="2040" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4425" daytime="10:34" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1250" daytime="10:40" gender="F" number="34" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1251" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2826" />
                    <RANKING order="2" place="2" resultid="2334" />
                    <RANKING order="3" place="3" resultid="2399" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1252" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2725" />
                    <RANKING order="2" place="2" resultid="2137" />
                    <RANKING order="3" place="3" resultid="2715" />
                    <RANKING order="4" place="4" resultid="2685" />
                    <RANKING order="5" place="5" resultid="3613" />
                    <RANKING order="6" place="6" resultid="2736" />
                    <RANKING order="7" place="7" resultid="3325" />
                    <RANKING order="8" place="8" resultid="3139" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1253" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2523" />
                    <RANKING order="2" place="2" resultid="2451" />
                    <RANKING order="3" place="3" resultid="2628" />
                    <RANKING order="4" place="4" resultid="3533" />
                    <RANKING order="5" place="5" resultid="1611" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1254" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2046" />
                    <RANKING order="2" place="2" resultid="3354" />
                    <RANKING order="3" place="3" resultid="3264" />
                    <RANKING order="4" place="4" resultid="1833" />
                    <RANKING order="5" place="-1" resultid="2966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1255" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2544" />
                    <RANKING order="2" place="2" resultid="1424" />
                    <RANKING order="3" place="3" resultid="2245" />
                    <RANKING order="4" place="4" resultid="3216" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1256" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1257" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2937" />
                    <RANKING order="2" place="2" resultid="3004" />
                    <RANKING order="3" place="3" resultid="2976" />
                    <RANKING order="4" place="4" resultid="3349" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4426" daytime="10:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4427" daytime="10:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4428" daytime="11:06" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1258" daytime="11:18" gender="M" number="35" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1259" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2772" />
                    <RANKING order="2" place="2" resultid="2754" />
                    <RANKING order="3" place="3" resultid="2795" />
                    <RANKING order="4" place="4" resultid="3367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2697" />
                    <RANKING order="2" place="2" resultid="2709" />
                    <RANKING order="3" place="3" resultid="2743" />
                    <RANKING order="4" place="4" resultid="3607" />
                    <RANKING order="5" place="5" resultid="3667" />
                    <RANKING order="6" place="6" resultid="2292" />
                    <RANKING order="7" place="7" resultid="3282" />
                    <RANKING order="8" place="-1" resultid="2382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1261" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2262" />
                    <RANKING order="2" place="2" resultid="3525" />
                    <RANKING order="3" place="3" resultid="3276" />
                    <RANKING order="4" place="4" resultid="2639" />
                    <RANKING order="5" place="5" resultid="1505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1262" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2854" />
                    <RANKING order="2" place="2" resultid="2358" />
                    <RANKING order="3" place="3" resultid="2125" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3731" />
                    <RANKING order="2" place="2" resultid="2107" />
                    <RANKING order="3" place="3" resultid="3362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1265" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3337" />
                    <RANKING order="2" place="2" resultid="1901" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4430" daytime="11:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4431" daytime="11:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4432" daytime="12:04" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-04-13" daytime="16:15" number="4" officialmeeting="16:30" warmupfrom="15:00" warmupuntil="16:00">
          <EVENTS>
            <EVENT eventid="1266" daytime="16:16" gender="F" number="36" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1267" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2884" />
                    <RANKING order="2" place="2" resultid="2827" />
                    <RANKING order="3" place="3" resultid="2329" />
                    <RANKING order="4" place="4" resultid="2779" />
                    <RANKING order="5" place="5" resultid="2955" />
                    <RANKING order="6" place="6" resultid="2413" />
                    <RANKING order="7" place="7" resultid="2371" />
                    <RANKING order="8" place="8" resultid="3108" />
                    <RANKING order="9" place="-1" resultid="1712" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1268" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2726" />
                    <RANKING order="2" place="2" resultid="2274" />
                    <RANKING order="3" place="3" resultid="2530" />
                    <RANKING order="4" place="4" resultid="3292" />
                    <RANKING order="5" place="5" resultid="3327" />
                    <RANKING order="6" place="6" resultid="1438" />
                    <RANKING order="7" place="7" resultid="2843" />
                    <RANKING order="8" place="8" resultid="2868" />
                    <RANKING order="9" place="9" resultid="2150" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1269" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3157" />
                    <RANKING order="2" place="2" resultid="2619" />
                    <RANKING order="3" place="3" resultid="2614" />
                    <RANKING order="4" place="4" resultid="2281" />
                    <RANKING order="5" place="5" resultid="1947" />
                    <RANKING order="6" place="6" resultid="3103" />
                    <RANKING order="7" place="-1" resultid="2629" />
                    <RANKING order="8" place="-1" resultid="2193" />
                    <RANKING order="9" place="-1" resultid="2535" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1270" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2457" />
                    <RANKING order="2" place="2" resultid="2448" />
                    <RANKING order="3" place="3" resultid="2270" />
                    <RANKING order="4" place="4" resultid="1419" />
                    <RANKING order="5" place="5" resultid="3399" />
                    <RANKING order="6" place="-1" resultid="2317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1271" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1449" />
                    <RANKING order="2" place="2" resultid="3217" />
                    <RANKING order="3" place="3" resultid="1970" />
                    <RANKING order="4" place="-1" resultid="2502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1272" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1473" />
                    <RANKING order="2" place="2" resultid="3309" />
                    <RANKING order="3" place="3" resultid="3315" />
                    <RANKING order="4" place="4" resultid="3089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1273" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3350" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4434" daytime="16:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4435" daytime="16:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4436" daytime="16:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4437" daytime="16:28" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4438" daytime="16:32" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4439" daytime="16:36" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1274" daytime="16:42" gender="M" number="37" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1275" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2323" />
                    <RANKING order="2" place="2" resultid="2311" />
                    <RANKING order="3" place="3" resultid="2832" />
                    <RANKING order="4" place="4" resultid="2395" />
                    <RANKING order="5" place="5" resultid="2816" />
                    <RANKING order="6" place="6" resultid="2796" />
                    <RANKING order="7" place="7" resultid="3596" />
                    <RANKING order="8" place="8" resultid="2900" />
                    <RANKING order="9" place="9" resultid="1658" />
                    <RANKING order="10" place="10" resultid="2820" />
                    <RANKING order="11" place="11" resultid="3187" />
                    <RANKING order="12" place="12" resultid="1597" />
                    <RANKING order="13" place="13" resultid="3127" />
                    <RANKING order="14" place="14" resultid="3438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2287" />
                    <RANKING order="2" place="2" resultid="1572" />
                    <RANKING order="3" place="3" resultid="1927" />
                    <RANKING order="4" place="4" resultid="2722" />
                    <RANKING order="5" place="5" resultid="3163" />
                    <RANKING order="6" place="6" resultid="2733" />
                    <RANKING order="7" place="7" resultid="3287" />
                    <RANKING order="8" place="-1" resultid="2698" />
                    <RANKING order="9" place="-1" resultid="2383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1877" />
                    <RANKING order="2" place="2" resultid="1464" />
                    <RANKING order="3" place="3" resultid="3675" />
                    <RANKING order="4" place="4" resultid="2540" />
                    <RANKING order="5" place="5" resultid="3277" />
                    <RANKING order="6" place="6" resultid="2347" />
                    <RANKING order="7" place="7" resultid="2624" />
                    <RANKING order="8" place="8" resultid="1918" />
                    <RANKING order="9" place="9" resultid="1981" />
                    <RANKING order="10" place="10" resultid="1584" />
                    <RANKING order="11" place="11" resultid="2120" />
                    <RANKING order="12" place="12" resultid="1676" />
                    <RANKING order="13" place="13" resultid="3426" />
                    <RANKING order="14" place="-1" resultid="2263" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1278" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2251" />
                    <RANKING order="2" place="2" resultid="2482" />
                    <RANKING order="3" place="3" resultid="2492" />
                    <RANKING order="4" place="4" resultid="2962" />
                    <RANKING order="5" place="5" resultid="1623" />
                    <RANKING order="6" place="6" resultid="2895" />
                    <RANKING order="7" place="7" resultid="3151" />
                    <RANKING order="8" place="8" resultid="1590" />
                    <RANKING order="9" place="9" resultid="3146" />
                    <RANKING order="10" place="10" resultid="3098" />
                    <RANKING order="11" place="-1" resultid="3321" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2511" />
                    <RANKING order="2" place="2" resultid="1408" />
                    <RANKING order="3" place="3" resultid="2557" />
                    <RANKING order="4" place="4" resultid="2300" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1280" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2233" />
                    <RANKING order="2" place="2" resultid="1602" />
                    <RANKING order="3" place="3" resultid="1607" />
                    <RANKING order="4" place="4" resultid="3256" />
                    <RANKING order="5" place="5" resultid="2197" />
                    <RANKING order="6" place="-1" resultid="3377" />
                    <RANKING order="7" place="-1" resultid="2472" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2657" />
                    <RANKING order="2" place="2" resultid="1887" />
                    <RANKING order="3" place="3" resultid="3338" />
                    <RANKING order="4" place="4" resultid="2090" />
                    <RANKING order="5" place="5" resultid="1907" />
                    <RANKING order="6" place="-1" resultid="2563" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4440" daytime="16:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4441" daytime="16:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4442" daytime="16:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4443" daytime="16:54" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4444" daytime="16:58" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4445" daytime="17:02" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4446" daytime="17:06" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4447" daytime="17:10" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4448" daytime="17:14" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1282" daytime="17:18" gender="F" number="38" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1283" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2809" />
                    <RANKING order="2" place="2" resultid="2804" />
                    <RANKING order="3" place="3" resultid="2335" />
                    <RANKING order="4" place="4" resultid="2400" />
                    <RANKING order="5" place="5" resultid="2873" />
                    <RANKING order="6" place="6" resultid="2954" />
                    <RANKING order="7" place="7" resultid="3819" />
                    <RANKING order="8" place="8" resultid="3211" />
                    <RANKING order="9" place="9" resultid="3169" />
                    <RANKING order="10" place="10" resultid="2792" />
                    <RANKING order="11" place="11" resultid="3303" />
                    <RANKING order="12" place="12" resultid="1663" />
                    <RANKING order="13" place="13" resultid="3644" />
                    <RANKING order="14" place="14" resultid="2005" />
                    <RANKING order="15" place="15" resultid="3702" />
                    <RANKING order="16" place="16" resultid="1442" />
                    <RANKING order="17" place="17" resultid="2162" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1284" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2679" />
                    <RANKING order="2" place="2" resultid="2691" />
                    <RANKING order="3" place="3" resultid="3614" />
                    <RANKING order="4" place="4" resultid="1687" />
                    <RANKING order="5" place="5" resultid="2377" />
                    <RANKING order="6" place="6" resultid="2716" />
                    <RANKING order="7" place="7" resultid="2996" />
                    <RANKING order="8" place="8" resultid="2138" />
                    <RANKING order="9" place="9" resultid="3708" />
                    <RANKING order="10" place="10" resultid="3662" />
                    <RANKING order="11" place="11" resultid="1437" />
                    <RANKING order="12" place="12" resultid="3657" />
                    <RANKING order="13" place="13" resultid="3326" />
                    <RANKING order="14" place="14" resultid="2921" />
                    <RANKING order="15" place="15" resultid="2737" />
                    <RANKING order="16" place="16" resultid="2419" />
                    <RANKING order="17" place="17" resultid="1817" />
                    <RANKING order="18" place="18" resultid="2842" />
                    <RANKING order="19" place="19" resultid="3720" />
                    <RANKING order="20" place="20" resultid="1744" />
                    <RANKING order="21" place="21" resultid="3725" />
                    <RANKING order="22" place="22" resultid="3393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3485" />
                    <RANKING order="2" place="2" resultid="2524" />
                    <RANKING order="3" place="3" resultid="2464" />
                    <RANKING order="4" place="4" resultid="2452" />
                    <RANKING order="5" place="5" resultid="3638" />
                    <RANKING order="6" place="6" resultid="3544" />
                    <RANKING order="7" place="7" resultid="3568" />
                    <RANKING order="8" place="8" resultid="1952" />
                    <RANKING order="9" place="9" resultid="3534" />
                    <RANKING order="10" place="10" resultid="2113" />
                    <RANKING order="11" place="11" resultid="2192" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1286" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1749" />
                    <RANKING order="2" place="2" resultid="3414" />
                    <RANKING order="3" place="3" resultid="3355" />
                    <RANKING order="4" place="4" resultid="2269" />
                    <RANKING order="5" place="5" resultid="1834" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1287" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2545" />
                    <RANKING order="2" place="2" resultid="2059" />
                    <RANKING order="3" place="3" resultid="1425" />
                    <RANKING order="4" place="4" resultid="1975" />
                    <RANKING order="5" place="5" resultid="1760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3502" />
                    <RANKING order="2" place="2" resultid="3371" />
                    <RANKING order="3" place="-1" resultid="2072" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1289" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2938" />
                    <RANKING order="2" place="2" resultid="2240" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4449" daytime="17:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4450" daytime="17:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4451" daytime="17:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4452" daytime="17:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4453" daytime="17:34" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4454" daytime="17:38" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4455" daytime="17:42" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4456" daytime="17:44" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4457" daytime="17:48" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4977" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1290" daytime="17:52" gender="M" number="39" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1291" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2861" />
                    <RANKING order="2" place="2" resultid="2305" />
                    <RANKING order="3" place="3" resultid="2755" />
                    <RANKING order="4" place="4" resultid="2760" />
                    <RANKING order="5" place="5" resultid="3632" />
                    <RANKING order="6" place="6" resultid="3602" />
                    <RANKING order="7" place="7" resultid="2341" />
                    <RANKING order="8" place="8" resultid="2207" />
                    <RANKING order="9" place="9" resultid="2408" />
                    <RANKING order="10" place="10" resultid="2773" />
                    <RANKING order="11" place="11" resultid="2910" />
                    <RANKING order="12" place="12" resultid="3175" />
                    <RANKING order="13" place="13" resultid="2174" />
                    <RANKING order="14" place="14" resultid="3650" />
                    <RANKING order="15" place="15" resultid="3193" />
                    <RANKING order="16" place="16" resultid="2365" />
                    <RANKING order="17" place="17" resultid="1923" />
                    <RANKING order="18" place="18" resultid="1846" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2849" />
                    <RANKING order="2" place="2" resultid="2704" />
                    <RANKING order="3" place="3" resultid="2932" />
                    <RANKING order="4" place="4" resultid="2744" />
                    <RANKING order="5" place="5" resultid="2286" />
                    <RANKING order="6" place="6" resultid="2710" />
                    <RANKING order="7" place="7" resultid="2663" />
                    <RANKING order="8" place="8" resultid="3586" />
                    <RANKING order="9" place="9" resultid="2667" />
                    <RANKING order="10" place="10" resultid="3668" />
                    <RANKING order="11" place="11" resultid="3608" />
                    <RANKING order="12" place="12" resultid="2293" />
                    <RANKING order="13" place="13" resultid="1717" />
                    <RANKING order="14" place="14" resultid="2017" />
                    <RANKING order="15" place="15" resultid="3283" />
                    <RANKING order="16" place="16" resultid="3680" />
                    <RANKING order="17" place="17" resultid="3222" />
                    <RANKING order="18" place="18" resultid="2029" />
                    <RANKING order="19" place="-1" resultid="1958" />
                    <RANKING order="20" place="-1" resultid="2156" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1293" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1566" />
                    <RANKING order="2" place="2" resultid="1456" />
                    <RANKING order="3" place="3" resultid="2487" />
                    <RANKING order="4" place="4" resultid="3527" />
                    <RANKING order="5" place="5" resultid="2609" />
                    <RANKING order="6" place="6" resultid="3552" />
                    <RANKING order="7" place="7" resultid="3180" />
                    <RANKING order="8" place="8" resultid="3345" />
                    <RANKING order="9" place="9" resultid="3714" />
                    <RANKING order="10" place="10" resultid="1934" />
                    <RANKING order="11" place="11" resultid="2010" />
                    <RANKING order="12" place="12" resultid="2221" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1294" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2855" />
                    <RANKING order="2" place="2" resultid="2389" />
                    <RANKING order="3" place="3" resultid="2915" />
                    <RANKING order="4" place="4" resultid="3539" />
                    <RANKING order="5" place="5" resultid="2102" />
                    <RANKING order="6" place="6" resultid="2359" />
                    <RANKING order="7" place="7" resultid="2594" />
                    <RANKING order="8" place="8" resultid="1840" />
                    <RANKING order="9" place="9" resultid="3509" />
                    <RANKING order="10" place="10" resultid="2126" />
                    <RANKING order="11" place="11" resultid="2132" />
                    <RANKING order="12" place="12" resultid="1999" />
                    <RANKING order="13" place="13" resultid="2065" />
                    <RANKING order="14" place="14" resultid="3461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1295" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2551" />
                    <RANKING order="2" place="2" resultid="3497" />
                    <RANKING order="3" place="3" resultid="3408" />
                    <RANKING order="4" place="4" resultid="3741" />
                    <RANKING order="5" place="5" resultid="2108" />
                    <RANKING order="6" place="6" resultid="3732" />
                    <RANKING order="7" place="7" resultid="3455" />
                    <RANKING order="8" place="8" resultid="3205" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1296" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2505" />
                    <RANKING order="2" place="2" resultid="2985" />
                    <RANKING order="3" place="3" resultid="2519" />
                    <RANKING order="4" place="4" resultid="2517" />
                    <RANKING order="5" place="5" resultid="3561" />
                    <RANKING order="6" place="6" resultid="1557" />
                    <RANKING order="7" place="7" resultid="2749" />
                    <RANKING order="8" place="8" resultid="3015" />
                    <RANKING order="9" place="9" resultid="2084" />
                    <RANKING order="10" place="10" resultid="3626" />
                    <RANKING order="11" place="11" resultid="2096" />
                    <RANKING order="12" place="12" resultid="3259" />
                    <RANKING order="13" place="13" resultid="1897" />
                    <RANKING order="14" place="14" resultid="1640" />
                    <RANKING order="15" place="15" resultid="3805" />
                    <RANKING order="16" place="16" resultid="2568" />
                    <RANKING order="17" place="17" resultid="3376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1297" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2926" />
                    <RANKING order="2" place="2" resultid="1911" />
                    <RANKING order="3" place="3" resultid="1892" />
                    <RANKING order="4" place="4" resultid="1902" />
                    <RANKING order="5" place="5" resultid="3132" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4458" daytime="17:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4459" daytime="17:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4460" daytime="18:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4461" daytime="18:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4462" daytime="18:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4463" daytime="18:12" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4464" daytime="18:16" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4465" daytime="18:18" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4466" daytime="18:22" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="4467" daytime="18:26" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="4468" daytime="18:28" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="4469" daytime="18:32" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1298" daytime="18:36" gender="F" number="40" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1299" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1541" />
                    <RANKING order="2" place="2" resultid="2948" />
                    <RANKING order="3" place="3" resultid="1699" />
                    <RANKING order="4" place="4" resultid="3304" />
                    <RANKING order="5" place="5" resultid="2202" />
                    <RANKING order="6" place="6" resultid="1669" />
                    <RANKING order="7" place="7" resultid="3645" />
                    <RANKING order="8" place="8" resultid="1810" />
                    <RANKING order="9" place="9" resultid="1443" />
                    <RANKING order="10" place="10" resultid="3703" />
                    <RANKING order="11" place="11" resultid="2163" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1300" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3810" />
                    <RANKING order="2" place="2" resultid="1770" />
                    <RANKING order="3" place="3" resultid="2674" />
                    <RANKING order="4" place="4" resultid="1681" />
                    <RANKING order="5" place="5" resultid="3726" />
                    <RANKING order="6" place="6" resultid="1518" />
                    <RANKING order="7" place="7" resultid="3241" />
                    <RANKING order="8" place="8" resultid="3387" />
                    <RANKING order="9" place="9" resultid="1801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1301" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1872" />
                    <RANKING order="2" place="2" resultid="1479" />
                    <RANKING order="3" place="3" resultid="3639" />
                    <RANKING order="4" place="4" resultid="1612" />
                    <RANKING order="5" place="5" resultid="3545" />
                    <RANKING order="6" place="6" resultid="1495" />
                    <RANKING order="7" place="7" resultid="3420" />
                    <RANKING order="8" place="8" resultid="1618" />
                    <RANKING order="9" place="9" resultid="1946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1302" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2967" />
                    <RANKING order="2" place="2" resultid="3265" />
                    <RANKING order="3" place="3" resultid="1634" />
                    <RANKING order="4" place="4" resultid="3398" />
                    <RANKING order="5" place="5" resultid="1781" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1303" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3491" />
                    <RANKING order="2" place="2" resultid="1489" />
                    <RANKING order="3" place="3" resultid="1484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1304" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1738" />
                    <RANKING order="2" place="2" resultid="2051" />
                    <RANKING order="3" place="3" resultid="3798" />
                    <RANKING order="4" place="4" resultid="3314" />
                    <RANKING order="5" place="5" resultid="3088" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1305" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2257" />
                    <RANKING order="2" place="2" resultid="3792" />
                    <RANKING order="3" place="3" resultid="3381" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4470" daytime="18:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4471" daytime="18:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4472" daytime="18:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4473" daytime="18:44" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4474" daytime="18:46" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4475" daytime="18:48" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1306" daytime="18:50" gender="M" number="41" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1307" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1651" />
                    <RANKING order="2" place="2" resultid="1796" />
                    <RANKING order="3" place="3" resultid="3580" />
                    <RANKING order="4" place="4" resultid="1530" />
                    <RANKING order="5" place="5" resultid="1856" />
                    <RANKING order="6" place="6" resultid="3369" />
                    <RANKING order="7" place="7" resultid="3126" />
                    <RANKING order="8" place="8" resultid="3686" />
                    <RANKING order="9" place="9" resultid="3229" />
                    <RANKING order="10" place="10" resultid="1806" />
                    <RANKING order="11" place="11" resultid="1862" />
                    <RANKING order="12" place="12" resultid="1693" />
                    <RANKING order="13" place="13" resultid="3236" />
                    <RANKING order="14" place="14" resultid="2168" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1308" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2144" />
                    <RANKING order="2" place="2" resultid="1645" />
                    <RANKING order="3" place="3" resultid="3223" />
                    <RANKING order="4" place="4" resultid="3286" />
                    <RANKING order="5" place="5" resultid="1985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1309" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3009" />
                    <RANKING order="2" place="2" resultid="1457" />
                    <RANKING order="3" place="3" resultid="3298" />
                    <RANKING order="4" place="4" resultid="3521" />
                    <RANKING order="5" place="5" resultid="1940" />
                    <RANKING order="6" place="6" resultid="3181" />
                    <RANKING order="7" place="7" resultid="2119" />
                    <RANKING order="8" place="8" resultid="3068" />
                    <RANKING order="9" place="9" resultid="2011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1310" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2476" />
                    <RANKING order="2" place="2" resultid="2645" />
                    <RANKING order="3" place="3" resultid="3786" />
                    <RANKING order="4" place="4" resultid="2598" />
                    <RANKING order="5" place="5" resultid="2066" />
                    <RANKING order="6" place="5" resultid="2579" />
                    <RANKING order="7" place="7" resultid="1578" />
                    <RANKING order="8" place="8" resultid="2573" />
                    <RANKING order="9" place="9" resultid="1867" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1311" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2990" />
                    <RANKING order="2" place="2" resultid="3199" />
                    <RANKING order="3" place="3" resultid="3432" />
                    <RANKING order="4" place="4" resultid="3206" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1312" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3562" />
                    <RANKING order="2" place="2" resultid="1883" />
                    <RANKING order="3" place="3" resultid="1512" />
                    <RANKING order="4" place="4" resultid="2353" />
                    <RANKING order="5" place="5" resultid="1851" />
                    <RANKING order="6" place="6" resultid="2189" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1313" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2837" />
                    <RANKING order="2" place="2" resultid="3746" />
                    <RANKING order="3" place="3" resultid="1822" />
                    <RANKING order="4" place="4" resultid="2423" />
                    <RANKING order="5" place="5" resultid="2077" />
                    <RANKING order="6" place="6" resultid="2055" />
                    <RANKING order="7" place="7" resultid="2089" />
                    <RANKING order="8" place="8" resultid="1829" />
                    <RANKING order="9" place="9" resultid="3133" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4476" daytime="18:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4477" daytime="18:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4478" daytime="18:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4479" daytime="18:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4480" daytime="19:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4481" daytime="19:02" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4482" daytime="19:04" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1314" daytime="19:06" gender="F" number="42" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1315" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3020" />
                    <RANKING order="2" place="2" resultid="2427" />
                    <RANKING order="3" place="-1" resultid="3048" />
                    <RANKING order="4" place="-1" resultid="1719" />
                    <RANKING order="5" place="-1" resultid="3767" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4483" daytime="19:06" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1316" daytime="19:14" gender="F" number="43" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1317" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3021" />
                    <RANKING order="2" place="2" resultid="3049" />
                    <RANKING order="3" place="3" resultid="2428" />
                    <RANKING order="4" place="4" resultid="3768" />
                    <RANKING order="5" place="5" resultid="3827" />
                    <RANKING order="6" place="6" resultid="3465" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4484" daytime="19:14" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1318" daytime="19:20" gender="F" number="44" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1319" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3023" />
                    <RANKING order="2" place="2" resultid="3748" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4485" daytime="19:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1320" daytime="19:26" gender="F" number="45" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1321" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3022" />
                    <RANKING order="2" place="2" resultid="2031" />
                    <RANKING order="3" place="3" resultid="3466" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4486" daytime="19:26" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1322" daytime="19:32" gender="F" number="46" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1323" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3024" />
                    <RANKING order="2" place="-1" resultid="3749" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4487" daytime="19:32" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1324" daytime="19:40" gender="M" number="47" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1325" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2433" />
                    <RANKING order="2" place="2" resultid="3772" />
                    <RANKING order="3" place="3" resultid="3052" />
                    <RANKING order="4" place="4" resultid="1721" />
                    <RANKING order="5" place="5" resultid="3245" />
                    <RANKING order="6" place="6" resultid="3761" />
                    <RANKING order="7" place="-1" resultid="3033" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4488" daytime="19:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1326" daytime="19:46" gender="M" number="48" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1327" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3034" />
                    <RANKING order="2" place="2" resultid="3053" />
                    <RANKING order="3" place="3" resultid="2434" />
                    <RANKING order="4" place="4" resultid="3773" />
                    <RANKING order="5" place="5" resultid="2034" />
                    <RANKING order="6" place="6" resultid="3473" />
                    <RANKING order="7" place="7" resultid="3246" />
                    <RANKING order="8" place="-1" resultid="2177" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4489" daytime="19:46" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1328" daytime="19:54" gender="M" number="49" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1329" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3036" />
                    <RANKING order="2" place="2" resultid="1548" />
                    <RANKING order="3" place="3" resultid="3754" />
                    <RANKING order="4" place="4" resultid="2035" />
                    <RANKING order="5" place="5" resultid="1723" />
                    <RANKING order="6" place="6" resultid="3474" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4490" daytime="19:54" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1330" daytime="20:00" gender="M" number="50" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1331" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3035" />
                    <RANKING order="2" place="2" resultid="2435" />
                    <RANKING order="3" place="3" resultid="1722" />
                    <RANKING order="4" place="-1" resultid="2178" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4491" daytime="20:00" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1332" daytime="20:06" gender="M" number="51" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1333" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3037" />
                    <RANKING order="2" place="2" resultid="1724" />
                    <RANKING order="3" place="3" resultid="3755" />
                    <RANKING order="4" place="4" resultid="2036" />
                    <RANKING order="5" place="5" resultid="2179" />
                    <RANKING order="6" place="6" resultid="3475" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4492" daytime="20:06" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="4970" gender="F" number="68" order="17" round="TIMETRIAL" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4971" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4973" />
                    <RANKING order="2" place="2" resultid="4976" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4972" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-04-14" daytime="08:45" endtime="12:56" number="5" officialmeeting="08:00" warmupfrom="07:30" warmupuntil="08:30">
          <EVENTS>
            <EVENT eventid="1334" daytime="08:46" gender="F" number="52" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1335" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2885" />
                    <RANKING order="2" place="2" resultid="3170" />
                    <RANKING order="3" place="3" resultid="2330" />
                    <RANKING order="4" place="4" resultid="2956" />
                    <RANKING order="5" place="5" resultid="2414" />
                    <RANKING order="6" place="6" resultid="3820" />
                    <RANKING order="7" place="7" resultid="2372" />
                    <RANKING order="8" place="8" resultid="1664" />
                    <RANKING order="9" place="9" resultid="3109" />
                    <RANKING order="10" place="-1" resultid="1787" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1336" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1688" />
                    <RANKING order="2" place="2" resultid="2727" />
                    <RANKING order="3" place="3" resultid="3615" />
                    <RANKING order="4" place="4" resultid="2275" />
                    <RANKING order="5" place="5" resultid="2680" />
                    <RANKING order="6" place="6" resultid="1431" />
                    <RANKING order="7" place="7" resultid="3709" />
                    <RANKING order="8" place="8" resultid="2738" />
                    <RANKING order="9" place="9" resultid="3394" />
                    <RANKING order="10" place="-1" resultid="3293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1337" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3486" />
                    <RANKING order="2" place="2" resultid="3158" />
                    <RANKING order="3" place="3" resultid="1953" />
                    <RANKING order="4" place="4" resultid="3104" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1338" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2458" />
                    <RANKING order="2" place="2" resultid="2318" />
                    <RANKING order="3" place="3" resultid="2047" />
                    <RANKING order="4" place="4" resultid="1750" />
                    <RANKING order="5" place="5" resultid="3415" />
                    <RANKING order="6" place="6" resultid="1994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1339" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2060" />
                    <RANKING order="2" place="2" resultid="1450" />
                    <RANKING order="3" place="3" resultid="2246" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1340" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3503" />
                    <RANKING order="2" place="2" resultid="1474" />
                    <RANKING order="3" place="3" resultid="3316" />
                    <RANKING order="4" place="4" resultid="3372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1341" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3382" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4493" daytime="08:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4494" daytime="08:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4495" daytime="08:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4496" daytime="08:54" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4497" daytime="08:56" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1342" daytime="08:58" gender="M" number="53" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1343" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2306" />
                    <RANKING order="2" place="2" resultid="2762" />
                    <RANKING order="3" place="3" resultid="1652" />
                    <RANKING order="4" place="4" resultid="3633" />
                    <RANKING order="5" place="5" resultid="2342" />
                    <RANKING order="6" place="6" resultid="2798" />
                    <RANKING order="7" place="7" resultid="3687" />
                    <RANKING order="8" place="8" resultid="3597" />
                    <RANKING order="9" place="9" resultid="3188" />
                    <RANKING order="10" place="10" resultid="2785" />
                    <RANKING order="11" place="11" resultid="3651" />
                    <RANKING order="12" place="-1" resultid="2366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1344" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1573" />
                    <RANKING order="2" place="2" resultid="1928" />
                    <RANKING order="3" place="3" resultid="3587" />
                    <RANKING order="4" place="4" resultid="2288" />
                    <RANKING order="5" place="5" resultid="3609" />
                    <RANKING order="6" place="6" resultid="2734" />
                    <RANKING order="7" place="7" resultid="3669" />
                    <RANKING order="8" place="8" resultid="3444" />
                    <RANKING order="9" place="9" resultid="2294" />
                    <RANKING order="10" place="-1" resultid="2018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1345" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1567" />
                    <RANKING order="2" place="2" resultid="2973" />
                    <RANKING order="3" place="3" resultid="3522" />
                    <RANKING order="4" place="4" resultid="1629" />
                    <RANKING order="5" place="5" resultid="2348" />
                    <RANKING order="6" place="6" resultid="1501" />
                    <RANKING order="7" place="7" resultid="1585" />
                    <RANKING order="8" place="8" resultid="1935" />
                    <RANKING order="9" place="9" resultid="3715" />
                    <RANKING order="10" place="10" resultid="2634" />
                    <RANKING order="11" place="11" resultid="3427" />
                    <RANKING order="12" place="-1" resultid="2651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1346" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2493" />
                    <RANKING order="2" place="2" resultid="2585" />
                    <RANKING order="3" place="3" resultid="2390" />
                    <RANKING order="4" place="4" resultid="2944" />
                    <RANKING order="5" place="5" resultid="3510" />
                    <RANKING order="6" place="6" resultid="1579" />
                    <RANKING order="7" place="7" resultid="2000" />
                    <RANKING order="8" place="8" resultid="1990" />
                    <RANKING order="9" place="-1" resultid="3152" />
                    <RANKING order="10" place="-1" resultid="3462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1347" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2512" />
                    <RANKING order="2" place="2" resultid="1409" />
                    <RANKING order="3" place="3" resultid="2558" />
                    <RANKING order="4" place="4" resultid="3272" />
                    <RANKING order="5" place="5" resultid="2109" />
                    <RANKING order="6" place="6" resultid="3433" />
                    <RANKING order="7" place="-1" resultid="3456" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1348" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2750" />
                    <RANKING order="2" place="2" resultid="2085" />
                    <RANKING order="3" place="3" resultid="3016" />
                    <RANKING order="4" place="4" resultid="3627" />
                    <RANKING order="5" place="5" resultid="2234" />
                    <RANKING order="6" place="6" resultid="3333" />
                    <RANKING order="7" place="7" resultid="1608" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1349" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1823" />
                    <RANKING order="2" place="2" resultid="2078" />
                    <RANKING order="3" place="3" resultid="1912" />
                    <RANKING order="4" place="4" resultid="1414" />
                    <RANKING order="5" place="5" resultid="1888" />
                    <RANKING order="6" place="6" resultid="1893" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4498" daytime="08:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4499" daytime="09:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4500" daytime="09:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4501" daytime="09:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4502" daytime="09:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4503" daytime="09:12" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4504" daytime="09:14" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4505" daytime="09:16" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1350" daytime="09:18" gender="F" number="54" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1351" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2886" />
                    <RANKING order="2" place="2" resultid="2828" />
                    <RANKING order="3" place="3" resultid="2780" />
                    <RANKING order="4" place="4" resultid="2336" />
                    <RANKING order="5" place="5" resultid="2402" />
                    <RANKING order="6" place="6" resultid="2950" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1352" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2681" />
                    <RANKING order="2" place="2" resultid="2728" />
                    <RANKING order="3" place="3" resultid="2693" />
                    <RANKING order="4" place="4" resultid="2687" />
                    <RANKING order="5" place="5" resultid="2139" />
                    <RANKING order="6" place="6" resultid="2717" />
                    <RANKING order="7" place="7" resultid="2378" />
                    <RANKING order="8" place="8" resultid="2739" />
                    <RANKING order="9" place="9" resultid="1818" />
                    <RANKING order="10" place="10" resultid="2844" />
                    <RANKING order="11" place="11" resultid="3140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1353" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2525" />
                    <RANKING order="2" place="2" resultid="2453" />
                    <RANKING order="3" place="3" resultid="2630" />
                    <RANKING order="4" place="4" resultid="2115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1354" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3357" />
                    <RANKING order="2" place="2" resultid="1835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1355" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2546" />
                    <RANKING order="2" place="2" resultid="2061" />
                    <RANKING order="3" place="3" resultid="1426" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1356" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2890" />
                    <RANKING order="2" place="2" resultid="3504" />
                    <RANKING order="3" place="3" resultid="3311" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1357" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2939" />
                    <RANKING order="2" place="2" resultid="3005" />
                    <RANKING order="3" place="3" resultid="3351" />
                    <RANKING order="4" place="-1" resultid="2977" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4506" daytime="09:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4507" daytime="09:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4508" daytime="09:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4509" daytime="09:38" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4510" daytime="09:44" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1358" daytime="09:52" gender="M" number="55" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1359" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2862" />
                    <RANKING order="2" place="2" resultid="2324" />
                    <RANKING order="3" place="3" resultid="2756" />
                    <RANKING order="4" place="4" resultid="2761" />
                    <RANKING order="5" place="5" resultid="2768" />
                    <RANKING order="6" place="6" resultid="2774" />
                    <RANKING order="7" place="7" resultid="2833" />
                    <RANKING order="8" place="8" resultid="2797" />
                    <RANKING order="9" place="9" resultid="2208" />
                    <RANKING order="10" place="10" resultid="2821" />
                    <RANKING order="11" place="11" resultid="3603" />
                    <RANKING order="12" place="12" resultid="2901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1360" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2850" />
                    <RANKING order="2" place="2" resultid="2711" />
                    <RANKING order="3" place="3" resultid="2745" />
                    <RANKING order="4" place="4" resultid="2668" />
                    <RANKING order="5" place="5" resultid="3164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1361" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2264" />
                    <RANKING order="2" place="2" resultid="2541" />
                    <RANKING order="3" place="3" resultid="3278" />
                    <RANKING order="4" place="4" resultid="2488" />
                    <RANKING order="5" place="5" resultid="1507" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1362" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2252" />
                    <RANKING order="2" place="2" resultid="2856" />
                    <RANKING order="3" place="3" resultid="2103" />
                    <RANKING order="4" place="4" resultid="3540" />
                    <RANKING order="5" place="5" resultid="2595" />
                    <RANKING order="6" place="6" resultid="2360" />
                    <RANKING order="7" place="7" resultid="1591" />
                    <RANKING order="8" place="8" resultid="2127" />
                    <RANKING order="9" place="9" resultid="3322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1363" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3498" />
                    <RANKING order="2" place="2" resultid="3409" />
                    <RANKING order="3" place="3" resultid="3733" />
                    <RANKING order="4" place="4" resultid="3363" />
                    <RANKING order="5" place="-1" resultid="2552" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1364" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2506" />
                    <RANKING order="2" place="2" resultid="2986" />
                    <RANKING order="3" place="3" resultid="3260" />
                    <RANKING order="4" place="4" resultid="1898" />
                    <RANKING order="5" place="5" resultid="2569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1365" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3339" />
                    <RANKING order="2" place="2" resultid="1903" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4511" daytime="09:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4512" daytime="09:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4513" daytime="10:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4514" daytime="10:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4515" daytime="10:16" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4516" daytime="10:22" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1366" daytime="10:28" gender="F" number="56" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1367" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2810" />
                    <RANKING order="2" place="2" resultid="2874" />
                    <RANKING order="3" place="3" resultid="2401" />
                    <RANKING order="4" place="4" resultid="1700" />
                    <RANKING order="5" place="5" resultid="2949" />
                    <RANKING order="6" place="6" resultid="3212" />
                    <RANKING order="7" place="7" resultid="2006" />
                    <RANKING order="8" place="8" resultid="3305" />
                    <RANKING order="9" place="9" resultid="1670" />
                    <RANKING order="10" place="-1" resultid="1444" />
                    <RANKING order="11" place="-1" resultid="1542" />
                    <RANKING order="12" place="-1" resultid="1811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1368" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2276" />
                    <RANKING order="2" place="2" resultid="3811" />
                    <RANKING order="3" place="3" resultid="2686" />
                    <RANKING order="4" place="4" resultid="1432" />
                    <RANKING order="5" place="5" resultid="2675" />
                    <RANKING order="6" place="6" resultid="1682" />
                    <RANKING order="7" place="7" resultid="1771" />
                    <RANKING order="8" place="8" resultid="2692" />
                    <RANKING order="9" place="9" resultid="2997" />
                    <RANKING order="10" place="10" resultid="2151" />
                    <RANKING order="11" place="11" resultid="3328" />
                    <RANKING order="12" place="12" resultid="3727" />
                    <RANKING order="13" place="13" resultid="3721" />
                    <RANKING order="14" place="14" resultid="2420" />
                    <RANKING order="15" place="15" resultid="3663" />
                    <RANKING order="16" place="16" resultid="1519" />
                    <RANKING order="17" place="17" resultid="3242" />
                    <RANKING order="18" place="18" resultid="3388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1369" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1873" />
                    <RANKING order="2" place="2" resultid="1480" />
                    <RANKING order="3" place="3" resultid="3546" />
                    <RANKING order="4" place="4" resultid="1613" />
                    <RANKING order="5" place="5" resultid="2282" />
                    <RANKING order="6" place="6" resultid="1496" />
                    <RANKING order="7" place="7" resultid="2114" />
                    <RANKING order="8" place="8" resultid="3569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1370" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2968" />
                    <RANKING order="2" place="2" resultid="2459" />
                    <RANKING order="3" place="3" resultid="2048" />
                    <RANKING order="4" place="4" resultid="3266" />
                    <RANKING order="5" place="5" resultid="3356" />
                    <RANKING order="6" place="6" resultid="1420" />
                    <RANKING order="7" place="7" resultid="1635" />
                    <RANKING order="8" place="8" resultid="3400" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1371" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3492" />
                    <RANKING order="2" place="2" resultid="1490" />
                    <RANKING order="3" place="3" resultid="3218" />
                    <RANKING order="4" place="4" resultid="1976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1372" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1739" />
                    <RANKING order="2" place="2" resultid="2052" />
                    <RANKING order="3" place="3" resultid="3799" />
                    <RANKING order="4" place="4" resultid="3310" />
                    <RANKING order="5" place="-1" resultid="2073" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1373" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2258" />
                    <RANKING order="2" place="2" resultid="3793" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4517" daytime="10:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4518" daytime="10:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4519" daytime="10:36" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4520" daytime="10:38" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4521" daytime="10:42" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4522" daytime="10:44" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4523" daytime="10:48" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4524" daytime="10:50" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1374" daytime="10:54" gender="M" number="57" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1375" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2312" />
                    <RANKING order="2" place="2" resultid="1797" />
                    <RANKING order="3" place="3" resultid="3581" />
                    <RANKING order="4" place="4" resultid="3128" />
                    <RANKING order="5" place="5" resultid="2396" />
                    <RANKING order="6" place="6" resultid="3176" />
                    <RANKING order="7" place="7" resultid="2175" />
                    <RANKING order="8" place="8" resultid="2822" />
                    <RANKING order="9" place="9" resultid="1857" />
                    <RANKING order="10" place="10" resultid="3230" />
                    <RANKING order="11" place="11" resultid="1863" />
                    <RANKING order="12" place="12" resultid="2786" />
                    <RANKING order="13" place="13" resultid="1694" />
                    <RANKING order="14" place="14" resultid="2169" />
                    <RANKING order="15" place="-1" resultid="3194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1376" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2145" />
                    <RANKING order="2" place="2" resultid="2933" />
                    <RANKING order="3" place="3" resultid="2705" />
                    <RANKING order="4" place="4" resultid="1929" />
                    <RANKING order="5" place="5" resultid="2699" />
                    <RANKING order="6" place="6" resultid="2669" />
                    <RANKING order="7" place="7" resultid="1646" />
                    <RANKING order="8" place="8" resultid="2384" />
                    <RANKING order="9" place="9" resultid="1718" />
                    <RANKING order="10" place="10" resultid="3681" />
                    <RANKING order="11" place="11" resultid="2030" />
                    <RANKING order="12" place="-1" resultid="3224" />
                    <RANKING order="13" place="-1" resultid="1959" />
                    <RANKING order="14" place="-1" resultid="2157" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1377" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1878" />
                    <RANKING order="2" place="2" resultid="1458" />
                    <RANKING order="3" place="3" resultid="3299" />
                    <RANKING order="4" place="4" resultid="2640" />
                    <RANKING order="5" place="5" resultid="3528" />
                    <RANKING order="6" place="6" resultid="1941" />
                    <RANKING order="7" place="7" resultid="3182" />
                    <RANKING order="8" place="8" resultid="1982" />
                    <RANKING order="9" place="9" resultid="2121" />
                    <RANKING order="10" place="10" resultid="2604" />
                    <RANKING order="11" place="-1" resultid="3010" />
                    <RANKING order="12" place="-1" resultid="2012" />
                    <RANKING order="13" place="-1" resultid="3069" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1378" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2477" />
                    <RANKING order="2" place="2" resultid="2646" />
                    <RANKING order="3" place="3" resultid="2483" />
                    <RANKING order="4" place="4" resultid="1624" />
                    <RANKING order="5" place="5" resultid="2599" />
                    <RANKING order="6" place="6" resultid="3787" />
                    <RANKING order="7" place="7" resultid="2580" />
                    <RANKING order="8" place="8" resultid="2574" />
                    <RANKING order="9" place="9" resultid="1765" />
                    <RANKING order="10" place="10" resultid="2067" />
                    <RANKING order="11" place="11" resultid="2133" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1379" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2991" />
                    <RANKING order="2" place="2" resultid="3742" />
                    <RANKING order="3" place="3" resultid="3200" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1380" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2467" />
                    <RANKING order="2" place="2" resultid="3563" />
                    <RANKING order="3" place="3" resultid="2097" />
                    <RANKING order="4" place="4" resultid="1513" />
                    <RANKING order="5" place="5" resultid="2354" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1381" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2838" />
                    <RANKING order="2" place="2" resultid="1824" />
                    <RANKING order="3" place="3" resultid="2927" />
                    <RANKING order="4" place="4" resultid="2079" />
                    <RANKING order="5" place="5" resultid="2424" />
                    <RANKING order="6" place="6" resultid="2091" />
                    <RANKING order="7" place="7" resultid="3134" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4525" daytime="10:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4526" daytime="10:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4527" daytime="11:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4528" daytime="11:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4529" daytime="11:06" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4530" daytime="11:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4531" daytime="11:12" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="4532" daytime="11:16" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="4533" daytime="11:18" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1382" daytime="11:20" gender="F" number="58" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1383" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3029" />
                    <RANKING order="2" place="2" resultid="3051" />
                    <RANKING order="3" place="3" resultid="2430" />
                    <RANKING order="4" place="4" resultid="1720" />
                    <RANKING order="5" place="5" resultid="3770" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4534" daytime="11:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1384" daytime="11:28" gender="F" number="59" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1385" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3027" />
                    <RANKING order="2" place="2" resultid="3769" />
                    <RANKING order="3" place="3" resultid="3050" />
                    <RANKING order="4" place="4" resultid="2429" />
                    <RANKING order="5" place="5" resultid="3828" />
                    <RANKING order="6" place="6" resultid="3243" />
                    <RANKING order="7" place="7" resultid="3469" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4535" daytime="11:28" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1386" daytime="11:34" gender="F" number="60" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1387" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3028" />
                    <RANKING order="2" place="2" resultid="3751" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4536" daytime="11:34" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1388" daytime="11:40" gender="F" number="61" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1389" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3025" />
                    <RANKING order="2" place="2" resultid="3467" />
                    <RANKING order="3" place="-1" resultid="2032" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4537" daytime="11:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1390" daytime="11:46" gender="F" number="62" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1391" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3750" />
                    <RANKING order="2" place="2" resultid="3468" />
                    <RANKING order="3" place="-1" resultid="3026" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4538" daytime="11:46" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1392" daytime="11:52" gender="M" number="63" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1393" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3038" />
                    <RANKING order="2" place="2" resultid="2436" />
                    <RANKING order="3" place="3" resultid="3774" />
                    <RANKING order="4" place="4" resultid="3054" />
                    <RANKING order="5" place="5" resultid="1725" />
                    <RANKING order="6" place="6" resultid="3247" />
                    <RANKING order="7" place="7" resultid="3762" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4539" daytime="11:52" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1394" daytime="11:58" gender="M" number="64" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1395" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3039" />
                    <RANKING order="2" place="2" resultid="3055" />
                    <RANKING order="3" place="3" resultid="3775" />
                    <RANKING order="4" place="4" resultid="2437" />
                    <RANKING order="5" place="5" resultid="2037" />
                    <RANKING order="6" place="-1" resultid="2180" />
                    <RANKING order="7" place="-1" resultid="3248" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4540" daytime="11:58" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1396" daytime="12:04" gender="M" number="65" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1397" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3041" />
                    <RANKING order="2" place="2" resultid="1549" />
                    <RANKING order="3" place="3" resultid="2039" />
                    <RANKING order="4" place="4" resultid="3757" />
                    <RANKING order="5" place="5" resultid="1727" />
                    <RANKING order="6" place="6" resultid="3477" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4541" daytime="12:04" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1398" daytime="12:10" gender="M" number="66" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1399" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3042" />
                    <RANKING order="2" place="2" resultid="2439" />
                    <RANKING order="3" place="3" resultid="2182" />
                    <RANKING order="4" place="4" resultid="1728" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4542" daytime="12:10" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1400" daytime="12:16" gender="M" number="67" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1401" agemax="-1" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3040" />
                    <RANKING order="2" place="2" resultid="3756" />
                    <RANKING order="3" place="3" resultid="1726" />
                    <RANKING order="4" place="4" resultid="3476" />
                    <RANKING order="5" place="5" resultid="2181" />
                    <RANKING order="6" place="6" resultid="2038" />
                    <RANKING order="7" place="7" resultid="2438" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4543" daytime="12:16" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="13038" nation="BRA" region="PR" clubid="1733" swrid="93759" name="Associação De Pais E Atletas De Natação Ws/Crb" shortname="Apan/Ws">
          <ATHLETES>
            <ATHLETE firstname="Heloisa" lastname="Daniele Silva" birthdate="2010-07-06" gender="F" nation="BRA" license="359593" swrid="5588628" athleteid="1766" externalid="359593">
              <RESULTS>
                <RESULT eventid="1064" points="354" swimtime="00:02:54.01" resultid="1767" heatid="4269" lane="3" entrytime="00:02:54.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="461" swimtime="00:01:06.91" resultid="1768" heatid="4326" lane="1" entrytime="00:01:09.94" entrycourse="LCM" />
                <RESULT eventid="1228" points="485" swimtime="00:00:30.03" resultid="1769" heatid="4403" lane="8" entrytime="00:00:30.78" entrycourse="LCM" />
                <RESULT eventid="1298" points="450" swimtime="00:00:35.05" resultid="1770" heatid="4474" lane="7" entrytime="00:00:37.29" entrycourse="LCM" />
                <RESULT eventid="1366" points="382" swimtime="00:01:18.97" resultid="1771" heatid="4523" lane="7" entrytime="00:01:17.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Zanatta Flizikowski" birthdate="2007-09-14" gender="F" nation="BRA" license="366835" swrid="5600281" athleteid="1756" externalid="366835">
              <RESULTS>
                <RESULT eventid="1180" points="247" swimtime="00:00:46.46" resultid="1757" heatid="4357" lane="8" entrytime="00:00:45.88" entrycourse="LCM" />
                <RESULT eventid="1228" points="261" swimtime="00:00:36.92" resultid="1758" heatid="4399" lane="8" entrytime="00:00:35.84" entrycourse="LCM" />
                <RESULT eventid="1212" points="244" swimtime="00:01:42.54" resultid="1759" heatid="4380" lane="6" entrytime="00:01:38.53" entrycourse="LCM" />
                <RESULT eventid="1282" points="236" swimtime="00:03:02.41" resultid="1760" heatid="4452" lane="8" entrytime="00:02:50.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabelly" lastname="Mendonca Bello" birthdate="2008-04-15" gender="F" nation="BRA" license="376996" swrid="5600217" athleteid="1751" externalid="376996">
              <RESULTS>
                <RESULT eventid="1080" points="353" swimtime="00:03:14.61" resultid="1752" heatid="4280" lane="2" entrytime="00:03:11.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="410" swimtime="00:00:39.25" resultid="1753" heatid="4357" lane="3" entrytime="00:00:41.92" entrycourse="LCM" />
                <RESULT eventid="1228" points="431" swimtime="00:00:31.24" resultid="1754" heatid="4402" lane="5" entrytime="00:00:31.05" entrycourse="LCM" />
                <RESULT eventid="1212" points="363" swimtime="00:01:29.83" resultid="1755" heatid="4382" lane="1" entrytime="00:01:29.32" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Arceli Silva" birthdate="2008-03-04" gender="M" nation="BRA" license="331565" swrid="5385686" athleteid="1761" externalid="331565">
              <RESULTS>
                <RESULT eventid="1104" points="395" swimtime="00:00:30.33" resultid="1762" heatid="4300" lane="3" entrytime="00:00:30.60" entrycourse="LCM" />
                <RESULT eventid="1156" points="423" swimtime="00:01:02.42" resultid="1763" heatid="4340" lane="7" entrytime="00:01:06.29" entrycourse="LCM" />
                <RESULT eventid="1236" points="369" swimtime="00:00:29.15" resultid="1764" heatid="4415" lane="1" entrytime="00:00:29.68" entrycourse="LCM" />
                <RESULT eventid="1374" points="399" swimtime="00:01:10.06" resultid="1765" heatid="4530" lane="3" entrytime="00:01:09.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Sieck" birthdate="2011-01-20" gender="F" nation="BRA" license="382234" swrid="5602584" athleteid="1782" externalid="382234">
              <RESULTS>
                <RESULT eventid="1096" points="164" swimtime="00:00:44.60" resultid="1783" heatid="4291" lane="4" entrytime="00:00:50.12" entrycourse="LCM" />
                <RESULT eventid="1164" points="110" swimtime="00:04:14.21" resultid="1784" heatid="4349" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:56.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="198" swimtime="00:01:28.61" resultid="1785" heatid="4320" lane="4" entrytime="00:01:28.51" entrycourse="LCM" />
                <RESULT eventid="1228" points="214" swimtime="00:00:39.42" resultid="1786" heatid="4398" lane="8" entrytime="00:00:40.14" entrycourse="LCM" />
                <RESULT eventid="1334" status="DSQ" swimtime="00:01:55.16" resultid="1787" heatid="4494" lane="5" entrytime="00:01:45.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Alexandre Azevedo" birthdate="2008-05-20" gender="M" nation="BRA" license="398694" swrid="5717240" athleteid="1772" externalid="398694">
              <RESULTS>
                <RESULT eventid="1156" points="280" swimtime="00:01:11.58" resultid="1773" heatid="4336" lane="4" entrytime="00:01:11.37" entrycourse="LCM" />
                <RESULT eventid="1188" points="231" swimtime="00:00:42.28" resultid="1774" heatid="4361" lane="4" />
                <RESULT eventid="1220" points="203" swimtime="00:01:36.66" resultid="1775" heatid="4387" lane="5" entrytime="00:01:40.53" entrycourse="LCM" />
                <RESULT eventid="1236" points="296" swimtime="00:00:31.35" resultid="1776" heatid="4409" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Reis" birthdate="2008-04-07" gender="F" nation="BRA" license="378820" swrid="5600243" athleteid="1777" externalid="378820">
              <RESULTS>
                <RESULT eventid="1096" points="178" swimtime="00:00:43.38" resultid="1778" heatid="4290" lane="4" />
                <RESULT eventid="1148" points="227" swimtime="00:01:24.70" resultid="1779" heatid="4322" lane="8" entrytime="00:01:22.05" entrycourse="LCM" />
                <RESULT eventid="1228" points="223" swimtime="00:00:38.89" resultid="1780" heatid="4398" lane="5" entrytime="00:00:36.71" entrycourse="LCM" />
                <RESULT eventid="1298" points="222" swimtime="00:00:44.31" resultid="1781" heatid="4472" lane="2" entrytime="00:00:43.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Cravcenco Marcondes" birthdate="2011-05-06" gender="M" nation="BRA" license="406867" swrid="5723023" athleteid="1802" externalid="406867">
              <RESULTS>
                <RESULT eventid="1156" points="192" swimtime="00:01:21.17" resultid="1803" heatid="4334" lane="3" entrytime="00:01:23.37" entrycourse="LCM" />
                <RESULT eventid="1188" points="147" swimtime="00:00:49.09" resultid="1804" heatid="4361" lane="7" />
                <RESULT eventid="1236" points="242" swimtime="00:00:33.54" resultid="1805" heatid="4408" lane="2" />
                <RESULT eventid="1306" points="170" swimtime="00:00:42.45" resultid="1806" heatid="4477" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Zeclhynski Silva" birthdate="2006-09-14" gender="F" nation="BRA" license="330727" swrid="5600283" athleteid="1734" externalid="330727">
              <RESULTS>
                <RESULT eventid="1064" points="505" swimtime="00:02:34.57" resultid="1735" heatid="4271" lane="6" entrytime="00:02:32.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="629" swimtime="00:01:00.34" resultid="1736" heatid="4330" lane="6" entrytime="00:01:01.02" entrycourse="LCM" />
                <RESULT eventid="1228" points="600" swimtime="00:00:27.99" resultid="1737" heatid="4405" lane="3" entrytime="00:00:27.83" entrycourse="LCM" />
                <RESULT eventid="1298" points="695" swimtime="00:00:30.32" resultid="1738" heatid="4475" lane="4" entrytime="00:00:30.32" entrycourse="LCM" />
                <RESULT eventid="1366" points="620" swimtime="00:01:07.23" resultid="1739" heatid="4524" lane="4" entrytime="00:01:06.10" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Rosa Silva" birthdate="2011-03-25" gender="F" nation="BRA" license="392120" swrid="5602579" athleteid="1788" externalid="392120">
              <RESULTS>
                <RESULT eventid="1148" points="240" swimtime="00:01:23.16" resultid="1789" heatid="4319" lane="5" />
                <RESULT eventid="1180" points="178" swimtime="00:00:51.77" resultid="1790" heatid="4356" lane="1" />
                <RESULT eventid="1228" points="236" swimtime="00:00:38.18" resultid="1791" heatid="4398" lane="1" entrytime="00:00:39.90" entrycourse="LCM" />
                <RESULT eventid="1212" points="176" swimtime="00:01:54.30" resultid="1792" heatid="4379" lane="2" entrytime="00:01:52.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="De Reginalda" birthdate="2011-07-22" gender="M" nation="BRA" license="400323" swrid="5717257" athleteid="1793" externalid="400323">
              <RESULTS>
                <RESULT eventid="1156" points="391" swimtime="00:01:04.08" resultid="1794" heatid="4339" lane="1" entrytime="00:01:07.31" entrycourse="LCM" />
                <RESULT eventid="1236" points="405" swimtime="00:00:28.25" resultid="1795" heatid="4408" lane="3" />
                <RESULT eventid="1306" points="364" swimtime="00:00:32.96" resultid="1796" heatid="4477" lane="4" />
                <RESULT eventid="1374" points="334" swimtime="00:01:14.30" resultid="1797" heatid="4528" lane="2" entrytime="00:01:17.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonia" lastname="Adam  Fracaro" birthdate="2010-04-27" gender="F" nation="BRA" license="382212" swrid="5588512" athleteid="1740" externalid="382212">
              <RESULTS>
                <RESULT eventid="1148" points="339" swimtime="00:01:14.16" resultid="1741" heatid="4324" lane="8" entrytime="00:01:13.40" entrycourse="LCM" />
                <RESULT eventid="1180" points="152" swimtime="00:00:54.53" resultid="1742" heatid="4355" lane="3" />
                <RESULT eventid="1212" status="DSQ" swimtime="00:02:00.49" resultid="1743" heatid="4378" lane="5" />
                <RESULT eventid="1282" points="303" swimtime="00:02:47.93" resultid="1744" heatid="4452" lane="7" entrytime="00:02:47.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Zanchetta Silva" birthdate="2010-08-05" gender="F" nation="BRA" license="406865" swrid="5717308" athleteid="1798" externalid="406865">
              <RESULTS>
                <RESULT eventid="1148" points="190" swimtime="00:01:29.89" resultid="1799" heatid="4320" lane="5" entrytime="00:01:36.50" entrycourse="LCM" />
                <RESULT eventid="1228" points="211" swimtime="00:00:39.64" resultid="1800" heatid="4396" lane="7" />
                <RESULT eventid="1298" points="195" swimtime="00:00:46.25" resultid="1801" heatid="4470" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Da Costa Riekes" birthdate="2008-06-19" gender="F" nation="BRA" license="331686" swrid="5600143" athleteid="1745" externalid="331686">
              <RESULTS>
                <RESULT eventid="1096" points="471" swimtime="00:00:31.38" resultid="1746" heatid="4294" lane="7" entrytime="00:00:32.02" entrycourse="LCM" />
                <RESULT eventid="1148" points="534" swimtime="00:01:03.73" resultid="1747" heatid="4329" lane="4" entrytime="00:01:04.00" entrycourse="LCM" />
                <RESULT eventid="1228" points="524" swimtime="00:00:29.28" resultid="1748" heatid="4404" lane="2" entrytime="00:00:29.74" entrycourse="LCM" />
                <RESULT eventid="1282" points="500" swimtime="00:02:22.15" resultid="1749" heatid="4456" lane="7" entrytime="00:02:24.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="432" swimtime="00:01:13.39" resultid="1750" heatid="4497" lane="8" entrytime="00:01:13.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marjori" lastname="Leticia Oliveira" birthdate="2011-05-23" gender="F" nation="BRA" license="406869" swrid="5717279" athleteid="1807" externalid="406869">
              <RESULTS>
                <RESULT eventid="1148" points="252" swimtime="00:01:21.78" resultid="1808" heatid="4321" lane="1" entrytime="00:01:26.97" entrycourse="LCM" />
                <RESULT eventid="1228" points="299" swimtime="00:00:35.29" resultid="1809" heatid="4397" lane="7" />
                <RESULT eventid="1298" points="218" swimtime="00:00:44.57" resultid="1810" heatid="4471" lane="6" />
                <RESULT eventid="1366" status="DNS" swimtime="00:00:00.00" resultid="1811" heatid="4518" lane="7" entrytime="00:01:42.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2416" nation="BRA" region="PR" clubid="1552" swrid="93758" name="Apan/Maringá">
          <ATHLETES>
            <ATHLETE firstname="Daniela" lastname="Inoue" birthdate="2008-10-31" gender="F" nation="BRA" license="378348" swrid="5603856" athleteid="1630" externalid="378348">
              <RESULTS>
                <RESULT eventid="1096" points="318" swimtime="00:00:35.76" resultid="1631" heatid="4292" lane="4" entrytime="00:00:37.06" entrycourse="LCM" />
                <RESULT eventid="1148" points="389" swimtime="00:01:10.78" resultid="1632" heatid="4324" lane="2" entrytime="00:01:12.28" entrycourse="LCM" />
                <RESULT eventid="1228" points="414" swimtime="00:00:31.67" resultid="1633" heatid="4401" lane="7" entrytime="00:00:32.51" entrycourse="LCM" />
                <RESULT eventid="1298" points="354" swimtime="00:00:37.96" resultid="1634" heatid="4473" lane="1" entrytime="00:00:41.25" entrycourse="LCM" />
                <RESULT eventid="1366" points="313" swimtime="00:01:24.40" resultid="1635" heatid="4519" lane="6" entrytime="00:01:29.94" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietro" lastname="Nabas De Assis" birthdate="2011-07-09" gender="M" nation="BRA" license="366968" swrid="5603878" athleteid="1653" externalid="366968">
              <RESULTS>
                <RESULT eventid="1088" points="338" swimtime="00:03:00.13" resultid="1654" heatid="4284" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="367" swimtime="00:00:36.22" resultid="1655" heatid="4365" lane="4" entrytime="00:00:37.50" entrycourse="LCM" />
                <RESULT eventid="1220" points="331" swimtime="00:01:22.16" resultid="1656" heatid="4391" lane="2" entrytime="00:01:22.78" entrycourse="LCM" />
                <RESULT eventid="1236" points="291" swimtime="00:00:31.54" resultid="1657" heatid="4411" lane="5" entrytime="00:00:33.56" entrycourse="LCM" />
                <RESULT eventid="1274" points="262" swimtime="00:02:58.15" resultid="1658" heatid="4440" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Sossai Altoe" birthdate="2006-09-04" gender="M" nation="BRA" license="296488" swrid="5603915" athleteid="1553" externalid="296488">
              <RESULTS>
                <RESULT eventid="1104" points="580" swimtime="00:00:26.69" resultid="1554" heatid="4304" lane="8" entrytime="00:00:27.28" entrycourse="LCM" />
                <RESULT eventid="1156" points="716" swimtime="00:00:52.37" resultid="1555" heatid="4348" lane="6" entrytime="00:00:52.41" entrycourse="LCM" />
                <RESULT eventid="1236" points="585" swimtime="00:00:24.99" resultid="1556" heatid="4421" lane="1" entrytime="00:00:25.03" entrycourse="LCM" />
                <RESULT eventid="1290" points="635" swimtime="00:01:58.66" resultid="1557" heatid="4469" lane="8" entrytime="00:02:01.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felype" lastname="Gongora Zago" birthdate="2011-09-14" gender="M" nation="BRA" license="392099" swrid="5603848" athleteid="1689" externalid="392099">
              <RESULTS>
                <RESULT eventid="1104" status="DSQ" swimtime="00:00:42.00" resultid="1690" heatid="4297" lane="4" entrytime="00:00:51.80" entrycourse="LCM" />
                <RESULT eventid="1156" points="222" swimtime="00:01:17.30" resultid="1691" heatid="4334" lane="2" entrytime="00:01:27.75" entrycourse="LCM" />
                <RESULT eventid="1236" points="218" swimtime="00:00:34.71" resultid="1692" heatid="4410" lane="5" entrytime="00:00:37.78" entrycourse="LCM" />
                <RESULT eventid="1306" points="146" swimtime="00:00:44.70" resultid="1693" heatid="4478" lane="6" entrytime="00:00:47.68" entrycourse="LCM" />
                <RESULT eventid="1374" points="156" swimtime="00:01:35.80" resultid="1694" heatid="4526" lane="2" entrytime="00:01:47.57" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Biason Santana" birthdate="2009-01-21" gender="M" nation="BRA" license="366969" swrid="5317765" athleteid="1625" externalid="366969">
              <RESULTS>
                <RESULT eventid="1104" points="466" swimtime="00:00:28.72" resultid="1626" heatid="4301" lane="5" entrytime="00:00:29.53" entrycourse="LCM" />
                <RESULT eventid="1172" points="326" swimtime="00:02:40.19" resultid="1627" heatid="4351" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="415" swimtime="00:00:28.03" resultid="1628" heatid="4416" lane="5" entrytime="00:00:27.68" entrycourse="LCM" />
                <RESULT eventid="1342" points="417" swimtime="00:01:06.14" resultid="1629" heatid="4503" lane="8" entrytime="00:01:04.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wellington" lastname="De Lima" birthdate="2008-03-01" gender="M" nation="BRA" license="370024" swrid="5470912" athleteid="1574" externalid="370024">
              <RESULTS>
                <RESULT eventid="1104" points="460" swimtime="00:00:28.83" resultid="1575" heatid="4301" lane="2" entrytime="00:00:30.03" entrycourse="LCM" />
                <RESULT eventid="1156" points="542" swimtime="00:00:57.45" resultid="1576" heatid="4345" lane="4" entrytime="00:00:58.49" entrycourse="LCM" />
                <RESULT eventid="1236" points="502" swimtime="00:00:26.30" resultid="1577" heatid="4418" lane="5" entrytime="00:00:26.85" entrycourse="LCM" />
                <RESULT eventid="1306" points="389" swimtime="00:00:32.24" resultid="1578" heatid="4480" lane="7" entrytime="00:00:33.17" entrycourse="LCM" />
                <RESULT eventid="1342" points="385" swimtime="00:01:07.95" resultid="1579" heatid="4502" lane="7" entrytime="00:01:09.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Furuchi Martins" birthdate="2011-10-05" gender="F" nation="BRA" license="367001" swrid="5602616" athleteid="1707" externalid="367001">
              <RESULTS>
                <RESULT eventid="1080" points="281" swimtime="00:03:29.89" resultid="1708" heatid="4278" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="181" swimtime="00:00:43.18" resultid="1709" heatid="4290" lane="6" />
                <RESULT eventid="1180" points="294" swimtime="00:00:43.83" resultid="1710" heatid="4356" lane="5" entrytime="00:00:49.50" entrycourse="LCM" />
                <RESULT eventid="1212" points="285" swimtime="00:01:37.40" resultid="1711" heatid="4379" lane="3" entrytime="00:01:51.04" entrycourse="LCM" />
                <RESULT eventid="1266" status="DSQ" swimtime="00:03:22.16" resultid="1712" heatid="4434" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Garcia Cavalcante" birthdate="2011-11-21" gender="M" nation="BRA" license="378200" swrid="5603840" athleteid="1592" externalid="378200">
              <RESULTS>
                <RESULT eventid="1088" points="270" swimtime="00:03:13.97" resultid="1593" heatid="4283" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="200" swimtime="00:00:38.02" resultid="1594" heatid="4297" lane="8" />
                <RESULT eventid="1188" points="261" swimtime="00:00:40.56" resultid="1595" heatid="4364" lane="4" entrytime="00:00:42.18" entrycourse="LCM" />
                <RESULT eventid="1220" points="265" swimtime="00:01:28.52" resultid="1596" heatid="4388" lane="4" entrytime="00:01:33.46" entrycourse="LCM" />
                <RESULT eventid="1274" points="233" swimtime="00:03:05.19" resultid="1597" heatid="4443" lane="8" entrytime="00:03:14.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Sol Reolon Gomes" birthdate="2011-02-28" gender="F" nation="BRA" license="392100" swrid="5603914" athleteid="1695" externalid="392100">
              <RESULTS>
                <RESULT eventid="1096" points="319" swimtime="00:00:35.74" resultid="1696" heatid="4290" lane="5" />
                <RESULT eventid="1148" points="420" swimtime="00:01:09.01" resultid="1697" heatid="4323" lane="8" entrytime="00:01:14.75" entrycourse="LCM" />
                <RESULT eventid="1228" points="430" swimtime="00:00:31.28" resultid="1698" heatid="4400" lane="7" entrytime="00:00:33.10" entrycourse="LCM" />
                <RESULT eventid="1298" points="386" swimtime="00:00:36.89" resultid="1699" heatid="4473" lane="6" entrytime="00:00:38.23" entrycourse="LCM" />
                <RESULT eventid="1366" points="319" swimtime="00:01:23.87" resultid="1700" heatid="4519" lane="1" entrytime="00:01:32.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Gabriel Oliveira" birthdate="2006-05-31" gender="M" nation="BRA" license="345589" swrid="5603838" athleteid="1636" externalid="345589">
              <RESULTS>
                <RESULT eventid="1104" points="399" swimtime="00:00:30.25" resultid="1637" heatid="4300" lane="6" entrytime="00:00:31.15" entrycourse="LCM" />
                <RESULT eventid="1156" points="492" swimtime="00:00:59.34" resultid="1638" heatid="4345" lane="8" entrytime="00:00:59.56" entrycourse="LCM" />
                <RESULT eventid="1236" points="458" swimtime="00:00:27.12" resultid="1639" heatid="4417" lane="4" entrytime="00:00:27.25" entrycourse="LCM" />
                <RESULT eventid="1290" points="431" swimtime="00:02:14.97" resultid="1640" heatid="4464" lane="6" entrytime="00:02:21.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Corsine Ferreira" birthdate="2010-03-10" gender="F" nation="BRA" license="353591" swrid="5588608" athleteid="1677" externalid="353591">
              <RESULTS>
                <RESULT eventid="1064" points="386" swimtime="00:02:49.08" resultid="1678" heatid="4270" lane="3" entrytime="00:02:46.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="381" swimtime="00:00:40.21" resultid="1679" heatid="4355" lane="8" />
                <RESULT eventid="1228" points="403" swimtime="00:00:31.94" resultid="1680" heatid="4402" lane="2" entrytime="00:00:31.19" entrycourse="LCM" />
                <RESULT eventid="1298" points="420" swimtime="00:00:35.86" resultid="1681" heatid="4475" lane="1" entrytime="00:00:35.38" entrycourse="LCM" />
                <RESULT eventid="1366" points="391" swimtime="00:01:18.38" resultid="1682" heatid="4523" lane="6" entrytime="00:01:16.89" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Schuch Pimpao" birthdate="2010-12-31" gender="M" nation="BRA" license="355586" swrid="5588908" athleteid="1641" externalid="355586">
              <RESULTS>
                <RESULT eventid="1072" points="324" swimtime="00:02:42.94" resultid="1642" heatid="4274" lane="3" entrytime="00:02:43.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="298" swimtime="00:00:38.81" resultid="1643" heatid="4362" lane="6" />
                <RESULT eventid="1220" points="290" swimtime="00:01:25.87" resultid="1644" heatid="4386" lane="4" />
                <RESULT eventid="1306" points="332" swimtime="00:00:33.99" resultid="1645" heatid="4479" lane="3" entrytime="00:00:34.86" entrycourse="LCM" />
                <RESULT eventid="1374" points="342" swimtime="00:01:13.76" resultid="1646" heatid="4529" lane="6" entrytime="00:01:13.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Batista Sanchez" birthdate="2009-05-22" gender="M" nation="BRA" license="370668" swrid="5255779" athleteid="1580" externalid="370668">
              <RESULTS>
                <RESULT eventid="1088" points="346" swimtime="00:02:58.67" resultid="1581" heatid="4286" lane="6" entrytime="00:02:55.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="385" swimtime="00:00:35.65" resultid="1582" heatid="4366" lane="4" entrytime="00:00:35.90" entrycourse="LCM" />
                <RESULT eventid="1220" status="DSQ" swimtime="00:00:00.00" resultid="1583" heatid="4392" lane="7" entrytime="00:01:17.76" entrycourse="LCM" />
                <RESULT eventid="1274" points="337" swimtime="00:02:43.72" resultid="1584" heatid="4444" lane="6" entrytime="00:02:52.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="293" swimtime="00:01:14.37" resultid="1585" heatid="4498" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Marques Picolo Vinha" birthdate="2010-07-01" gender="M" nation="BRA" license="366990" swrid="5603869" athleteid="1713" externalid="366990">
              <RESULTS>
                <RESULT eventid="1104" points="243" swimtime="00:00:35.68" resultid="1714" heatid="4299" lane="8" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1156" points="340" swimtime="00:01:07.10" resultid="1715" heatid="4339" lane="8" entrytime="00:01:07.45" entrycourse="LCM" />
                <RESULT eventid="1236" points="328" swimtime="00:00:30.31" resultid="1716" heatid="4414" lane="2" entrytime="00:00:30.22" entrycourse="LCM" />
                <RESULT eventid="1290" points="313" swimtime="00:02:30.13" resultid="1717" heatid="4460" lane="4" entrytime="00:02:43.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="281" swimtime="00:01:18.76" resultid="1718" heatid="4527" lane="2" entrytime="00:01:24.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ghelere" birthdate="2011-04-03" gender="F" nation="BRA" license="368146" swrid="5603843" athleteid="1659" externalid="368146">
              <RESULTS>
                <RESULT eventid="1096" points="295" swimtime="00:00:36.66" resultid="1660" heatid="4292" lane="3" entrytime="00:00:37.46" entrycourse="LCM" />
                <RESULT eventid="1148" points="317" swimtime="00:01:15.77" resultid="1661" heatid="4322" lane="4" entrytime="00:01:15.19" entrycourse="LCM" />
                <RESULT eventid="1228" points="337" swimtime="00:00:33.91" resultid="1662" heatid="4399" lane="2" entrytime="00:00:34.40" entrycourse="LCM" />
                <RESULT eventid="1282" points="316" swimtime="00:02:45.57" resultid="1663" heatid="4450" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="173" swimtime="00:01:39.41" resultid="1664" heatid="4493" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Casavechia Carraro" birthdate="2009-07-28" gender="M" nation="BRA" license="368150" swrid="5384752" athleteid="1562" externalid="368150">
              <RESULTS>
                <RESULT eventid="1104" points="559" swimtime="00:00:27.02" resultid="1563" heatid="4303" lane="2" entrytime="00:00:28.03" entrycourse="LCM" />
                <RESULT eventid="1156" points="620" swimtime="00:00:54.93" resultid="1564" heatid="4347" lane="3" entrytime="00:00:54.99" entrycourse="LCM" />
                <RESULT eventid="1236" points="545" swimtime="00:00:25.59" resultid="1565" heatid="4420" lane="5" entrytime="00:00:25.52" entrycourse="LCM" />
                <RESULT eventid="1290" points="574" swimtime="00:02:02.71" resultid="1566" heatid="4468" lane="3" entrytime="00:02:02.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="561" swimtime="00:00:59.93" resultid="1567" heatid="4504" lane="5" entrytime="00:01:01.47" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanni" lastname="Lazzari Mariotti" birthdate="2006-08-14" gender="M" nation="BRA" license="341929" swrid="5615873" athleteid="1598" externalid="341929">
              <RESULTS>
                <RESULT eventid="1088" points="523" swimtime="00:02:35.67" resultid="1599" heatid="4288" lane="3" entrytime="00:02:36.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="556" swimtime="00:00:31.55" resultid="1600" heatid="4368" lane="3" entrytime="00:00:32.28" entrycourse="LCM" />
                <RESULT eventid="1220" points="536" swimtime="00:01:10.00" resultid="1601" heatid="4394" lane="4" entrytime="00:01:09.42" entrycourse="LCM" />
                <RESULT eventid="1274" points="462" swimtime="00:02:27.38" resultid="1602" heatid="4447" lane="3" entrytime="00:02:25.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Pacheco" birthdate="2006-12-20" gender="M" nation="BRA" license="336850" swrid="5603854" athleteid="1603" externalid="336850">
              <RESULTS>
                <RESULT eventid="1104" points="492" swimtime="00:00:28.20" resultid="1604" heatid="4302" lane="7" entrytime="00:00:28.96" entrycourse="LCM" />
                <RESULT eventid="1140" points="407" swimtime="00:05:27.06" resultid="1605" heatid="4317" lane="6" entrytime="00:05:34.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.86" />
                    <SPLIT distance="200" swimtime="00:02:35.97" />
                    <SPLIT distance="300" swimtime="00:04:13.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="453" swimtime="00:00:27.21" resultid="1606" heatid="4418" lane="8" entrytime="00:00:27.07" entrycourse="LCM" />
                <RESULT eventid="1274" points="412" swimtime="00:02:33.12" resultid="1607" heatid="4446" lane="8" entrytime="00:02:36.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="468" swimtime="00:01:03.65" resultid="1608" heatid="4503" lane="2" entrytime="00:01:04.26" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Campelo" birthdate="2011-09-12" gender="M" nation="BRA" license="366963" swrid="5588742" athleteid="1647" externalid="366963">
              <RESULTS>
                <RESULT eventid="1104" points="402" swimtime="00:00:30.16" resultid="1648" heatid="4300" lane="1" entrytime="00:00:32.30" entrycourse="LCM" />
                <RESULT eventid="1156" points="450" swimtime="00:01:01.11" resultid="1649" heatid="4338" lane="4" entrytime="00:01:07.47" entrycourse="LCM" />
                <RESULT eventid="1236" points="449" swimtime="00:00:27.29" resultid="1650" heatid="4415" lane="5" entrytime="00:00:28.66" entrycourse="LCM" />
                <RESULT eventid="1306" points="399" swimtime="00:00:31.97" resultid="1651" heatid="4479" lane="6" entrytime="00:00:35.18" entrycourse="LCM" />
                <RESULT eventid="1342" points="311" swimtime="00:01:12.98" resultid="1652" heatid="4498" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Chaim" birthdate="2011-05-29" gender="F" nation="BRA" license="370662" swrid="5409721" athleteid="1665" externalid="370662">
              <RESULTS>
                <RESULT eventid="1096" points="233" swimtime="00:00:39.65" resultid="1666" heatid="4292" lane="8" entrytime="00:00:45.43" entrycourse="LCM" />
                <RESULT eventid="1148" points="310" swimtime="00:01:16.38" resultid="1667" heatid="4321" lane="3" entrytime="00:01:23.31" entrycourse="LCM" />
                <RESULT eventid="1228" points="307" swimtime="00:00:34.97" resultid="1668" heatid="4398" lane="2" entrytime="00:00:38.45" entrycourse="LCM" />
                <RESULT eventid="1298" points="243" swimtime="00:00:42.99" resultid="1669" heatid="4471" lane="4" entrytime="00:00:47.61" entrycourse="LCM" />
                <RESULT eventid="1366" points="216" swimtime="00:01:35.49" resultid="1670" heatid="4518" lane="2" entrytime="00:01:39.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Passafaro" birthdate="2009-02-01" gender="F" nation="BRA" license="370673" swrid="5603885" athleteid="1614" externalid="370673">
              <RESULTS>
                <RESULT eventid="1096" points="351" swimtime="00:00:34.61" resultid="1615" heatid="4293" lane="3" entrytime="00:00:34.94" entrycourse="LCM" />
                <RESULT eventid="1148" points="337" swimtime="00:01:14.28" resultid="1616" heatid="4325" lane="6" entrytime="00:01:10.85" entrycourse="LCM" />
                <RESULT eventid="1228" points="416" swimtime="00:00:31.62" resultid="1617" heatid="4403" lane="4" entrytime="00:00:30.34" entrycourse="LCM" />
                <RESULT eventid="1298" points="278" swimtime="00:00:41.11" resultid="1618" heatid="4472" lane="4" entrytime="00:00:41.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Quental De Meireles" birthdate="2008-11-20" gender="M" nation="BRA" license="392103" swrid="5603898" athleteid="1701" externalid="392103">
              <RESULTS>
                <RESULT eventid="1104" points="410" swimtime="00:00:29.96" resultid="1702" heatid="4297" lane="6" />
                <RESULT eventid="1156" points="361" swimtime="00:01:05.79" resultid="1703" heatid="4338" lane="5" entrytime="00:01:07.51" entrycourse="LCM" />
                <RESULT eventid="1188" points="350" swimtime="00:00:36.80" resultid="1704" heatid="4366" lane="8" entrytime="00:00:37.40" entrycourse="LCM" />
                <RESULT eventid="1220" points="297" swimtime="00:01:25.25" resultid="1705" heatid="4391" lane="7" entrytime="00:01:22.80" entrycourse="LCM" />
                <RESULT eventid="1236" points="315" swimtime="00:00:30.71" resultid="1706" heatid="4414" lane="7" entrytime="00:00:30.32" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mochiutti Carneiro" birthdate="2010-04-22" gender="F" nation="BRA" license="370670" swrid="5588817" athleteid="1683" externalid="370670">
              <RESULTS>
                <RESULT eventid="1096" points="403" swimtime="00:00:33.06" resultid="1684" heatid="4294" lane="8" entrytime="00:00:33.10" entrycourse="LCM" />
                <RESULT eventid="1148" points="457" swimtime="00:01:07.12" resultid="1685" heatid="4328" lane="1" entrytime="00:01:06.60" entrycourse="LCM" />
                <RESULT eventid="1228" points="446" swimtime="00:00:30.89" resultid="1686" heatid="4404" lane="7" entrytime="00:00:30.18" entrycourse="LCM" />
                <RESULT eventid="1282" points="456" swimtime="00:02:26.58" resultid="1687" heatid="4455" lane="2" entrytime="00:02:28.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="408" swimtime="00:01:14.76" resultid="1688" heatid="4496" lane="6" entrytime="00:01:17.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Ficher Delmont Pais" birthdate="2010-07-15" gender="M" nation="BRA" license="338533" swrid="5588701" athleteid="1568" externalid="338533">
              <RESULTS>
                <RESULT eventid="1104" points="544" swimtime="00:00:27.28" resultid="1569" heatid="4303" lane="6" entrytime="00:00:27.70" entrycourse="LCM" />
                <RESULT eventid="1156" points="599" swimtime="00:00:55.56" resultid="1570" heatid="4346" lane="7" entrytime="00:00:57.93" entrycourse="LCM" />
                <RESULT eventid="1236" points="511" swimtime="00:00:26.14" resultid="1571" heatid="4419" lane="3" entrytime="00:00:26.36" entrycourse="LCM" />
                <RESULT eventid="1274" points="447" swimtime="00:02:29.09" resultid="1572" heatid="4446" lane="1" entrytime="00:02:36.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="531" swimtime="00:01:01.04" resultid="1573" heatid="4504" lane="6" entrytime="00:01:01.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Antonio Mendes" birthdate="2008-12-04" gender="M" nation="BRA" license="366962" swrid="5196287" athleteid="1619" externalid="366962">
              <RESULTS>
                <RESULT eventid="1088" points="498" swimtime="00:02:38.25" resultid="1620" heatid="4287" lane="2" entrytime="00:02:50.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="587" swimtime="00:00:30.98" resultid="1621" heatid="4368" lane="2" entrytime="00:00:32.84" entrycourse="LCM" />
                <RESULT eventid="1220" points="550" swimtime="00:01:09.42" resultid="1622" heatid="4393" lane="5" entrytime="00:01:12.52" entrycourse="LCM" />
                <RESULT eventid="1274" points="453" swimtime="00:02:28.42" resultid="1623" heatid="4440" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="446" swimtime="00:01:07.53" resultid="1624" heatid="4530" lane="6" entrytime="00:01:10.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Otavio Costa" birthdate="2009-01-28" gender="M" nation="BRA" license="370666" swrid="5603881" athleteid="1671" externalid="370666">
              <RESULTS>
                <RESULT eventid="1088" points="278" swimtime="00:03:12.13" resultid="1672" heatid="4285" lane="1" entrytime="00:03:17.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="282" swimtime="00:00:39.54" resultid="1673" heatid="4365" lane="7" entrytime="00:00:41.24" entrycourse="LCM" />
                <RESULT eventid="1220" points="271" swimtime="00:01:27.83" resultid="1674" heatid="4390" lane="8" entrytime="00:01:30.23" entrycourse="LCM" />
                <RESULT eventid="1236" points="265" swimtime="00:00:32.52" resultid="1675" heatid="4408" lane="4" />
                <RESULT eventid="1274" points="243" swimtime="00:03:02.53" resultid="1676" heatid="4443" lane="1" entrytime="00:03:06.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Donato De Morais" birthdate="2009-03-28" gender="F" nation="BRA" license="345588" swrid="5485198" athleteid="1609" externalid="345588">
              <RESULTS>
                <RESULT eventid="1064" points="365" swimtime="00:02:52.19" resultid="1610" heatid="4270" lane="8" entrytime="00:02:50.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="282" swimtime="00:12:19.06" resultid="1611" heatid="4426" lane="6" entrytime="00:11:36.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.32" />
                    <SPLIT distance="200" swimtime="00:02:49.90" />
                    <SPLIT distance="300" swimtime="00:04:24.70" />
                    <SPLIT distance="400" swimtime="00:06:00.37" />
                    <SPLIT distance="500" swimtime="00:07:36.22" />
                    <SPLIT distance="600" swimtime="00:09:12.81" />
                    <SPLIT distance="700" swimtime="00:10:48.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="400" swimtime="00:00:36.43" resultid="1612" heatid="4474" lane="1" entrytime="00:00:37.48" entrycourse="LCM" />
                <RESULT eventid="1366" points="379" swimtime="00:01:19.17" resultid="1613" heatid="4522" lane="5" entrytime="00:01:18.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Bessa" birthdate="2003-06-19" gender="M" nation="BRA" license="317841" swrid="5312237" athleteid="1558" externalid="317841">
              <RESULTS>
                <RESULT eventid="1088" points="555" swimtime="00:02:32.60" resultid="1559" heatid="4289" lane="7" entrytime="00:02:27.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="689" swimtime="00:00:29.38" resultid="1560" heatid="4369" lane="7" entrytime="00:00:29.55" entrycourse="LCM" />
                <RESULT eventid="1220" points="677" swimtime="00:01:04.77" resultid="1561" heatid="4395" lane="2" entrytime="00:01:05.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Garcia Cavalcante" birthdate="2008-08-11" gender="M" nation="BRA" license="369676" swrid="5603841" athleteid="1586" externalid="369676">
              <RESULTS>
                <RESULT eventid="1088" points="424" swimtime="00:02:47.00" resultid="1587" heatid="4288" lane="1" entrytime="00:02:43.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="405" swimtime="00:00:35.06" resultid="1588" heatid="4366" lane="6" entrytime="00:00:36.34" entrycourse="LCM" />
                <RESULT eventid="1220" points="396" swimtime="00:01:17.42" resultid="1589" heatid="4392" lane="3" entrytime="00:01:16.94" entrycourse="LCM" />
                <RESULT eventid="1274" points="380" swimtime="00:02:37.31" resultid="1590" heatid="4445" lane="2" entrytime="00:02:42.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="399" swimtime="00:04:58.71" resultid="1591" heatid="4512" lane="4" entrytime="00:05:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.71" />
                    <SPLIT distance="200" swimtime="00:02:25.16" />
                    <SPLIT distance="300" swimtime="00:03:41.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1324" points="261" swimtime="00:05:23.55" resultid="1721" heatid="4488" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.29" />
                    <SPLIT distance="200" swimtime="00:02:36.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1647" number="1" />
                    <RELAYPOSITION athleteid="1653" number="2" />
                    <RELAYPOSITION athleteid="1592" number="3" />
                    <RELAYPOSITION athleteid="1689" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1392" points="308" swimtime="00:04:38.72" resultid="1725" heatid="4539" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1647" number="1" />
                    <RELAYPOSITION athleteid="1592" number="2" />
                    <RELAYPOSITION athleteid="1689" number="3" />
                    <RELAYPOSITION athleteid="1653" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1330" points="428" swimtime="00:04:34.34" resultid="1722" heatid="4491" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.38" />
                    <SPLIT distance="200" swimtime="00:02:20.74" />
                    <SPLIT distance="300" swimtime="00:03:31.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1574" number="1" />
                    <RELAYPOSITION athleteid="1619" number="2" />
                    <RELAYPOSITION athleteid="1701" number="3" />
                    <RELAYPOSITION athleteid="1586" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1398" points="452" swimtime="00:04:05.24" resultid="1728" heatid="4542" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.67" />
                    <SPLIT distance="200" swimtime="00:01:58.24" />
                    <SPLIT distance="300" swimtime="00:02:59.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1574" number="1" />
                    <RELAYPOSITION athleteid="1619" number="2" />
                    <RELAYPOSITION athleteid="1586" number="3" />
                    <RELAYPOSITION athleteid="1701" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1328" points="362" swimtime="00:04:50.04" resultid="1723" heatid="4490" lane="5" entrytime="00:04:26.66">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.74" />
                    <SPLIT distance="200" swimtime="00:02:31.46" />
                    <SPLIT distance="300" swimtime="00:03:37.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1562" number="1" />
                    <RELAYPOSITION athleteid="1580" number="2" />
                    <RELAYPOSITION athleteid="1625" number="3" />
                    <RELAYPOSITION athleteid="1671" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1396" points="397" swimtime="00:04:15.94" resultid="1727" heatid="4541" lane="5" entrytime="00:04:00.62">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.39" />
                    <SPLIT distance="200" swimtime="00:01:58.23" />
                    <SPLIT distance="300" swimtime="00:03:10.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1562" number="1" />
                    <RELAYPOSITION athleteid="1625" number="2" />
                    <RELAYPOSITION athleteid="1671" number="3" />
                    <RELAYPOSITION athleteid="1580" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1332" points="540" swimtime="00:04:13.87" resultid="1724" heatid="4492" lane="5" entrytime="00:04:04.97">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.37" />
                    <SPLIT distance="200" swimtime="00:02:11.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1553" number="1" />
                    <RELAYPOSITION athleteid="1558" number="2" />
                    <RELAYPOSITION athleteid="1603" number="3" />
                    <RELAYPOSITION athleteid="1598" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1400" points="566" swimtime="00:03:47.51" resultid="1726" heatid="4543" lane="3" entrytime="00:03:48.18">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1553" number="1" />
                    <RELAYPOSITION athleteid="1603" number="2" />
                    <RELAYPOSITION athleteid="1598" number="3" />
                    <RELAYPOSITION athleteid="1636" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1314" status="DSQ" swimtime="00:05:50.22" resultid="1719" heatid="4483" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.09" />
                    <SPLIT distance="200" swimtime="00:02:59.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1695" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="1707" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="1659" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="1665" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1382" points="330" swimtime="00:05:00.80" resultid="1720" heatid="4534" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1695" number="1" />
                    <RELAYPOSITION athleteid="1659" number="2" />
                    <RELAYPOSITION athleteid="1707" number="3" />
                    <RELAYPOSITION athleteid="1665" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1112" points="336" swimtime="00:05:12.93" resultid="1729" heatid="4306" lane="5" entrytime="00:04:58.04">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.25" />
                    <SPLIT distance="200" swimtime="00:02:48.60" />
                    <SPLIT distance="300" swimtime="00:03:58.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1695" number="1" />
                    <RELAYPOSITION athleteid="1653" number="2" />
                    <RELAYPOSITION athleteid="1647" number="3" />
                    <RELAYPOSITION athleteid="1659" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1114" points="409" swimtime="00:04:52.99" resultid="1730" heatid="4307" lane="2" entrytime="00:04:56.80">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:02:44.40" />
                    <SPLIT distance="300" swimtime="00:03:45.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1677" number="1" />
                    <RELAYPOSITION athleteid="1641" number="2" />
                    <RELAYPOSITION athleteid="1568" number="3" />
                    <RELAYPOSITION athleteid="1683" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1244" points="388" swimtime="00:04:58.24" resultid="1731" heatid="4423" lane="5" entrytime="00:04:38.17">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.43" />
                    <SPLIT distance="200" swimtime="00:02:36.72" />
                    <SPLIT distance="300" swimtime="00:03:42.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1609" number="1" />
                    <RELAYPOSITION athleteid="1580" number="2" />
                    <RELAYPOSITION athleteid="1625" number="3" />
                    <RELAYPOSITION athleteid="1614" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/MARINGÁ &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1112" points="211" swimtime="00:06:05.22" resultid="1732" heatid="4306" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.25" />
                    <SPLIT distance="200" swimtime="00:03:14.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1689" number="1" />
                    <RELAYPOSITION athleteid="1707" number="2" />
                    <RELAYPOSITION athleteid="1592" number="3" />
                    <RELAYPOSITION athleteid="1665" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="11303" nation="BRA" region="PR" clubid="1868" swrid="93760" name="Associação De Talentos Da Natação" shortname="Atn/Curitiba">
          <ATHLETES>
            <ATHLETE firstname="Marcos" lastname="Demchuk" birthdate="2011-06-15" gender="M" nation="BRA" license="388540" swrid="5602530" athleteid="1960" externalid="388540">
              <RESULTS>
                <RESULT eventid="1156" points="234" swimtime="00:01:16.04" resultid="1961" heatid="4335" lane="2" entrytime="00:01:17.76" entrycourse="LCM" />
                <RESULT eventid="1188" points="245" swimtime="00:00:41.45" resultid="1962" heatid="4364" lane="8" entrytime="00:00:50.45" entrycourse="LCM" />
                <RESULT eventid="1220" status="DSQ" swimtime="00:01:34.90" resultid="1963" heatid="4388" lane="7" entrytime="00:01:38.13" entrycourse="LCM" />
                <RESULT eventid="1236" points="282" swimtime="00:00:31.87" resultid="1964" heatid="4411" lane="8" entrytime="00:00:35.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Ocanha" birthdate="2005-06-21" gender="M" nation="BRA" license="313769" swrid="5600231" athleteid="1879" externalid="313769">
              <RESULTS>
                <RESULT eventid="1188" points="582" swimtime="00:00:31.07" resultid="1880" heatid="4369" lane="1" entrytime="00:00:31.13" entrycourse="LCM" />
                <RESULT eventid="1220" points="502" swimtime="00:01:11.56" resultid="1881" heatid="4394" lane="1" entrytime="00:01:11.79" entrycourse="LCM" />
                <RESULT eventid="1236" points="583" swimtime="00:00:25.03" resultid="1882" heatid="4421" lane="5" entrytime="00:00:24.74" entrycourse="LCM" />
                <RESULT eventid="1306" points="459" swimtime="00:00:30.52" resultid="1883" heatid="4476" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Kerniski Demantova" birthdate="1982-05-25" gender="M" nation="BRA" license="398222" swrid="5653293" athleteid="1899" externalid="398222">
              <RESULTS>
                <RESULT eventid="1124" points="385" swimtime="00:10:20.99" resultid="1900" heatid="4311" lane="6" entrytime="00:10:29.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.91" />
                    <SPLIT distance="200" swimtime="00:02:28.51" />
                    <SPLIT distance="300" swimtime="00:03:46.05" />
                    <SPLIT distance="400" swimtime="00:05:04.21" />
                    <SPLIT distance="500" swimtime="00:06:23.85" />
                    <SPLIT distance="600" swimtime="00:07:42.89" />
                    <SPLIT distance="700" swimtime="00:09:02.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="369" swimtime="00:20:14.03" resultid="1901" heatid="4431" lane="3" entrytime="00:20:15.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.49" />
                    <SPLIT distance="200" swimtime="00:02:32.92" />
                    <SPLIT distance="300" swimtime="00:03:54.50" />
                    <SPLIT distance="400" swimtime="00:05:15.19" />
                    <SPLIT distance="500" swimtime="00:06:35.86" />
                    <SPLIT distance="600" swimtime="00:07:56.50" />
                    <SPLIT distance="700" swimtime="00:09:17.47" />
                    <SPLIT distance="800" swimtime="00:10:39.03" />
                    <SPLIT distance="900" swimtime="00:12:01.17" />
                    <SPLIT distance="1000" swimtime="00:13:23.22" />
                    <SPLIT distance="1100" swimtime="00:14:45.15" />
                    <SPLIT distance="1200" swimtime="00:16:07.87" />
                    <SPLIT distance="1300" swimtime="00:17:31.98" />
                    <SPLIT distance="1400" swimtime="00:18:54.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="377" swimtime="00:02:21.08" resultid="1902" heatid="4464" lane="4" entrytime="00:02:20.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="397" swimtime="00:04:59.33" resultid="1903" heatid="4514" lane="2" entrytime="00:05:01.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                    <SPLIT distance="200" swimtime="00:02:26.24" />
                    <SPLIT distance="300" swimtime="00:03:43.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Yuji Yamazato" birthdate="2008-10-01" gender="M" nation="BRA" license="392664" swrid="5622313" athleteid="1986" externalid="392664">
              <RESULTS>
                <RESULT eventid="1104" points="370" swimtime="00:00:31.01" resultid="1987" heatid="4299" lane="6" entrytime="00:00:34.11" entrycourse="LCM" />
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="1988" heatid="4340" lane="2" entrytime="00:01:06.10" entrycourse="LCM" />
                <RESULT eventid="1236" points="373" swimtime="00:00:29.03" resultid="1989" heatid="4415" lane="2" entrytime="00:00:29.48" entrycourse="LCM" />
                <RESULT eventid="1342" points="183" swimtime="00:01:27.05" resultid="1990" heatid="4499" lane="6" entrytime="00:01:29.94" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Angelo" lastname="De Queiroz Neto" birthdate="2003-10-31" gender="M" nation="BRA" license="342814" swrid="5600149" athleteid="1889" externalid="342814">
              <RESULTS>
                <RESULT eventid="1104" points="382" swimtime="00:00:30.67" resultid="1890" heatid="4300" lane="4" entrytime="00:00:30.33" entrycourse="LCM" />
                <RESULT eventid="1156" points="427" swimtime="00:01:02.20" resultid="1891" heatid="4344" lane="1" entrytime="00:01:00.52" entrycourse="LCM" />
                <RESULT eventid="1290" points="395" swimtime="00:02:18.92" resultid="1892" heatid="4465" lane="4" entrytime="00:02:15.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="362" swimtime="00:01:09.33" resultid="1893" heatid="4502" lane="6" entrytime="00:01:07.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Iglesias Prado" birthdate="2010-06-15" gender="M" nation="BRA" license="408052" swrid="5723025" athleteid="2025" externalid="408052">
              <RESULTS>
                <RESULT eventid="1104" points="149" swimtime="00:00:41.95" resultid="2026" heatid="4295" lane="2" />
                <RESULT eventid="1156" points="292" swimtime="00:01:10.59" resultid="2027" heatid="4336" lane="6" entrytime="00:01:12.35" entrycourse="LCM" />
                <RESULT eventid="1236" points="318" swimtime="00:00:30.61" resultid="2028" heatid="4408" lane="6" />
                <RESULT eventid="1290" points="239" swimtime="00:02:44.34" resultid="2029" heatid="4460" lane="2" entrytime="00:02:46.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="170" swimtime="00:01:33.00" resultid="2030" heatid="4526" lane="6" entrytime="00:01:34.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Neves Vianna" birthdate="2007-12-30" gender="F" nation="BRA" license="391106" swrid="5600223" athleteid="1971" externalid="391106">
              <RESULTS>
                <RESULT eventid="1064" points="231" swimtime="00:03:20.61" resultid="1972" heatid="4266" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="123" swimtime="00:00:49.01" resultid="1973" heatid="4292" lane="1" entrytime="00:00:44.66" entrycourse="LCM" />
                <RESULT eventid="1148" points="253" swimtime="00:01:21.68" resultid="1974" heatid="4321" lane="6" entrytime="00:01:23.58" entrycourse="LCM" />
                <RESULT eventid="1282" points="238" swimtime="00:03:02.04" resultid="1975" heatid="4451" lane="7" entrytime="00:03:00.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="223" swimtime="00:01:34.49" resultid="1976" heatid="4518" lane="3" entrytime="00:01:36.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="James" lastname="Roberto Zoschke" birthdate="1976-02-08" gender="M" nation="BRA" license="312251" swrid="5688617" athleteid="1904" externalid="312251">
              <RESULTS>
                <RESULT eventid="1188" points="465" swimtime="00:00:33.49" resultid="1905" heatid="4363" lane="1" />
                <RESULT eventid="1220" points="435" swimtime="00:01:15.05" resultid="1906" heatid="4393" lane="3" entrytime="00:01:14.18" entrycourse="LCM" />
                <RESULT eventid="1274" points="379" swimtime="00:02:37.42" resultid="1907" heatid="4442" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabiana" lastname="Zaleski Dallazem" birthdate="2009-05-16" gender="F" nation="BRA" license="344287" swrid="5600279" athleteid="1869" externalid="344287">
              <RESULTS>
                <RESULT eventid="1064" points="480" swimtime="00:02:37.25" resultid="1870" heatid="4271" lane="2" entrytime="00:02:38.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="488" swimtime="00:01:05.65" resultid="1871" heatid="4328" lane="5" entrytime="00:01:05.60" entrycourse="LCM" />
                <RESULT eventid="1298" points="546" swimtime="00:00:32.86" resultid="1872" heatid="4475" lane="6" entrytime="00:00:32.81" entrycourse="LCM" />
                <RESULT eventid="1366" points="497" swimtime="00:01:12.36" resultid="1873" heatid="4524" lane="2" entrytime="00:01:10.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Camila" lastname="Duarte De Almeida" birthdate="2009-11-26" gender="F" nation="BRA" license="378819" swrid="5600152" athleteid="1948" externalid="378819">
              <RESULTS>
                <RESULT eventid="1096" points="349" swimtime="00:00:34.69" resultid="1949" heatid="4293" lane="2" entrytime="00:00:36.70" entrycourse="LCM" />
                <RESULT eventid="1148" points="470" swimtime="00:01:06.47" resultid="1950" heatid="4327" lane="3" entrytime="00:01:07.85" entrycourse="LCM" />
                <RESULT eventid="1228" points="474" swimtime="00:00:30.26" resultid="1951" heatid="4402" lane="4" entrytime="00:00:31.04" entrycourse="LCM" />
                <RESULT eventid="1282" points="419" swimtime="00:02:30.73" resultid="1952" heatid="4453" lane="3" entrytime="00:02:34.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="233" swimtime="00:01:30.04" resultid="1953" heatid="4494" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Kerppers Kreia" birthdate="2006-12-01" gender="M" nation="BRA" license="366815" swrid="5600195" athleteid="1894" externalid="366815">
              <RESULTS>
                <RESULT eventid="1156" points="509" swimtime="00:00:58.68" resultid="1895" heatid="4345" lane="2" entrytime="00:00:59.28" entrycourse="LCM" />
                <RESULT eventid="1236" points="437" swimtime="00:00:27.54" resultid="1896" heatid="4417" lane="2" entrytime="00:00:27.47" entrycourse="LCM" />
                <RESULT eventid="1290" points="460" swimtime="00:02:12.05" resultid="1897" heatid="4467" lane="8" entrytime="00:02:11.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="425" swimtime="00:04:52.61" resultid="1898" heatid="4514" lane="6" entrytime="00:05:01.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.38" />
                    <SPLIT distance="200" swimtime="00:02:24.99" />
                    <SPLIT distance="300" swimtime="00:03:40.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Araujo Do Rego Barros" birthdate="2009-04-30" gender="M" nation="BRA" license="376325" swrid="5377739" athleteid="1930" externalid="376325">
              <RESULTS>
                <RESULT eventid="1104" points="313" swimtime="00:00:32.77" resultid="1931" heatid="4299" lane="1" entrytime="00:00:34.74" entrycourse="LCM" />
                <RESULT eventid="1156" points="303" swimtime="00:01:09.76" resultid="1932" heatid="4338" lane="2" entrytime="00:01:08.19" entrycourse="LCM" />
                <RESULT eventid="1172" points="224" swimtime="00:03:01.49" resultid="1933" heatid="4352" lane="7" entrytime="00:02:59.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="280" swimtime="00:02:35.75" resultid="1934" heatid="4461" lane="6" entrytime="00:02:39.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="289" swimtime="00:01:14.73" resultid="1935" heatid="4500" lane="5" entrytime="00:01:16.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Garcia Fraga" birthdate="2003-10-07" gender="M" nation="BRA" license="283467" swrid="5717265" athleteid="1884" externalid="283467">
              <RESULTS>
                <RESULT eventid="1072" points="435" swimtime="00:02:27.63" resultid="1885" heatid="4272" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="458" swimtime="00:01:13.75" resultid="1886" heatid="4385" lane="4" />
                <RESULT eventid="1274" points="511" swimtime="00:02:22.54" resultid="1887" heatid="4440" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="440" swimtime="00:01:04.97" resultid="1888" heatid="4503" lane="1" entrytime="00:01:04.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Dallastra" birthdate="2010-08-21" gender="M" nation="BRA" license="408024" swrid="5723028" athleteid="2013" externalid="408024">
              <RESULTS>
                <RESULT eventid="1104" points="236" swimtime="00:00:35.99" resultid="2014" heatid="4295" lane="3" />
                <RESULT eventid="1156" points="299" swimtime="00:01:10.02" resultid="2015" heatid="4336" lane="5" entrytime="00:01:11.52" entrycourse="LCM" />
                <RESULT eventid="1236" points="266" swimtime="00:00:32.49" resultid="2016" heatid="4409" lane="8" />
                <RESULT eventid="1290" points="275" swimtime="00:02:36.69" resultid="2017" heatid="4462" lane="2" entrytime="00:02:33.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" status="DNS" swimtime="00:00:00.00" resultid="2018" heatid="4498" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Bortoleto" birthdate="2008-09-05" gender="M" nation="BRA" license="406709" swrid="5717249" athleteid="1995" externalid="406709">
              <RESULTS>
                <RESULT eventid="1104" points="368" swimtime="00:00:31.05" resultid="1996" heatid="4296" lane="3" />
                <RESULT eventid="1156" points="411" swimtime="00:01:02.99" resultid="1997" heatid="4341" lane="3" entrytime="00:01:04.50" entrycourse="LCM" />
                <RESULT eventid="1236" points="417" swimtime="00:00:27.97" resultid="1998" heatid="4409" lane="3" />
                <RESULT eventid="1290" points="363" swimtime="00:02:22.94" resultid="1999" heatid="4458" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="334" swimtime="00:01:11.23" resultid="2000" heatid="4501" lane="4" entrytime="00:01:13.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelo" lastname="Correia Bonfim" birthdate="2009-06-21" gender="M" nation="BRA" license="391663" swrid="5622271" athleteid="1977" externalid="391663">
              <RESULTS>
                <RESULT eventid="1104" points="343" swimtime="00:00:31.80" resultid="1978" heatid="4296" lane="8" />
                <RESULT eventid="1156" points="424" swimtime="00:01:02.36" resultid="1979" heatid="4342" lane="1" entrytime="00:01:03.44" entrycourse="LCM" />
                <RESULT eventid="1236" points="416" swimtime="00:00:28.01" resultid="1980" heatid="4407" lane="4" />
                <RESULT eventid="1274" points="338" swimtime="00:02:43.64" resultid="1981" heatid="4443" lane="4" entrytime="00:02:59.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="325" swimtime="00:01:15.01" resultid="1982" heatid="4525" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Garcia De Fraga" birthdate="2009-03-24" gender="M" nation="BRA" license="342147" swrid="5600172" athleteid="1874" externalid="342147">
              <RESULTS>
                <RESULT eventid="1072" points="574" swimtime="00:02:14.61" resultid="1875" heatid="4277" lane="6" entrytime="00:02:17.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="512" swimtime="00:05:02.95" resultid="1876" heatid="4318" lane="2" entrytime="00:05:02.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.31" />
                    <SPLIT distance="200" swimtime="00:02:21.89" />
                    <SPLIT distance="300" swimtime="00:03:51.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1274" points="579" swimtime="00:02:16.76" resultid="1877" heatid="4448" lane="2" entrytime="00:02:16.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="577" swimtime="00:01:01.98" resultid="1878" heatid="4533" lane="8" entrytime="00:01:01.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Zaleski Dallazem" birthdate="2009-05-16" gender="M" nation="BRA" license="344286" swrid="5600280" athleteid="1913" externalid="344286">
              <RESULTS>
                <RESULT eventid="1088" points="382" swimtime="00:02:52.91" resultid="1914" heatid="4286" lane="5" entrytime="00:02:53.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="457" swimtime="00:01:00.82" resultid="1915" heatid="4332" lane="1" />
                <RESULT eventid="1220" points="390" swimtime="00:01:17.82" resultid="1916" heatid="4392" lane="2" entrytime="00:01:17.44" entrycourse="LCM" />
                <RESULT eventid="1236" points="411" swimtime="00:00:28.11" resultid="1917" heatid="4414" lane="5" entrytime="00:00:30.14" entrycourse="LCM" />
                <RESULT eventid="1274" points="384" swimtime="00:02:36.75" resultid="1918" heatid="4445" lane="8" entrytime="00:02:47.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Faria Del Valle" birthdate="2009-08-28" gender="M" nation="BRA" license="376328" swrid="5600155" athleteid="1936" externalid="376328">
              <RESULTS>
                <RESULT eventid="1156" points="535" swimtime="00:00:57.69" resultid="1937" heatid="4345" lane="1" entrytime="00:00:59.47" entrycourse="LCM" />
                <RESULT eventid="1188" points="438" swimtime="00:00:34.15" resultid="1938" heatid="4366" lane="2" entrytime="00:00:36.50" entrycourse="LCM" />
                <RESULT eventid="1236" points="551" swimtime="00:00:25.50" resultid="1939" heatid="4419" lane="4" entrytime="00:00:26.20" entrycourse="LCM" />
                <RESULT eventid="1306" points="419" swimtime="00:00:31.45" resultid="1940" heatid="4480" lane="3" entrytime="00:00:32.28" entrycourse="LCM" />
                <RESULT eventid="1374" points="392" swimtime="00:01:10.48" resultid="1941" heatid="4529" lane="2" entrytime="00:01:13.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Castellano Purkot" birthdate="2010-01-25" gender="M" nation="BRA" license="392484" swrid="5622268" athleteid="1983" externalid="392484">
              <RESULTS>
                <RESULT eventid="1236" points="268" swimtime="00:00:32.42" resultid="1984" heatid="4414" lane="8" entrytime="00:00:30.44" entrycourse="LCM" />
                <RESULT eventid="1306" points="168" swimtime="00:00:42.61" resultid="1985" heatid="4476" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Fonseca Vendramin" birthdate="2008-09-28" gender="F" nation="BRA" license="393918" swrid="5622282" athleteid="1991" externalid="393918">
              <RESULTS>
                <RESULT eventid="1096" points="303" swimtime="00:00:36.37" resultid="1992" heatid="4292" lane="5" entrytime="00:00:37.29" entrycourse="LCM" />
                <RESULT eventid="1228" status="DSQ" swimtime="00:00:31.62" resultid="1993" heatid="4400" lane="2" entrytime="00:00:33.06" entrycourse="LCM" />
                <RESULT eventid="1334" points="226" swimtime="00:01:31.03" resultid="1994" heatid="4495" lane="5" entrytime="00:01:25.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Freitas Szucs" birthdate="2011-10-02" gender="M" nation="BRA" license="377272" swrid="5588708" athleteid="1919" externalid="377272">
              <RESULTS>
                <RESULT eventid="1104" points="182" swimtime="00:00:39.25" resultid="1920" heatid="4298" lane="1" entrytime="00:00:41.08" entrycourse="LCM" />
                <RESULT eventid="1156" points="208" swimtime="00:01:19.06" resultid="1921" heatid="4335" lane="1" entrytime="00:01:18.83" entrycourse="LCM" />
                <RESULT eventid="1236" points="215" swimtime="00:00:34.87" resultid="1922" heatid="4411" lane="1" entrytime="00:00:35.74" entrycourse="LCM" />
                <RESULT eventid="1290" points="196" swimtime="00:02:55.38" resultid="1923" heatid="4460" lane="1" entrytime="00:02:58.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Sofia Silva" birthdate="2007-05-28" gender="F" nation="BRA" license="390921" swrid="5600260" athleteid="1965" externalid="390921">
              <RESULTS>
                <RESULT eventid="1080" points="235" swimtime="00:03:42.87" resultid="1966" heatid="4278" lane="2" entrytime="00:04:15.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="226" swimtime="00:01:24.78" resultid="1967" heatid="4319" lane="6" />
                <RESULT eventid="1180" points="205" swimtime="00:00:49.39" resultid="1968" heatid="4356" lane="6" entrytime="00:00:50.90" entrycourse="LCM" />
                <RESULT eventid="1212" points="236" swimtime="00:01:43.68" resultid="1969" heatid="4379" lane="6" entrytime="00:01:51.65" entrycourse="LCM" />
                <RESULT eventid="1266" points="238" swimtime="00:03:23.23" resultid="1970" heatid="4435" lane="6" entrytime="00:03:40.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Riccieri" lastname="Rodrigues Muzolon" birthdate="2010-11-08" gender="M" nation="BRA" license="385439" swrid="5588887" athleteid="1954" externalid="385439">
              <RESULTS>
                <RESULT eventid="1072" points="273" swimtime="00:02:52.41" resultid="1955" heatid="4272" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="283" swimtime="00:00:33.92" resultid="1956" heatid="4298" lane="3" entrytime="00:00:37.64" entrycourse="LCM" />
                <RESULT eventid="1156" points="332" swimtime="00:01:07.61" resultid="1957" heatid="4337" lane="4" entrytime="00:01:09.08" entrycourse="LCM" />
                <RESULT eventid="1290" status="DNS" swimtime="00:00:00.00" resultid="1958" heatid="4461" lane="7" entrytime="00:02:40.53" entrycourse="LCM" />
                <RESULT eventid="1374" status="DNS" swimtime="00:00:00.00" resultid="1959" heatid="4527" lane="5" entrytime="00:01:22.03" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Navarro Silva" birthdate="2011-01-10" gender="F" nation="BRA" license="406711" swrid="5717284" athleteid="2001" externalid="406711">
              <RESULTS>
                <RESULT eventid="1064" points="287" swimtime="00:03:06.63" resultid="2002" heatid="4267" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="295" swimtime="00:01:17.63" resultid="2003" heatid="4320" lane="8" />
                <RESULT eventid="1228" points="274" swimtime="00:00:36.33" resultid="2004" heatid="4397" lane="6" />
                <RESULT eventid="1282" points="281" swimtime="00:02:52.27" resultid="2005" heatid="4451" lane="6" entrytime="00:02:53.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="283" swimtime="00:01:27.27" resultid="2006" heatid="4519" lane="3" entrytime="00:01:29.62" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mauricio" lastname="Furtado Niwa" birthdate="1978-05-30" gender="M" nation="BRA" license="398757" swrid="5653291" athleteid="1908" externalid="398757">
              <RESULTS>
                <RESULT eventid="1172" points="366" swimtime="00:02:34.18" resultid="1909" heatid="4353" lane="3" entrytime="00:02:31.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="473" swimtime="00:00:26.83" resultid="1910" heatid="4410" lane="7" />
                <RESULT eventid="1290" points="461" swimtime="00:02:11.96" resultid="1911" heatid="4458" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="501" swimtime="00:01:02.26" resultid="1912" heatid="4504" lane="2" entrytime="00:01:01.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Arthur Ribeiro" birthdate="2010-02-05" gender="M" nation="BRA" license="408025" swrid="5723020" athleteid="2019" externalid="408025">
              <RESULTS>
                <RESULT eventid="1104" points="212" swimtime="00:00:37.30" resultid="2020" heatid="4296" lane="7" />
                <RESULT eventid="1156" points="257" swimtime="00:01:13.61" resultid="2021" heatid="4335" lane="8" entrytime="00:01:19.52" entrycourse="LCM" />
                <RESULT eventid="1188" points="298" swimtime="00:00:38.85" resultid="2022" heatid="4360" lane="3" />
                <RESULT eventid="1220" points="249" swimtime="00:01:30.36" resultid="2023" heatid="4388" lane="2" entrytime="00:01:35.86" entrycourse="LCM" />
                <RESULT eventid="1236" points="266" swimtime="00:00:32.49" resultid="2024" heatid="4406" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jhon" lastname="Caleb Dos Santos" birthdate="2010-03-02" gender="M" nation="BRA" license="359020" swrid="5588574" athleteid="1924" externalid="359020">
              <RESULTS>
                <RESULT eventid="1140" points="437" swimtime="00:05:19.42" resultid="1925" heatid="4317" lane="3" entrytime="00:05:24.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.26" />
                    <SPLIT distance="200" swimtime="00:02:34.07" />
                    <SPLIT distance="300" swimtime="00:04:08.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="386" swimtime="00:01:18.08" resultid="1926" heatid="4392" lane="1" entrytime="00:01:18.40" entrycourse="LCM" />
                <RESULT eventid="1274" points="442" swimtime="00:02:29.55" resultid="1927" heatid="4446" lane="4" entrytime="00:02:31.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="427" swimtime="00:01:05.62" resultid="1928" heatid="4502" lane="5" entrytime="00:01:05.68" entrycourse="LCM" />
                <RESULT eventid="1374" points="377" swimtime="00:01:11.40" resultid="1929" heatid="4526" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Inacio Carneiro" birthdate="2009-09-09" gender="M" nation="BRA" license="408023" swrid="5723026" athleteid="2007" externalid="408023">
              <RESULTS>
                <RESULT eventid="1156" points="252" swimtime="00:01:14.10" resultid="2008" heatid="4336" lane="1" entrytime="00:01:14.15" entrycourse="LCM" />
                <RESULT eventid="1236" points="298" swimtime="00:00:31.29" resultid="2009" heatid="4407" lane="2" />
                <RESULT eventid="1290" points="212" swimtime="00:02:50.93" resultid="2010" heatid="4460" lane="7" entrytime="00:02:57.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1306" points="146" swimtime="00:00:44.69" resultid="2011" heatid="4476" lane="8" />
                <RESULT eventid="1374" status="DSQ" swimtime="00:01:38.86" resultid="2012" heatid="4526" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Muller" birthdate="2009-10-10" gender="F" nation="BRA" license="376952" swrid="5600221" athleteid="1942" externalid="376952">
              <RESULTS>
                <RESULT eventid="1080" points="434" swimtime="00:03:01.63" resultid="1943" heatid="4281" lane="4" entrytime="00:02:59.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="471" swimtime="00:00:37.46" resultid="1944" heatid="4359" lane="6" entrytime="00:00:36.62" entrycourse="LCM" />
                <RESULT eventid="1212" points="452" swimtime="00:01:23.56" resultid="1945" heatid="4384" lane="8" entrytime="00:01:21.69" entrycourse="LCM" />
                <RESULT eventid="1298" points="261" swimtime="00:00:41.99" resultid="1946" heatid="4473" lane="2" entrytime="00:00:40.07" entrycourse="LCM" />
                <RESULT eventid="1266" points="376" swimtime="00:02:54.67" resultid="1947" heatid="4436" lane="6" entrytime="00:03:06.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="20" agetotalmax="-1" agetotalmin="-1" gender="M" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1210" points="429" swimtime="00:09:14.71" resultid="2033" heatid="4376" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.67" />
                    <SPLIT distance="300" swimtime="00:03:17.35" />
                    <SPLIT distance="400" swimtime="00:04:32.03" />
                    <SPLIT distance="500" swimtime="00:05:38.54" />
                    <SPLIT distance="600" swimtime="00:06:48.27" />
                    <SPLIT distance="700" swimtime="00:07:59.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1884" number="1" />
                    <RELAYPOSITION athleteid="1889" number="2" />
                    <RELAYPOSITION athleteid="1908" number="3" />
                    <RELAYPOSITION athleteid="1899" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1326" points="278" swimtime="00:05:16.56" resultid="2034" heatid="4489" lane="3" entrytime="00:04:46.17">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.47" />
                    <SPLIT distance="200" swimtime="00:02:59.64" />
                    <SPLIT distance="300" swimtime="00:04:05.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1983" number="1" />
                    <RELAYPOSITION athleteid="2019" number="2" />
                    <RELAYPOSITION athleteid="1924" number="3" />
                    <RELAYPOSITION athleteid="2025" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1394" points="339" swimtime="00:04:29.96" resultid="2037" heatid="4540" lane="5" entrytime="00:04:20.49">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.85" />
                    <SPLIT distance="200" swimtime="00:02:11.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1924" number="1" />
                    <RELAYPOSITION athleteid="2019" number="2" />
                    <RELAYPOSITION athleteid="2013" number="3" />
                    <RELAYPOSITION athleteid="2025" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1328" points="434" swimtime="00:04:32.98" resultid="2035" heatid="4490" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.06" />
                    <SPLIT distance="200" swimtime="00:02:32.23" />
                    <SPLIT distance="300" swimtime="00:03:33.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1977" number="1" />
                    <RELAYPOSITION athleteid="1913" number="2" />
                    <RELAYPOSITION athleteid="1874" number="3" />
                    <RELAYPOSITION athleteid="1936" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1396" points="493" swimtime="00:03:58.28" resultid="2039" heatid="4541" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.52" />
                    <SPLIT distance="200" swimtime="00:01:58.70" />
                    <SPLIT distance="300" swimtime="00:02:56.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1913" number="1" />
                    <RELAYPOSITION athleteid="1874" number="2" />
                    <RELAYPOSITION athleteid="1936" number="3" />
                    <RELAYPOSITION athleteid="1977" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1332" points="503" swimtime="00:04:19.97" resultid="2036" heatid="4492" lane="6" entrytime="00:04:55.22">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.14" />
                    <SPLIT distance="200" swimtime="00:02:22.02" />
                    <SPLIT distance="300" swimtime="00:03:25.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1884" number="1" />
                    <RELAYPOSITION athleteid="1904" number="2" />
                    <RELAYPOSITION athleteid="1908" number="3" />
                    <RELAYPOSITION athleteid="1879" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1400" points="507" swimtime="00:03:56.02" resultid="2038" heatid="4543" lane="2" entrytime="00:04:07.59">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.50" />
                    <SPLIT distance="200" swimtime="00:01:55.91" />
                    <SPLIT distance="300" swimtime="00:02:53.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1884" number="1" />
                    <RELAYPOSITION athleteid="1894" number="2" />
                    <RELAYPOSITION athleteid="1908" number="3" />
                    <RELAYPOSITION athleteid="1889" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1320" points="406" swimtime="00:05:11.02" resultid="2031" heatid="4486" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.71" />
                    <SPLIT distance="200" swimtime="00:02:38.41" />
                    <SPLIT distance="300" swimtime="00:04:04.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1869" number="1" />
                    <RELAYPOSITION athleteid="1942" number="2" />
                    <RELAYPOSITION athleteid="1991" number="3" />
                    <RELAYPOSITION athleteid="1948" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1388" status="DSQ" swimtime="00:04:34.86" resultid="2032" heatid="4537" lane="5" entrytime="00:05:32.92">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.53" />
                    <SPLIT distance="200" swimtime="00:02:12.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1948" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="1869" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="1991" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="1942" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1248" points="291" swimtime="00:05:28.20" resultid="2040" heatid="4425" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.47" />
                    <SPLIT distance="200" swimtime="00:03:18.08" />
                    <SPLIT distance="300" swimtime="00:04:28.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1971" number="1" />
                    <RELAYPOSITION athleteid="1965" number="2" />
                    <RELAYPOSITION athleteid="1889" number="3" />
                    <RELAYPOSITION athleteid="1894" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1244" points="499" swimtime="00:04:34.31" resultid="2041" heatid="4423" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.18" />
                    <SPLIT distance="200" swimtime="00:02:35.59" />
                    <SPLIT distance="300" swimtime="00:03:35.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1869" number="1" />
                    <RELAYPOSITION athleteid="1942" number="2" />
                    <RELAYPOSITION athleteid="1874" number="3" />
                    <RELAYPOSITION athleteid="1936" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="2539" nation="BRA" region="PR" clubid="2186" swrid="93771" name="Círculo Militar Do Paraná" shortname="Círculo Militar">
          <ATHLETES>
            <ATHLETE firstname="Nathan" lastname="Torres Oliveira" birthdate="2008-04-10" gender="M" nation="BRA" license="400274" swrid="5653303" athleteid="2212" externalid="400274">
              <RESULTS>
                <RESULT eventid="1088" points="235" swimtime="00:03:23.13" resultid="2213" heatid="4284" lane="5" entrytime="00:03:25.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="314" swimtime="00:01:08.93" resultid="2214" heatid="4338" lane="1" entrytime="00:01:08.46" entrycourse="LCM" />
                <RESULT eventid="1188" points="273" swimtime="00:00:39.96" resultid="2215" heatid="4365" lane="8" entrytime="00:00:41.48" entrycourse="LCM" />
                <RESULT eventid="1220" points="251" swimtime="00:01:30.10" resultid="2216" heatid="4389" lane="5" entrytime="00:01:30.32" entrycourse="LCM" />
                <RESULT eventid="1236" points="365" swimtime="00:00:29.24" resultid="2217" heatid="4414" lane="1" entrytime="00:00:30.44" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Maria Romanelli" birthdate="2011-04-18" gender="F" nation="BRA" license="378335" swrid="5588803" athleteid="2198" externalid="378335">
              <RESULTS>
                <RESULT eventid="1148" points="402" swimtime="00:01:10.02" resultid="2199" heatid="4325" lane="1" entrytime="00:01:11.42" entrycourse="LCM" />
                <RESULT eventid="1180" points="225" swimtime="00:00:47.90" resultid="2200" heatid="4356" lane="4" entrytime="00:00:48.39" entrycourse="LCM" />
                <RESULT eventid="1228" points="378" swimtime="00:00:32.63" resultid="2201" heatid="4400" lane="8" entrytime="00:00:33.27" entrycourse="LCM" />
                <RESULT eventid="1298" points="249" swimtime="00:00:42.66" resultid="2202" heatid="4472" lane="5" entrytime="00:00:41.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Cavalcante Pierin" birthdate="2010-12-28" gender="M" nation="BRA" license="391227" swrid="5622269" athleteid="2209" externalid="391227">
              <RESULTS>
                <RESULT eventid="1156" points="252" swimtime="00:01:14.12" resultid="2210" heatid="4335" lane="5" entrytime="00:01:16.19" entrycourse="LCM" />
                <RESULT eventid="1188" points="172" swimtime="00:00:46.66" resultid="2211" heatid="4361" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Vieira De Macedo Brasil" birthdate="2009-12-19" gender="F" nation="BRA" license="344143" swrid="5622311" athleteid="2190" externalid="344143">
              <RESULTS>
                <RESULT eventid="1228" points="399" swimtime="00:00:32.05" resultid="2191" heatid="4400" lane="5" entrytime="00:00:32.80" entrycourse="LCM" />
                <RESULT eventid="1282" points="384" swimtime="00:02:35.25" resultid="2192" heatid="4453" lane="1" entrytime="00:02:36.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" status="DSQ" swimtime="00:03:12.59" resultid="2193" heatid="4434" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Yamamoto" birthdate="2006-04-22" gender="M" nation="BRA" license="336569" swrid="5717304" athleteid="2187" externalid="336569">
              <RESULTS>
                <RESULT eventid="1236" points="432" swimtime="00:00:27.65" resultid="2188" heatid="4409" lane="5" />
                <RESULT eventid="1306" points="285" swimtime="00:00:35.75" resultid="2189" heatid="4476" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernando" lastname="Jun Melo Ogima" birthdate="2006-07-05" gender="M" nation="BRA" license="378332" swrid="5622284" athleteid="2194" externalid="378332">
              <RESULTS>
                <RESULT eventid="1156" points="413" swimtime="00:01:02.91" resultid="2195" heatid="4342" lane="3" entrytime="00:01:02.12" entrycourse="LCM" />
                <RESULT eventid="1220" points="261" swimtime="00:01:28.95" resultid="2196" heatid="4390" lane="7" entrytime="00:01:27.49" entrycourse="LCM" />
                <RESULT eventid="1274" points="272" swimtime="00:02:55.75" resultid="2197" heatid="4443" lane="5" entrytime="00:03:00.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Manocchio" birthdate="2011-07-28" gender="M" nation="BRA" license="384916" swrid="5588573" athleteid="2203" externalid="384916">
              <RESULTS>
                <RESULT eventid="1156" points="345" swimtime="00:01:06.81" resultid="2204" heatid="4339" lane="6" entrytime="00:01:06.82" entrycourse="LCM" />
                <RESULT eventid="1220" points="223" swimtime="00:01:33.76" resultid="2205" heatid="4388" lane="6" entrytime="00:01:34.96" entrycourse="LCM" />
                <RESULT eventid="1236" points="311" swimtime="00:00:30.84" resultid="2206" heatid="4412" lane="3" entrytime="00:00:31.69" entrycourse="LCM" />
                <RESULT eventid="1290" points="315" swimtime="00:02:29.82" resultid="2207" heatid="4463" lane="2" entrytime="00:02:27.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="330" swimtime="00:05:18.44" resultid="2208" heatid="4512" lane="6" entrytime="00:05:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.27" />
                    <SPLIT distance="200" swimtime="00:02:36.84" />
                    <SPLIT distance="300" swimtime="00:04:00.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thomas" lastname="Gomes" birthdate="2009-06-15" gender="M" nation="BRA" license="406948" swrid="5717268" athleteid="2218" externalid="406948">
              <RESULTS>
                <RESULT eventid="1156" points="216" swimtime="00:01:18.05" resultid="2219" heatid="4334" lane="4" entrytime="00:01:20.37" entrycourse="LCM" />
                <RESULT eventid="1236" points="207" swimtime="00:00:35.30" resultid="2220" heatid="4408" lane="5" />
                <RESULT eventid="1290" points="184" swimtime="00:02:59.25" resultid="2221" heatid="4460" lane="8" entrytime="00:03:01.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vicente" lastname="Bileski" birthdate="2011-06-29" gender="M" nation="BRA" license="406950" swrid="5717248" athleteid="2222" externalid="406950">
              <RESULTS>
                <RESULT eventid="1104" points="139" swimtime="00:00:42.95" resultid="2223" heatid="4297" lane="2" />
                <RESULT eventid="1156" points="182" swimtime="00:01:22.57" resultid="2224" heatid="4334" lane="6" entrytime="00:01:24.86" entrycourse="LCM" />
                <RESULT eventid="1188" points="154" swimtime="00:00:48.33" resultid="2225" heatid="4360" lane="5" />
                <RESULT eventid="1220" points="140" swimtime="00:01:49.51" resultid="2226" heatid="4387" lane="2" entrytime="00:01:49.98" entrycourse="LCM" />
                <RESULT eventid="1236" points="170" swimtime="00:00:37.69" resultid="2227" heatid="4406" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="12782" nation="BRA" region="PR" clubid="3058" swrid="93773" name="Clube Duque De Caxias" shortname="Duque De Caxias">
          <ATHLETES>
            <ATHLETE firstname="Lucas" lastname="Bulgarelli Castro" birthdate="2009-04-20" gender="M" nation="BRA" license="401867" swrid="5658058" athleteid="3074" externalid="401867">
              <RESULTS>
                <RESULT eventid="1156" points="342" swimtime="00:01:06.99" resultid="3075" heatid="4338" lane="3" entrytime="00:01:07.54" entrycourse="LCM" />
                <RESULT eventid="1188" status="DNS" swimtime="00:00:00.00" resultid="3076" heatid="4363" lane="3" />
                <RESULT eventid="1236" points="333" swimtime="00:00:30.15" resultid="3077" heatid="4413" lane="3" entrytime="00:00:30.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Vitor Girelli" birthdate="2009-08-01" gender="M" nation="BRA" license="387965" swrid="5622312" athleteid="3064" externalid="387965">
              <RESULTS>
                <RESULT eventid="1104" points="320" swimtime="00:00:32.55" resultid="3065" heatid="4299" lane="3" entrytime="00:00:33.51" entrycourse="LCM" />
                <RESULT eventid="1156" points="413" swimtime="00:01:02.90" resultid="3066" heatid="4342" lane="2" entrytime="00:01:02.36" entrycourse="LCM" />
                <RESULT eventid="1236" points="372" swimtime="00:00:29.06" resultid="3067" heatid="4415" lane="7" entrytime="00:00:29.55" entrycourse="LCM" />
                <RESULT eventid="1306" points="294" swimtime="00:00:35.39" resultid="3068" heatid="4479" lane="7" entrytime="00:00:35.71" entrycourse="LCM" />
                <RESULT eventid="1374" status="DNS" swimtime="00:00:00.00" resultid="3069" heatid="4528" lane="5" entrytime="00:01:15.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Flavia Braz" birthdate="2004-10-25" gender="F" nation="BRA" license="280573" swrid="5622281" athleteid="3059" externalid="280573">
              <RESULTS>
                <RESULT eventid="1080" points="405" swimtime="00:03:05.80" resultid="3060" heatid="4280" lane="7" entrytime="00:03:14.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="336" swimtime="00:00:35.14" resultid="3061" heatid="4291" lane="8" />
                <RESULT eventid="1228" points="467" swimtime="00:00:30.42" resultid="3062" heatid="4396" lane="1" />
                <RESULT eventid="1212" points="454" swimtime="00:01:23.43" resultid="3063" heatid="4383" lane="7" entrytime="00:01:24.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Bochi Conte" birthdate="2009-04-20" gender="M" nation="BRA" license="401868" swrid="5658057" athleteid="3078" externalid="401868">
              <RESULTS>
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="3079" heatid="4333" lane="6" />
                <RESULT eventid="1236" points="305" swimtime="00:00:31.04" resultid="3080" heatid="4413" lane="7" entrytime="00:00:31.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ian" lastname="Berger" birthdate="2011-07-27" gender="M" nation="BRA" license="387966" swrid="5652879" athleteid="3070" externalid="387966">
              <RESULTS>
                <RESULT eventid="1156" points="268" swimtime="00:01:12.61" resultid="3071" heatid="4336" lane="8" entrytime="00:01:14.95" entrycourse="LCM" />
                <RESULT eventid="1188" points="178" swimtime="00:00:46.07" resultid="3072" heatid="4361" lane="6" />
                <RESULT eventid="1236" points="254" swimtime="00:00:33.00" resultid="3073" heatid="4411" lane="3" entrytime="00:00:34.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3501" nation="BRA" region="PR" clubid="1812" swrid="93752" name="Ortega &amp; De Souza Jesus" shortname="Aquafoz">
          <ATHLETES>
            <ATHLETE firstname="Julio" lastname="Heck" birthdate="1998-02-15" gender="M" nation="BRA" license="185880" swrid="5596906" athleteid="1825" externalid="185880">
              <RESULTS>
                <RESULT eventid="1104" points="534" swimtime="00:00:27.44" resultid="1826" heatid="4296" lane="2" />
                <RESULT eventid="1156" points="635" swimtime="00:00:54.49" resultid="1827" heatid="4348" lane="8" entrytime="00:00:53.71" entrycourse="LCM" />
                <RESULT eventid="1236" points="612" swimtime="00:00:24.62" resultid="1828" heatid="4422" lane="1" entrytime="00:00:24.19" entrycourse="LCM" />
                <RESULT eventid="1306" points="415" swimtime="00:00:31.55" resultid="1829" heatid="4480" lane="6" entrytime="00:00:32.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Dominguez Olivieski" birthdate="2011-04-27" gender="M" nation="BRA" license="405717" swrid="5664737" athleteid="1858" externalid="405717">
              <RESULTS>
                <RESULT eventid="1088" status="DSQ" swimtime="00:03:46.25" resultid="1859" heatid="4284" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="200" swimtime="00:01:20.04" resultid="1860" heatid="4331" lane="5" />
                <RESULT eventid="1220" points="147" swimtime="00:01:47.62" resultid="1861" heatid="4387" lane="1" />
                <RESULT eventid="1306" points="167" swimtime="00:00:42.69" resultid="1862" heatid="4478" lane="1" />
                <RESULT eventid="1374" points="180" swimtime="00:01:31.26" resultid="1863" heatid="4525" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Geórgia" lastname="Adeli Jesus" birthdate="2008-03-27" gender="F" nation="BRA" license="312649" swrid="5596864" athleteid="1830" externalid="312649">
              <RESULTS>
                <RESULT eventid="1116" points="351" swimtime="00:21:44.66" resultid="1831" heatid="4309" lane="1" entrytime="00:21:35.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.83" />
                    <SPLIT distance="200" swimtime="00:02:39.14" />
                    <SPLIT distance="300" swimtime="00:04:03.73" />
                    <SPLIT distance="400" swimtime="00:05:30.81" />
                    <SPLIT distance="500" swimtime="00:06:59.99" />
                    <SPLIT distance="600" swimtime="00:08:29.39" />
                    <SPLIT distance="700" swimtime="00:09:56.52" />
                    <SPLIT distance="800" swimtime="00:11:25.29" />
                    <SPLIT distance="900" swimtime="00:12:54.01" />
                    <SPLIT distance="1000" swimtime="00:14:22.97" />
                    <SPLIT distance="1100" swimtime="00:15:52.37" />
                    <SPLIT distance="1200" swimtime="00:17:23.22" />
                    <SPLIT distance="1300" swimtime="00:18:52.99" />
                    <SPLIT distance="1400" swimtime="00:20:20.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="398" swimtime="00:01:10.24" resultid="1832" heatid="4319" lane="3" />
                <RESULT eventid="1250" points="352" swimtime="00:11:26.01" resultid="1833" heatid="4426" lane="5" entrytime="00:11:17.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.27" />
                    <SPLIT distance="200" swimtime="00:02:39.07" />
                    <SPLIT distance="300" swimtime="00:04:06.62" />
                    <SPLIT distance="400" swimtime="00:05:34.72" />
                    <SPLIT distance="500" swimtime="00:07:03.79" />
                    <SPLIT distance="600" swimtime="00:08:32.57" />
                    <SPLIT distance="700" swimtime="00:10:00.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="380" swimtime="00:02:35.68" resultid="1834" heatid="4454" lane="5" entrytime="00:02:31.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="377" swimtime="00:05:25.57" resultid="1835" heatid="4508" lane="3" entrytime="00:05:28.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.39" />
                    <SPLIT distance="200" swimtime="00:02:36.46" />
                    <SPLIT distance="300" swimtime="00:04:02.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Franco" birthdate="2010-06-09" gender="F" nation="BRA" license="383849" swrid="5596896" athleteid="1813" externalid="383849">
              <RESULTS>
                <RESULT eventid="1096" points="299" swimtime="00:00:36.53" resultid="1814" heatid="4293" lane="7" entrytime="00:00:36.75" entrycourse="LCM" />
                <RESULT eventid="1148" points="367" swimtime="00:01:12.19" resultid="1815" heatid="4323" lane="4" entrytime="00:01:13.61" entrycourse="LCM" />
                <RESULT eventid="1228" points="363" swimtime="00:00:33.08" resultid="1816" heatid="4399" lane="3" entrytime="00:00:33.93" entrycourse="LCM" />
                <RESULT eventid="1282" points="348" swimtime="00:02:40.39" resultid="1817" heatid="4452" lane="4" entrytime="00:02:40.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="321" swimtime="00:05:43.49" resultid="1818" heatid="4507" lane="3" entrytime="00:05:46.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.32" />
                    <SPLIT distance="200" swimtime="00:02:46.94" />
                    <SPLIT distance="300" swimtime="00:04:17.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Xavier" birthdate="2011-10-14" gender="M" nation="BRA" license="370564" swrid="5596949" athleteid="1841" externalid="370564">
              <RESULTS>
                <RESULT eventid="1088" points="218" swimtime="00:03:28.20" resultid="1842" heatid="4283" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="165" swimtime="00:01:25.41" resultid="1843" heatid="4332" lane="5" />
                <RESULT eventid="1220" points="200" swimtime="00:01:37.15" resultid="1844" heatid="4387" lane="3" entrytime="00:01:41.93" entrycourse="LCM" />
                <RESULT eventid="1236" points="171" swimtime="00:00:37.63" resultid="1845" heatid="4410" lane="1" />
                <RESULT eventid="1290" points="182" swimtime="00:02:59.69" resultid="1846" heatid="4459" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Mussi" birthdate="2006-12-31" gender="M" nation="BRA" license="370567" swrid="5596917" athleteid="1847" externalid="370567">
              <RESULTS>
                <RESULT eventid="1104" points="424" swimtime="00:00:29.63" resultid="1848" heatid="4300" lane="5" entrytime="00:00:30.35" entrycourse="LCM" />
                <RESULT eventid="1188" points="465" swimtime="00:00:33.49" resultid="1849" heatid="4368" lane="8" entrytime="00:00:33.86" entrycourse="LCM" />
                <RESULT eventid="1220" points="394" swimtime="00:01:17.57" resultid="1850" heatid="4391" lane="5" entrytime="00:01:20.71" entrycourse="LCM" />
                <RESULT eventid="1306" points="336" swimtime="00:00:33.87" resultid="1851" heatid="4479" lane="4" entrytime="00:00:33.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yago" lastname="Simon Pires" birthdate="2008-10-29" gender="M" nation="BRA" license="328942" swrid="5596939" athleteid="1836" externalid="328942">
              <RESULTS>
                <RESULT eventid="1156" points="510" swimtime="00:00:58.65" resultid="1837" heatid="4341" lane="5" entrytime="00:01:04.47" entrycourse="LCM" />
                <RESULT eventid="1188" points="387" swimtime="00:00:35.59" resultid="1838" heatid="4366" lane="3" entrytime="00:00:36.25" entrycourse="LCM" />
                <RESULT eventid="1236" points="474" swimtime="00:00:26.80" resultid="1839" heatid="4416" lane="8" entrytime="00:00:28.51" entrycourse="LCM" />
                <RESULT eventid="1290" points="432" swimtime="00:02:14.86" resultid="1840" heatid="4464" lane="1" entrytime="00:02:24.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Afonso Proteti" birthdate="2002-03-19" gender="M" nation="BRA" license="190464" swrid="5596865" athleteid="1819" externalid="190464">
              <RESULTS>
                <RESULT eventid="1104" points="690" swimtime="00:00:25.19" resultid="1820" heatid="4304" lane="3" entrytime="00:00:25.51" entrycourse="LCM" />
                <RESULT eventid="1156" points="590" swimtime="00:00:55.86" resultid="1821" heatid="4333" lane="2" />
                <RESULT eventid="1306" points="536" swimtime="00:00:28.98" resultid="1822" heatid="4482" lane="6" entrytime="00:00:28.76" entrycourse="LCM" />
                <RESULT eventid="1342" points="634" swimtime="00:00:57.54" resultid="1823" heatid="4505" lane="5" entrytime="00:00:57.08" entrycourse="LCM" />
                <RESULT eventid="1374" points="567" swimtime="00:01:02.33" resultid="1824" heatid="4533" lane="3" entrytime="00:01:01.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Wirtti" birthdate="2011-01-14" gender="M" nation="BRA" license="383854" swrid="4917570" athleteid="1852" externalid="383854">
              <RESULTS>
                <RESULT eventid="1104" points="239" swimtime="00:00:35.88" resultid="1853" heatid="4298" lane="8" entrytime="00:00:43.02" entrycourse="LCM" />
                <RESULT eventid="1156" points="304" swimtime="00:01:09.68" resultid="1854" heatid="4333" lane="4" />
                <RESULT eventid="1236" points="302" swimtime="00:00:31.16" resultid="1855" heatid="4411" lane="4" entrytime="00:00:33.45" entrycourse="LCM" />
                <RESULT eventid="1306" points="286" swimtime="00:00:35.71" resultid="1856" heatid="4478" lane="4" entrytime="00:00:39.69" entrycourse="LCM" />
                <RESULT eventid="1374" points="221" swimtime="00:01:25.34" resultid="1857" heatid="4526" lane="3" entrytime="00:01:32.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13025" nation="BRA" region="PR" clubid="2042" swrid="93779" name="Instituto Desportos Aquáticos De Foz Do Iguaçu" shortname="Cataratas Natação">
          <ATHLETES>
            <ATHLETE firstname="Vinicius" lastname="Monteiro Viebrantz" birthdate="2003-01-09" gender="M" nation="BRA" license="291175" swrid="5600219" athleteid="2053" externalid="291175">
              <RESULTS>
                <RESULT eventid="1236" points="614" swimtime="00:00:24.59" resultid="2054" heatid="4422" lane="3" entrytime="00:00:23.44" entrycourse="LCM" />
                <RESULT eventid="1306" points="474" swimtime="00:00:30.20" resultid="2055" heatid="4478" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="De Souza Tulio" birthdate="2006-06-23" gender="F" nation="BRA" license="342344" swrid="5030980" athleteid="2068" externalid="342344">
              <RESULTS>
                <RESULT eventid="1064" points="533" swimtime="00:02:31.80" resultid="2069" heatid="4271" lane="5" entrytime="00:02:31.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="584" swimtime="00:01:01.84" resultid="2070" heatid="4330" lane="4" entrytime="00:01:00.16" entrycourse="LCM" />
                <RESULT eventid="1228" points="569" swimtime="00:00:28.49" resultid="2071" heatid="4405" lane="5" entrytime="00:00:27.80" entrycourse="LCM" />
                <RESULT eventid="1282" status="DNS" swimtime="00:00:00.00" resultid="2072" heatid="4457" lane="3" entrytime="00:02:10.02" entrycourse="LCM" />
                <RESULT eventid="1366" status="DNS" swimtime="00:00:00.00" resultid="2073" heatid="4524" lane="5" entrytime="00:01:08.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Axel" lastname="Ariel Giménez González" birthdate="2011-06-01" gender="M" nation="BRA" license="365755" swrid="5676299" athleteid="2170" externalid="365755">
              <RESULTS>
                <RESULT eventid="1156" points="372" swimtime="00:01:05.15" resultid="2171" heatid="4333" lane="8" />
                <RESULT eventid="1188" points="296" swimtime="00:00:38.90" resultid="2172" heatid="4362" lane="3" />
                <RESULT eventid="1236" points="346" swimtime="00:00:29.77" resultid="2173" heatid="4410" lane="8" />
                <RESULT eventid="1290" points="281" swimtime="00:02:35.71" resultid="2174" heatid="4459" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="259" swimtime="00:01:20.88" resultid="2175" heatid="4525" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Christopher" lastname="De Araujo" birthdate="2008-08-09" gender="M" nation="BRA" license="366376" swrid="5596884" athleteid="2098" externalid="366376">
              <RESULTS>
                <RESULT eventid="1088" points="435" swimtime="00:02:45.59" resultid="2099" heatid="4288" lane="6" entrytime="00:02:41.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="428" swimtime="00:05:21.77" resultid="2100" heatid="4318" lane="8" entrytime="00:05:15.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.94" />
                    <SPLIT distance="200" swimtime="00:02:40.24" />
                    <SPLIT distance="300" swimtime="00:04:11.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="440" swimtime="00:01:14.76" resultid="2101" heatid="4394" lane="8" entrytime="00:01:12.24" entrycourse="LCM" />
                <RESULT eventid="1290" points="488" swimtime="00:02:09.54" resultid="2102" heatid="4468" lane="8" entrytime="00:02:05.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="521" swimtime="00:04:33.48" resultid="2103" heatid="4511" lane="4" entrytime="00:05:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.29" />
                    <SPLIT distance="200" swimtime="00:02:13.44" />
                    <SPLIT distance="300" swimtime="00:03:24.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Resende Ames" birthdate="2006-02-10" gender="M" nation="BRA" license="365657" swrid="5596931" athleteid="2080" externalid="365657">
              <RESULTS>
                <RESULT eventid="1072" points="464" swimtime="00:02:24.51" resultid="2081" heatid="4273" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="524" swimtime="00:02:16.78" resultid="2082" heatid="4354" lane="6" entrytime="00:02:16.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="528" swimtime="00:00:25.86" resultid="2083" heatid="4420" lane="2" entrytime="00:00:25.59" entrycourse="LCM" />
                <RESULT eventid="1290" points="550" swimtime="00:02:04.43" resultid="2084" heatid="4468" lane="7" entrytime="00:02:04.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="575" swimtime="00:00:59.44" resultid="2085" heatid="4505" lane="2" entrytime="00:00:59.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Targat Pinheiro" birthdate="2008-09-04" gender="F" nation="BRA" license="331610" swrid="5596894" athleteid="2043" externalid="331610">
              <RESULTS>
                <RESULT eventid="1064" points="396" swimtime="00:02:47.67" resultid="2044" heatid="4267" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="441" swimtime="00:05:49.21" resultid="2045" heatid="4315" lane="6" entrytime="00:05:44.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.13" />
                    <SPLIT distance="200" swimtime="00:02:45.50" />
                    <SPLIT distance="300" swimtime="00:04:29.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="442" swimtime="00:10:35.98" resultid="2046" heatid="4427" lane="4" entrytime="00:10:36.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.38" />
                    <SPLIT distance="200" swimtime="00:02:31.81" />
                    <SPLIT distance="300" swimtime="00:03:51.88" />
                    <SPLIT distance="400" swimtime="00:05:12.96" />
                    <SPLIT distance="500" swimtime="00:06:34.19" />
                    <SPLIT distance="600" swimtime="00:07:57.25" />
                    <SPLIT distance="700" swimtime="00:09:19.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="441" swimtime="00:01:12.87" resultid="2047" heatid="4497" lane="1" entrytime="00:01:12.83" entrycourse="LCM" />
                <RESULT eventid="1366" points="386" swimtime="00:01:18.73" resultid="2048" heatid="4523" lane="1" entrytime="00:01:17.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Mattiello" birthdate="2009-04-11" gender="F" nation="BRA" license="367011" swrid="5596914" athleteid="2110" externalid="367011">
              <RESULTS>
                <RESULT eventid="1148" points="433" swimtime="00:01:08.35" resultid="2111" heatid="4325" lane="3" entrytime="00:01:10.76" entrycourse="LCM" />
                <RESULT eventid="1228" points="431" swimtime="00:00:31.25" resultid="2112" heatid="4401" lane="4" entrytime="00:00:31.90" entrycourse="LCM" />
                <RESULT eventid="1282" points="393" swimtime="00:02:33.94" resultid="2113" heatid="4453" lane="2" entrytime="00:02:35.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="312" swimtime="00:01:24.47" resultid="2114" heatid="4520" lane="8" entrytime="00:01:28.28" entrycourse="LCM" />
                <RESULT eventid="1350" points="372" swimtime="00:05:26.99" resultid="2115" heatid="4508" lane="1" entrytime="00:05:36.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.44" />
                    <SPLIT distance="200" swimtime="00:02:42.77" />
                    <SPLIT distance="300" swimtime="00:04:07.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Luiz Martinazzo" birthdate="2006-05-16" gender="M" nation="BRA" license="345593" swrid="5596910" athleteid="2092" externalid="345593">
              <RESULTS>
                <RESULT eventid="1072" points="385" swimtime="00:02:33.82" resultid="2093" heatid="4276" lane="1" entrytime="00:02:30.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="546" swimtime="00:00:57.33" resultid="2094" heatid="4345" lane="6" entrytime="00:00:59.14" entrycourse="LCM" />
                <RESULT eventid="1258" points="466" swimtime="00:18:43.29" resultid="2095" heatid="4430" lane="4" entrytime="00:21:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.20" />
                    <SPLIT distance="200" swimtime="00:02:17.20" />
                    <SPLIT distance="300" swimtime="00:03:29.64" />
                    <SPLIT distance="400" swimtime="00:04:43.71" />
                    <SPLIT distance="500" swimtime="00:06:00.70" />
                    <SPLIT distance="600" swimtime="00:07:18.55" />
                    <SPLIT distance="700" swimtime="00:08:35.81" />
                    <SPLIT distance="800" swimtime="00:09:52.20" />
                    <SPLIT distance="900" swimtime="00:11:08.91" />
                    <SPLIT distance="1000" swimtime="00:12:25.57" />
                    <SPLIT distance="1100" swimtime="00:13:42.72" />
                    <SPLIT distance="1200" swimtime="00:14:59.23" />
                    <SPLIT distance="1300" swimtime="00:16:15.98" />
                    <SPLIT distance="1400" swimtime="00:17:30.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="487" swimtime="00:02:09.60" resultid="2096" heatid="4467" lane="4" entrytime="00:02:06.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="440" swimtime="00:01:07.83" resultid="2097" heatid="4532" lane="7" entrytime="00:01:06.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Marques Petry" birthdate="2008-01-08" gender="M" nation="BRA" license="392351" swrid="4711489" athleteid="2122" externalid="392351">
              <RESULTS>
                <RESULT eventid="1124" points="367" swimtime="00:10:30.92" resultid="2123" heatid="4310" lane="2" entrytime="00:11:24.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.95" />
                    <SPLIT distance="200" swimtime="00:02:29.66" />
                    <SPLIT distance="300" swimtime="00:03:51.25" />
                    <SPLIT distance="400" swimtime="00:05:11.79" />
                    <SPLIT distance="500" swimtime="00:06:32.70" />
                    <SPLIT distance="600" swimtime="00:07:53.68" />
                    <SPLIT distance="700" swimtime="00:09:15.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="385" swimtime="00:01:04.38" resultid="2124" heatid="4337" lane="5" entrytime="00:01:09.36" entrycourse="LCM" />
                <RESULT eventid="1258" points="384" swimtime="00:19:57.47" resultid="2125" heatid="4431" lane="8" entrytime="00:21:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.07" />
                    <SPLIT distance="200" swimtime="00:02:32.09" />
                    <SPLIT distance="300" swimtime="00:03:52.36" />
                    <SPLIT distance="400" swimtime="00:05:13.13" />
                    <SPLIT distance="500" swimtime="00:06:33.96" />
                    <SPLIT distance="600" swimtime="00:07:54.68" />
                    <SPLIT distance="700" swimtime="00:09:14.62" />
                    <SPLIT distance="800" swimtime="00:10:34.90" />
                    <SPLIT distance="900" swimtime="00:11:54.35" />
                    <SPLIT distance="1000" swimtime="00:13:13.68" />
                    <SPLIT distance="1100" swimtime="00:14:34.31" />
                    <SPLIT distance="1200" swimtime="00:15:55.60" />
                    <SPLIT distance="1300" swimtime="00:17:16.84" />
                    <SPLIT distance="1400" swimtime="00:18:39.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="385" swimtime="00:02:20.21" resultid="2126" heatid="4462" lane="1" entrytime="00:02:34.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="378" swimtime="00:05:04.35" resultid="2127" heatid="4512" lane="2" entrytime="00:05:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.95" />
                    <SPLIT distance="200" swimtime="00:02:26.53" />
                    <SPLIT distance="300" swimtime="00:03:45.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ysadora" lastname="Bertoldo" birthdate="2010-04-09" gender="F" nation="BRA" license="376444" swrid="5588553" athleteid="2134" externalid="376444">
              <RESULTS>
                <RESULT eventid="1116" points="433" swimtime="00:20:16.26" resultid="2135" heatid="4309" lane="8" entrytime="00:22:39.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.84" />
                    <SPLIT distance="200" swimtime="00:02:37.20" />
                    <SPLIT distance="300" swimtime="00:03:58.11" />
                    <SPLIT distance="400" swimtime="00:05:20.03" />
                    <SPLIT distance="500" swimtime="00:06:42.26" />
                    <SPLIT distance="600" swimtime="00:08:03.04" />
                    <SPLIT distance="700" swimtime="00:09:25.05" />
                    <SPLIT distance="800" swimtime="00:10:46.84" />
                    <SPLIT distance="900" swimtime="00:12:08.13" />
                    <SPLIT distance="1000" swimtime="00:13:29.90" />
                    <SPLIT distance="1100" swimtime="00:14:51.93" />
                    <SPLIT distance="1200" swimtime="00:16:14.52" />
                    <SPLIT distance="1300" swimtime="00:17:36.18" />
                    <SPLIT distance="1400" swimtime="00:18:58.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="391" swimtime="00:01:10.68" resultid="2136" heatid="4322" lane="2" entrytime="00:01:19.05" entrycourse="LCM" />
                <RESULT eventid="1250" points="432" swimtime="00:10:41.22" resultid="2137" heatid="4426" lane="2" entrytime="00:11:45.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.43" />
                    <SPLIT distance="200" swimtime="00:02:35.23" />
                    <SPLIT distance="300" swimtime="00:03:56.63" />
                    <SPLIT distance="400" swimtime="00:05:18.08" />
                    <SPLIT distance="500" swimtime="00:06:39.96" />
                    <SPLIT distance="600" swimtime="00:08:01.53" />
                    <SPLIT distance="700" swimtime="00:09:22.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="412" swimtime="00:02:31.65" resultid="2138" heatid="4452" lane="2" entrytime="00:02:46.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="425" swimtime="00:05:13.03" resultid="2139" heatid="4507" lane="4" entrytime="00:05:41.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.29" />
                    <SPLIT distance="200" swimtime="00:02:34.55" />
                    <SPLIT distance="300" swimtime="00:03:55.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Rogge" birthdate="2008-09-02" gender="M" nation="BRA" license="383387" swrid="4883279" athleteid="2062" externalid="383387">
              <RESULTS>
                <RESULT eventid="1156" points="507" swimtime="00:00:58.75" resultid="2063" heatid="4343" lane="5" entrytime="00:01:00.59" entrycourse="LCM" />
                <RESULT eventid="1236" points="490" swimtime="00:00:26.52" resultid="2064" heatid="4418" lane="4" entrytime="00:00:26.82" entrycourse="LCM" />
                <RESULT eventid="1290" points="323" swimtime="00:02:28.56" resultid="2065" heatid="4459" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1306" points="406" swimtime="00:00:31.79" resultid="2066" heatid="4481" lane="8" entrytime="00:00:31.79" entrycourse="LCM" />
                <RESULT eventid="1374" points="338" swimtime="00:01:14.05" resultid="2067" heatid="4529" lane="3" entrytime="00:01:12.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Faisal" lastname="Basem Ghotme" birthdate="2010-12-18" gender="M" nation="BRA" license="390809" swrid="5596871" athleteid="2152" externalid="390809">
              <RESULTS>
                <RESULT eventid="1072" points="378" swimtime="00:02:34.72" resultid="2153" heatid="4274" lane="5" entrytime="00:02:40.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="399" swimtime="00:01:03.62" resultid="2154" heatid="4339" lane="4" entrytime="00:01:06.60" entrycourse="LCM" />
                <RESULT eventid="1236" points="431" swimtime="00:00:27.68" resultid="2155" heatid="4414" lane="4" entrytime="00:00:29.94" entrycourse="LCM" />
                <RESULT eventid="1290" status="DNS" swimtime="00:00:00.00" resultid="2156" heatid="4461" lane="3" entrytime="00:02:37.79" entrycourse="LCM" />
                <RESULT eventid="1374" status="DNS" swimtime="00:00:00.00" resultid="2157" heatid="4530" lane="8" entrytime="00:01:12.05" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Gabriel Dreher" birthdate="2011-12-05" gender="M" nation="BRA" license="403148" swrid="5676302" athleteid="2164" externalid="403148">
              <RESULTS>
                <RESULT eventid="1156" points="147" swimtime="00:01:28.67" resultid="2165" heatid="4333" lane="3" />
                <RESULT eventid="1188" points="116" swimtime="00:00:53.11" resultid="2166" heatid="4361" lane="8" />
                <RESULT eventid="1236" points="169" swimtime="00:00:37.75" resultid="2167" heatid="4408" lane="7" />
                <RESULT eventid="1306" points="124" swimtime="00:00:47.17" resultid="2168" heatid="4477" lane="1" />
                <RESULT eventid="1374" points="112" swimtime="00:01:46.83" resultid="2169" heatid="4526" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Oliveira" birthdate="2003-07-16" gender="M" nation="BRA" license="295723" swrid="5596944" athleteid="2074" externalid="295723">
              <RESULTS>
                <RESULT eventid="1072" points="483" swimtime="00:02:22.59" resultid="2075" heatid="4276" lane="5" entrytime="00:02:20.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="504" swimtime="00:00:26.26" resultid="2076" heatid="4418" lane="1" entrytime="00:00:27.05" entrycourse="LCM" />
                <RESULT eventid="1306" points="479" swimtime="00:00:30.08" resultid="2077" heatid="4482" lane="2" entrytime="00:00:28.82" entrycourse="LCM" />
                <RESULT eventid="1342" points="519" swimtime="00:01:01.50" resultid="2078" heatid="4505" lane="7" entrytime="00:00:59.84" entrycourse="LCM" />
                <RESULT eventid="1374" points="484" swimtime="00:01:05.71" resultid="2079" heatid="4532" lane="4" entrytime="00:01:02.33" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="De Assis Santos" birthdate="2003-02-21" gender="M" nation="BRA" license="342496" swrid="5596885" athleteid="2086" externalid="342496">
              <RESULTS>
                <RESULT eventid="1072" points="414" swimtime="00:02:30.06" resultid="2087" heatid="4276" lane="7" entrytime="00:02:28.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" status="DSQ" swimtime="00:05:41.90" resultid="2088" heatid="4317" lane="7" entrytime="00:05:46.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.29" />
                    <SPLIT distance="200" swimtime="00:02:41.54" />
                    <SPLIT distance="300" swimtime="00:04:22.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1306" points="438" swimtime="00:00:31.00" resultid="2089" heatid="4481" lane="6" entrytime="00:00:31.01" entrycourse="LCM" />
                <RESULT eventid="1274" points="385" swimtime="00:02:36.59" resultid="2090" heatid="4445" lane="5" entrytime="00:02:39.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="447" swimtime="00:01:07.46" resultid="2091" heatid="4532" lane="2" entrytime="00:01:05.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabrizzio" lastname="Paolo Cazzola" birthdate="2009-06-15" gender="M" nation="BRA" license="357168" swrid="5596922" athleteid="2116" externalid="357168">
              <RESULTS>
                <RESULT eventid="1072" points="319" swimtime="00:02:43.77" resultid="2117" heatid="4274" lane="6" entrytime="00:02:44.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="388" swimtime="00:01:04.20" resultid="2118" heatid="4332" lane="3" />
                <RESULT eventid="1306" points="315" swimtime="00:00:34.59" resultid="2119" heatid="4477" lane="3" />
                <RESULT eventid="1274" points="323" swimtime="00:02:46.02" resultid="2120" heatid="4444" lane="3" entrytime="00:02:52.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="314" swimtime="00:01:15.85" resultid="2121" heatid="4528" lane="3" entrytime="00:01:16.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Bailke" birthdate="2007-05-04" gender="M" nation="BRA" license="370566" swrid="5596869" athleteid="2104" externalid="370566">
              <RESULTS>
                <RESULT eventid="1124" points="345" swimtime="00:10:44.50" resultid="2105" heatid="4310" lane="1" entrytime="00:11:24.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.78" />
                    <SPLIT distance="200" swimtime="00:02:33.73" />
                    <SPLIT distance="300" swimtime="00:03:55.68" />
                    <SPLIT distance="400" swimtime="00:05:17.39" />
                    <SPLIT distance="500" swimtime="00:06:42.76" />
                    <SPLIT distance="600" swimtime="00:08:03.57" />
                    <SPLIT distance="700" swimtime="00:09:26.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="218" swimtime="00:03:03.32" resultid="2106" heatid="4352" lane="3" entrytime="00:02:54.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="353" swimtime="00:20:31.34" resultid="2107" heatid="4430" lane="7" entrytime="00:21:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.10" />
                    <SPLIT distance="200" swimtime="00:02:37.42" />
                    <SPLIT distance="300" swimtime="00:04:00.13" />
                    <SPLIT distance="400" swimtime="00:05:23.91" />
                    <SPLIT distance="500" swimtime="00:06:47.65" />
                    <SPLIT distance="600" swimtime="00:08:09.91" />
                    <SPLIT distance="700" swimtime="00:09:32.51" />
                    <SPLIT distance="800" swimtime="00:10:52.85" />
                    <SPLIT distance="900" swimtime="00:12:16.11" />
                    <SPLIT distance="1000" swimtime="00:13:40.51" />
                    <SPLIT distance="1100" swimtime="00:15:02.13" />
                    <SPLIT distance="1200" swimtime="00:16:25.79" />
                    <SPLIT distance="1300" swimtime="00:17:48.31" />
                    <SPLIT distance="1400" swimtime="00:19:10.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="387" swimtime="00:02:19.90" resultid="2108" heatid="4465" lane="1" entrytime="00:02:19.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="303" swimtime="00:01:13.61" resultid="2109" heatid="4501" lane="5" entrytime="00:01:13.22" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mayumi" lastname="Napole" birthdate="2010-02-01" gender="F" nation="BRA" license="376446" swrid="5596918" athleteid="2146" externalid="376446">
              <RESULTS>
                <RESULT eventid="1080" points="266" swimtime="00:03:33.68" resultid="2147" heatid="4280" lane="8" entrytime="00:03:19.92" entrycourse="LCM" />
                <RESULT eventid="1148" points="411" swimtime="00:01:09.51" resultid="2148" heatid="4324" lane="4" entrytime="00:01:11.78" entrycourse="LCM" />
                <RESULT eventid="1228" points="413" swimtime="00:00:31.70" resultid="2149" heatid="4400" lane="1" entrytime="00:00:33.15" entrycourse="LCM" />
                <RESULT eventid="1266" points="302" swimtime="00:03:07.90" resultid="2150" heatid="4435" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="335" swimtime="00:01:22.49" resultid="2151" heatid="4521" lane="1" entrytime="00:01:23.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Marques Petry" birthdate="2008-01-08" gender="M" nation="BRA" license="392352" swrid="4795316" athleteid="2128" externalid="392352">
              <RESULTS>
                <RESULT eventid="1088" points="260" swimtime="00:03:16.51" resultid="2129" heatid="4283" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="412" swimtime="00:01:02.95" resultid="2130" heatid="4340" lane="4" entrytime="00:01:05.68" entrycourse="LCM" />
                <RESULT eventid="1220" points="253" swimtime="00:01:29.89" resultid="2131" heatid="4389" lane="6" entrytime="00:01:30.83" entrycourse="LCM" />
                <RESULT eventid="1290" points="369" swimtime="00:02:22.13" resultid="2132" heatid="4459" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="298" swimtime="00:01:17.20" resultid="2133" heatid="4528" lane="8" entrytime="00:01:19.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Sermidi" birthdate="2005-06-15" gender="F" nation="BRA" license="283035" swrid="5596938" athleteid="2049" externalid="283035">
              <RESULTS>
                <RESULT eventid="1228" points="480" swimtime="00:00:30.14" resultid="2050" heatid="4403" lane="6" entrytime="00:00:30.56" entrycourse="LCM" />
                <RESULT eventid="1298" points="391" swimtime="00:00:36.71" resultid="2051" heatid="4475" lane="7" entrytime="00:00:35.27" entrycourse="LCM" />
                <RESULT eventid="1366" points="384" swimtime="00:01:18.82" resultid="2052" heatid="4523" lane="8" entrytime="00:01:18.42" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Leticia Sbardelatti" birthdate="2011-07-28" gender="F" nation="BRA" license="403147" swrid="5676303" athleteid="2158" externalid="403147">
              <RESULTS>
                <RESULT eventid="1148" points="217" swimtime="00:01:26.04" resultid="2159" heatid="4319" lane="2" />
                <RESULT eventid="1180" points="185" swimtime="00:00:51.16" resultid="2160" heatid="4355" lane="1" />
                <RESULT eventid="1228" points="253" swimtime="00:00:37.32" resultid="2161" heatid="4397" lane="1" />
                <RESULT eventid="1282" points="188" swimtime="00:03:16.81" resultid="2162" heatid="4450" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="125" swimtime="00:00:53.60" resultid="2163" heatid="4471" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Resende Ames" birthdate="2010-02-02" gender="M" nation="BRA" license="365505" swrid="5588876" athleteid="2140" externalid="365505">
              <RESULTS>
                <RESULT eventid="1072" points="427" swimtime="00:02:28.55" resultid="2141" heatid="4276" lane="3" entrytime="00:02:25.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="426" swimtime="00:01:02.23" resultid="2142" heatid="4338" lane="6" entrytime="00:01:07.83" entrycourse="LCM" />
                <RESULT eventid="1236" points="388" swimtime="00:00:28.66" resultid="2143" heatid="4408" lane="1" />
                <RESULT eventid="1306" points="406" swimtime="00:00:31.79" resultid="2144" heatid="4480" lane="2" entrytime="00:00:32.87" entrycourse="LCM" />
                <RESULT eventid="1374" points="434" swimtime="00:01:08.15" resultid="2145" heatid="4532" lane="8" entrytime="00:01:07.32" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Carolina Ghellere" birthdate="2007-06-05" gender="F" nation="BRA" license="312662" swrid="5596874" athleteid="2056" externalid="312662">
              <RESULTS>
                <RESULT eventid="1096" points="507" swimtime="00:00:30.62" resultid="2057" heatid="4294" lane="4" entrytime="00:00:29.29" entrycourse="LCM" />
                <RESULT eventid="1148" points="547" swimtime="00:01:03.22" resultid="2058" heatid="4330" lane="3" entrytime="00:01:00.70" entrycourse="LCM" />
                <RESULT eventid="1282" points="578" swimtime="00:02:15.46" resultid="2059" heatid="4457" lane="5" entrytime="00:02:07.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="529" swimtime="00:01:08.57" resultid="2060" heatid="4497" lane="4" entrytime="00:01:03.53" entrycourse="LCM" />
                <RESULT eventid="1350" points="538" swimtime="00:04:49.25" resultid="2061" heatid="4510" lane="5" entrytime="00:04:25.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.80" />
                    <SPLIT distance="200" swimtime="00:02:21.04" />
                    <SPLIT distance="300" swimtime="00:03:35.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="16" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1206" points="400" swimtime="00:09:27.89" resultid="2176" heatid="4374" lane="6" entrytime="00:09:11.79">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.88" />
                    <SPLIT distance="200" swimtime="00:02:07.56" />
                    <SPLIT distance="300" swimtime="00:03:18.16" />
                    <SPLIT distance="400" swimtime="00:04:37.34" />
                    <SPLIT distance="500" swimtime="00:05:51.06" />
                    <SPLIT distance="600" swimtime="00:07:07.97" />
                    <SPLIT distance="700" swimtime="00:08:14.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2098" number="1" />
                    <RELAYPOSITION athleteid="2062" number="2" />
                    <RELAYPOSITION athleteid="2128" number="3" />
                    <RELAYPOSITION athleteid="2122" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1326" status="WDR" swimtime="00:00:00.00" resultid="2177" heatid="4489" lane="2" entrytime="00:05:13.43" />
                <RESULT eventid="1394" status="WDR" swimtime="00:00:00.00" resultid="2180" heatid="4540" lane="6" entrytime="00:04:44.02" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1330" status="DSQ" swimtime="00:05:03.66" resultid="2178" heatid="4491" lane="3" entrytime="00:05:15.22">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.25" />
                    <SPLIT distance="200" swimtime="00:02:53.74" />
                    <SPLIT distance="300" swimtime="00:04:03.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2122" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2128" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="2098" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="2062" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1398" points="455" swimtime="00:04:04.70" resultid="2182" heatid="4542" lane="5" entrytime="00:04:16.87">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.26" />
                    <SPLIT distance="200" swimtime="00:01:57.68" />
                    <SPLIT distance="300" swimtime="00:03:02.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2062" number="1" />
                    <RELAYPOSITION athleteid="2098" number="2" />
                    <RELAYPOSITION athleteid="2122" number="3" />
                    <RELAYPOSITION athleteid="2128" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1332" points="472" swimtime="00:04:25.46" resultid="2179" heatid="4492" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.07" />
                    <SPLIT distance="300" swimtime="00:03:31.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2074" number="1" />
                    <RELAYPOSITION athleteid="2086" number="2" />
                    <RELAYPOSITION athleteid="2080" number="3" />
                    <RELAYPOSITION athleteid="2053" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1400" points="527" swimtime="00:03:52.98" resultid="2181" heatid="4543" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.59" />
                    <SPLIT distance="200" swimtime="00:01:58.03" />
                    <SPLIT distance="300" swimtime="00:02:54.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2080" number="1" />
                    <RELAYPOSITION athleteid="2086" number="2" />
                    <RELAYPOSITION athleteid="2092" number="3" />
                    <RELAYPOSITION athleteid="2074" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1114" status="DSQ" swimtime="00:05:08.79" resultid="2183" heatid="4307" lane="7" entrytime="00:05:26.20">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.25" />
                    <SPLIT distance="300" swimtime="00:03:59.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2152" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2146" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="2140" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="2134" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1248" points="518" swimtime="00:04:30.77" resultid="2184" heatid="4425" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.84" />
                    <SPLIT distance="200" swimtime="00:02:30.79" />
                    <SPLIT distance="300" swimtime="00:03:29.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2074" number="1" />
                    <RELAYPOSITION athleteid="2056" number="2" />
                    <RELAYPOSITION athleteid="2080" number="3" />
                    <RELAYPOSITION athleteid="2068" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1246" points="421" swimtime="00:04:50.27" resultid="2185" heatid="4424" lane="3" entrytime="00:04:42.42">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.42" />
                    <SPLIT distance="200" swimtime="00:02:27.83" />
                    <SPLIT distance="300" swimtime="00:03:41.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2062" number="1" />
                    <RELAYPOSITION athleteid="2098" number="2" />
                    <RELAYPOSITION athleteid="2043" number="3" />
                    <RELAYPOSITION athleteid="2110" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="1007" nation="BRA" region="PR" clubid="3480" swrid="93785" name="Santa Mônica Clube De Campo" shortname="Santa Mônica">
          <ATHLETES>
            <ATHLETE firstname="Juliana" lastname="Moreira Furtado" birthdate="2011-01-27" gender="F" nation="BRA" license="403783" swrid="5684587" athleteid="3699" externalid="403783">
              <RESULTS>
                <RESULT eventid="1148" points="232" swimtime="00:01:24.08" resultid="3700" heatid="4321" lane="8" entrytime="00:01:27.48" entrycourse="LCM" />
                <RESULT eventid="1228" points="235" swimtime="00:00:38.21" resultid="3701" heatid="4397" lane="3" entrytime="00:00:51.29" entrycourse="LCM" />
                <RESULT eventid="1282" points="240" swimtime="00:03:01.39" resultid="3702" heatid="4450" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="136" swimtime="00:00:52.18" resultid="3703" heatid="4471" lane="5" entrytime="00:01:10.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Cavassin Ieger" birthdate="2011-08-31" gender="M" nation="BRA" license="367149" swrid="5588743" athleteid="3592" externalid="367149">
              <RESULTS>
                <RESULT eventid="1088" points="259" swimtime="00:03:16.64" resultid="3593" heatid="4285" lane="7" entrytime="00:03:16.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="248" swimtime="00:00:41.26" resultid="3594" heatid="4364" lane="6" entrytime="00:00:43.89" entrycourse="LCM" />
                <RESULT eventid="1220" points="247" swimtime="00:01:30.59" resultid="3595" heatid="4388" lane="3" entrytime="00:01:34.32" entrycourse="LCM" />
                <RESULT eventid="1274" points="276" swimtime="00:02:54.94" resultid="3596" heatid="4443" lane="2" entrytime="00:03:04.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="213" swimtime="00:01:22.70" resultid="3597" heatid="4499" lane="4" entrytime="00:01:23.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Analyce" lastname="Nunes Porto Luz" birthdate="2006-10-29" gender="F" nation="BRA" license="369322" swrid="5600226" athleteid="3499" externalid="369322">
              <RESULTS>
                <RESULT eventid="1096" points="457" swimtime="00:00:31.71" resultid="3500" heatid="4294" lane="2" entrytime="00:00:32.01" entrycourse="LCM" />
                <RESULT eventid="1148" points="540" swimtime="00:01:03.48" resultid="3501" heatid="4330" lane="8" entrytime="00:01:03.42" entrycourse="LCM" />
                <RESULT eventid="1282" points="526" swimtime="00:02:19.76" resultid="3502" heatid="4457" lane="1" entrytime="00:02:16.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="421" swimtime="00:01:14.02" resultid="3503" heatid="4497" lane="7" entrytime="00:01:11.70" entrycourse="LCM" />
                <RESULT eventid="1350" points="455" swimtime="00:05:06.03" resultid="3504" heatid="4510" lane="8" entrytime="00:04:50.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.03" />
                    <SPLIT distance="200" swimtime="00:02:26.67" />
                    <SPLIT distance="300" swimtime="00:03:47.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="De Castro Paiva Maciel" birthdate="2008-04-10" gender="M" nation="BRA" license="378333" swrid="5622275" athleteid="3505" externalid="378333">
              <RESULTS>
                <RESULT eventid="1104" points="464" swimtime="00:00:28.75" resultid="3506" heatid="4301" lane="3" entrytime="00:00:29.54" entrycourse="LCM" />
                <RESULT eventid="1156" points="498" swimtime="00:00:59.09" resultid="3507" heatid="4343" lane="2" entrytime="00:01:01.00" entrycourse="LCM" />
                <RESULT eventid="1236" points="470" swimtime="00:00:26.88" resultid="3508" heatid="4416" lane="2" entrytime="00:00:28.07" entrycourse="LCM" />
                <RESULT eventid="1290" points="426" swimtime="00:02:15.54" resultid="3509" heatid="4465" lane="8" entrytime="00:02:20.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="390" swimtime="00:01:07.65" resultid="3510" heatid="4501" lane="3" entrytime="00:01:14.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diego" lastname="Brasil Caropreso" birthdate="2009-10-29" gender="M" nation="BRA" license="399502" swrid="5653287" athleteid="3710" externalid="399502">
              <RESULTS>
                <RESULT eventid="1104" points="347" swimtime="00:00:31.69" resultid="3711" heatid="4298" lane="4" entrytime="00:00:36.07" entrycourse="LCM" />
                <RESULT eventid="1156" points="393" swimtime="00:01:03.94" resultid="3712" heatid="4341" lane="8" entrytime="00:01:05.51" entrycourse="LCM" />
                <RESULT eventid="1236" points="397" swimtime="00:00:28.45" resultid="3713" heatid="4415" lane="3" entrytime="00:00:29.21" entrycourse="LCM" />
                <RESULT eventid="1290" points="309" swimtime="00:02:30.78" resultid="3714" heatid="4463" lane="6" entrytime="00:02:27.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="262" swimtime="00:01:17.20" resultid="3715" heatid="4500" lane="1" entrytime="00:01:18.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathalia" lastname="Lourenco Osorio" birthdate="2007-04-14" gender="F" nation="BRA" license="307465" swrid="5600203" athleteid="3487" externalid="307465">
              <RESULTS>
                <RESULT eventid="1064" points="511" swimtime="00:02:33.97" resultid="3488" heatid="4271" lane="4" entrytime="00:02:29.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="435" swimtime="00:00:38.47" resultid="3489" heatid="4358" lane="5" entrytime="00:00:38.77" entrycourse="LCM" />
                <RESULT eventid="1228" points="540" swimtime="00:00:28.98" resultid="3490" heatid="4405" lane="6" entrytime="00:00:28.10" entrycourse="LCM" />
                <RESULT eventid="1298" points="583" swimtime="00:00:32.14" resultid="3491" heatid="4475" lane="5" entrytime="00:00:31.80" entrycourse="LCM" />
                <RESULT eventid="1366" points="526" swimtime="00:01:10.99" resultid="3492" heatid="4524" lane="3" entrytime="00:01:08.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otto" lastname="Hedeke" birthdate="2011-03-24" gender="M" nation="BRA" license="372643" swrid="5588738" athleteid="3646" externalid="372643">
              <RESULTS>
                <RESULT eventid="1088" points="187" swimtime="00:03:39.22" resultid="3647" heatid="4284" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="129" swimtime="00:03:38.33" resultid="3648" heatid="4351" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="162" swimtime="00:01:44.17" resultid="3649" heatid="4385" lane="3" />
                <RESULT eventid="1290" points="275" swimtime="00:02:36.81" resultid="3650" heatid="4461" lane="2" entrytime="00:02:40.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="144" swimtime="00:01:34.21" resultid="3651" heatid="4498" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Augusto Vaz" birthdate="2011-06-25" gender="M" nation="BRA" license="401737" swrid="5661339" athleteid="3682" externalid="401737">
              <RESULTS>
                <RESULT eventid="1104" points="288" swimtime="00:00:33.69" resultid="3683" heatid="4296" lane="1" />
                <RESULT eventid="1156" points="310" swimtime="00:01:09.18" resultid="3684" heatid="4337" lane="1" entrytime="00:01:11.01" entrycourse="LCM" />
                <RESULT eventid="1236" points="310" swimtime="00:00:30.87" resultid="3685" heatid="4411" lane="2" entrytime="00:00:35.22" entrycourse="LCM" />
                <RESULT eventid="1306" points="235" swimtime="00:00:38.14" resultid="3686" heatid="4478" lane="3" entrytime="00:00:45.56" entrycourse="LCM" />
                <RESULT eventid="1342" points="248" swimtime="00:01:18.70" resultid="3687" heatid="4499" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietra" lastname="Vitoria Paczrowski" birthdate="2009-08-12" gender="F" nation="BRA" license="351253" swrid="5600275" athleteid="3541" externalid="351253">
              <RESULTS>
                <RESULT eventid="1148" points="457" swimtime="00:01:07.11" resultid="3542" heatid="4327" lane="4" entrytime="00:01:07.29" entrycourse="LCM" />
                <RESULT eventid="1228" points="467" swimtime="00:00:30.42" resultid="3543" heatid="4403" lane="5" entrytime="00:00:30.36" entrycourse="LCM" />
                <RESULT eventid="1282" points="433" swimtime="00:02:29.06" resultid="3544" heatid="4455" lane="6" entrytime="00:02:27.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="384" swimtime="00:00:36.93" resultid="3545" heatid="4475" lane="8" entrytime="00:00:36.09" entrycourse="LCM" />
                <RESULT eventid="1366" points="384" swimtime="00:01:18.81" resultid="3546" heatid="4522" lane="4" entrytime="00:01:18.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pamella" lastname="De Machado" birthdate="2002-11-11" gender="F" nation="BRA" license="289846" swrid="5622277" athleteid="3734" externalid="289846">
              <RESULTS>
                <RESULT eventid="1228" points="444" swimtime="00:00:30.93" resultid="3735" heatid="4396" lane="2" />
                <RESULT eventid="1212" points="385" swimtime="00:01:28.09" resultid="3736" heatid="4378" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wilson" lastname="Candido Souza" birthdate="2005-04-06" gender="M" nation="BRA" license="256803" swrid="5600129" athleteid="3616" externalid="256803">
              <RESULTS>
                <RESULT eventid="1088" status="DSQ" swimtime="00:02:54.14" resultid="3617" heatid="4287" lane="8" entrytime="00:02:52.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="516" swimtime="00:00:27.75" resultid="3618" heatid="4303" lane="1" entrytime="00:00:28.09" entrycourse="LCM" />
                <RESULT eventid="1188" points="473" swimtime="00:00:33.30" resultid="3619" heatid="4368" lane="1" entrytime="00:00:33.81" entrycourse="LCM" />
                <RESULT eventid="1220" status="DSQ" swimtime="00:01:16.18" resultid="3620" heatid="4393" lane="2" entrytime="00:01:15.05" entrycourse="LCM" />
                <RESULT eventid="1236" points="477" swimtime="00:00:26.76" resultid="3621" heatid="4418" lane="2" entrytime="00:00:26.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabio" lastname="C Burak" birthdate="2009-08-29" gender="M" nation="BRA" license="343297" swrid="5600126" athleteid="3670" externalid="343297">
              <RESULTS>
                <RESULT eventid="1088" points="459" swimtime="00:02:42.63" resultid="3671" heatid="4287" lane="3" entrytime="00:02:46.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="432" swimtime="00:01:01.95" resultid="3672" heatid="4341" lane="4" entrytime="00:01:03.55" entrycourse="LCM" />
                <RESULT eventid="1188" points="406" swimtime="00:00:35.04" resultid="3673" heatid="4367" lane="3" entrytime="00:00:34.53" entrycourse="LCM" />
                <RESULT eventid="1220" points="417" swimtime="00:01:16.08" resultid="3674" heatid="4392" lane="5" entrytime="00:01:16.01" entrycourse="LCM" />
                <RESULT eventid="1274" points="486" swimtime="00:02:24.96" resultid="3675" heatid="4446" lane="2" entrytime="00:02:33.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Araujo Felix" birthdate="2010-05-27" gender="F" nation="BRA" license="393157" swrid="5622260" athleteid="3716" externalid="393157">
              <RESULTS>
                <RESULT eventid="1064" points="262" swimtime="00:03:12.33" resultid="3717" heatid="4268" lane="1" entrytime="00:03:18.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="328" swimtime="00:01:14.98" resultid="3718" heatid="4323" lane="5" entrytime="00:01:13.62" entrycourse="LCM" />
                <RESULT eventid="1228" points="345" swimtime="00:00:33.64" resultid="3719" heatid="4399" lane="7" entrytime="00:00:34.63" entrycourse="LCM" />
                <RESULT eventid="1282" points="326" swimtime="00:02:43.83" resultid="3720" heatid="4452" lane="6" entrytime="00:02:43.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="265" swimtime="00:01:29.18" resultid="3721" heatid="4519" lane="2" entrytime="00:01:31.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carol" lastname="Nalle Bejes" birthdate="2010-04-20" gender="F" nation="BRA" license="377315" swrid="5588824" athleteid="3652" externalid="377315">
              <RESULTS>
                <RESULT eventid="1080" points="458" swimtime="00:02:58.32" resultid="3653" heatid="4281" lane="5" entrytime="00:02:59.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="412" swimtime="00:01:09.48" resultid="3654" heatid="4325" lane="2" entrytime="00:01:11.16" entrycourse="LCM" />
                <RESULT eventid="1228" points="396" swimtime="00:00:32.14" resultid="3655" heatid="4400" lane="3" entrytime="00:00:32.85" entrycourse="LCM" />
                <RESULT eventid="1212" status="DSQ" swimtime="00:01:24.04" resultid="3656" heatid="4383" lane="8" entrytime="00:01:26.38" entrycourse="LCM" />
                <RESULT eventid="1282" points="379" swimtime="00:02:35.90" resultid="3657" heatid="4455" lane="1" entrytime="00:02:31.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Nogueira Silva" birthdate="2011-08-13" gender="M" nation="BRA" license="367150" swrid="5588832" athleteid="3598" externalid="367150">
              <RESULTS>
                <RESULT eventid="1156" points="362" swimtime="00:01:05.73" resultid="3599" heatid="4337" lane="3" entrytime="00:01:09.44" entrycourse="LCM" />
                <RESULT eventid="1220" points="228" swimtime="00:01:33.03" resultid="3600" heatid="4389" lane="2" entrytime="00:01:31.86" entrycourse="LCM" />
                <RESULT eventid="1236" points="313" swimtime="00:00:30.78" resultid="3601" heatid="4412" lane="1" entrytime="00:00:32.72" entrycourse="LCM" />
                <RESULT eventid="1290" points="340" swimtime="00:02:26.03" resultid="3602" heatid="4462" lane="4" entrytime="00:02:27.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="305" swimtime="00:05:26.69" resultid="3603" heatid="4512" lane="1" entrytime="00:05:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.31" />
                    <SPLIT distance="200" swimtime="00:02:40.72" />
                    <SPLIT distance="300" swimtime="00:04:06.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Guizun Jannuzzi" birthdate="2011-12-27" gender="M" nation="BRA" license="367148" swrid="5588732" athleteid="3588" externalid="367148">
              <RESULTS>
                <RESULT eventid="1156" points="223" swimtime="00:01:17.22" resultid="3589" heatid="4335" lane="7" entrytime="00:01:18.32" entrycourse="LCM" />
                <RESULT eventid="1188" points="163" swimtime="00:00:47.50" resultid="3590" heatid="4363" lane="5" />
                <RESULT eventid="1236" points="208" swimtime="00:00:35.28" resultid="3591" heatid="4407" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Celli Schneider" birthdate="2011-02-21" gender="M" nation="BRA" license="367055" swrid="5588587" athleteid="3576" externalid="367055">
              <RESULTS>
                <RESULT eventid="1072" points="322" swimtime="00:02:43.23" resultid="3577" heatid="4273" lane="4" entrytime="00:02:53.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="225" swimtime="00:03:01.31" resultid="3578" heatid="4351" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="337" swimtime="00:00:30.04" resultid="3579" heatid="4413" lane="2" entrytime="00:00:30.97" entrycourse="LCM" />
                <RESULT eventid="1306" points="340" swimtime="00:00:33.74" resultid="3580" heatid="4479" lane="2" entrytime="00:00:35.28" entrycourse="LCM" />
                <RESULT eventid="1374" points="307" swimtime="00:01:16.45" resultid="3581" heatid="4529" lane="8" entrytime="00:01:14.57" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Fontoura Barros" birthdate="2011-08-04" gender="F" nation="BRA" license="403143" swrid="5676298" athleteid="3688" externalid="403143">
              <RESULTS>
                <RESULT eventid="1080" points="155" swimtime="00:04:15.75" resultid="3689" heatid="4278" lane="6" entrytime="00:04:09.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="168" swimtime="00:01:33.71" resultid="3690" heatid="4320" lane="2" entrytime="00:01:41.04" entrycourse="LCM" />
                <RESULT eventid="1180" points="138" swimtime="00:00:56.30" resultid="3691" heatid="4356" lane="7" entrytime="00:00:59.80" entrycourse="LCM" />
                <RESULT eventid="1228" points="187" swimtime="00:00:41.25" resultid="3692" heatid="4397" lane="5" entrytime="00:00:43.98" entrycourse="LCM" />
                <RESULT eventid="1212" points="149" swimtime="00:02:00.70" resultid="3693" heatid="4379" lane="1" entrytime="00:01:58.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucca" lastname="Maceno Araujo" birthdate="2010-09-29" gender="M" nation="BRA" license="367056" swrid="5588788" athleteid="3582" externalid="367056">
              <RESULTS>
                <RESULT eventid="1104" points="444" swimtime="00:00:29.18" resultid="3583" heatid="4299" lane="4" entrytime="00:00:32.69" entrycourse="LCM" />
                <RESULT eventid="1172" points="274" swimtime="00:02:49.83" resultid="3584" heatid="4351" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="378" swimtime="00:00:28.90" resultid="3585" heatid="4415" lane="8" entrytime="00:00:29.73" entrycourse="LCM" />
                <RESULT eventid="1290" points="375" swimtime="00:02:21.38" resultid="3586" heatid="4464" lane="5" entrytime="00:02:21.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="406" swimtime="00:01:06.73" resultid="3587" heatid="4502" lane="2" entrytime="00:01:09.42" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Ruschel" birthdate="2009-12-28" gender="F" nation="BRA" license="371384" swrid="5600251" athleteid="3634" externalid="371384">
              <RESULTS>
                <RESULT eventid="1096" points="385" swimtime="00:00:33.58" resultid="3635" heatid="4294" lane="1" entrytime="00:00:32.91" entrycourse="LCM" />
                <RESULT eventid="1148" points="542" swimtime="00:01:03.40" resultid="3636" heatid="4329" lane="6" entrytime="00:01:04.30" entrycourse="LCM" />
                <RESULT eventid="1228" points="525" swimtime="00:00:29.25" resultid="3637" heatid="4404" lane="6" entrytime="00:00:29.69" entrycourse="LCM" />
                <RESULT eventid="1282" points="497" swimtime="00:02:22.43" resultid="3638" heatid="4456" lane="2" entrytime="00:02:21.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="407" swimtime="00:00:36.23" resultid="3639" heatid="4474" lane="4" entrytime="00:00:36.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Giuseppe Bulla Lanaro" birthdate="2007-05-22" gender="M" nation="BRA" license="331630" swrid="5600174" athleteid="3493" externalid="331630">
              <RESULTS>
                <RESULT eventid="1124" points="614" swimtime="00:08:51.94" resultid="3494" heatid="4313" lane="5" entrytime="00:09:01.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.53" />
                    <SPLIT distance="200" swimtime="00:02:07.76" />
                    <SPLIT distance="300" swimtime="00:03:14.42" />
                    <SPLIT distance="400" swimtime="00:04:21.61" />
                    <SPLIT distance="500" swimtime="00:05:28.37" />
                    <SPLIT distance="600" swimtime="00:06:36.34" />
                    <SPLIT distance="700" swimtime="00:07:44.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="650" swimtime="00:00:54.09" resultid="3495" heatid="4347" lane="4" entrytime="00:00:54.15" entrycourse="LCM" />
                <RESULT eventid="1236" points="535" swimtime="00:00:25.75" resultid="3496" heatid="4421" lane="8" entrytime="00:00:25.08" entrycourse="LCM" />
                <RESULT eventid="1290" points="640" swimtime="00:01:58.31" resultid="3497" heatid="4469" lane="2" entrytime="00:01:57.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="664" swimtime="00:04:12.14" resultid="3498" heatid="4516" lane="3" entrytime="00:04:14.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.47" />
                    <SPLIT distance="200" swimtime="00:02:02.64" />
                    <SPLIT distance="300" swimtime="00:03:07.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Inoue Kuroda" birthdate="2009-04-18" gender="M" nation="BRA" license="324700" swrid="5600190" athleteid="3523" externalid="324700">
              <RESULTS>
                <RESULT eventid="1156" points="504" swimtime="00:00:58.88" resultid="3524" heatid="4344" lane="7" entrytime="00:00:59.89" entrycourse="LCM" />
                <RESULT eventid="1258" points="547" swimtime="00:17:44.87" resultid="3525" heatid="4432" lane="6" entrytime="00:18:32.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.77" />
                    <SPLIT distance="200" swimtime="00:02:16.54" />
                    <SPLIT distance="300" swimtime="00:03:27.38" />
                    <SPLIT distance="400" swimtime="00:04:38.92" />
                    <SPLIT distance="500" swimtime="00:05:50.62" />
                    <SPLIT distance="600" swimtime="00:07:03.19" />
                    <SPLIT distance="700" swimtime="00:08:15.30" />
                    <SPLIT distance="800" swimtime="00:09:27.52" />
                    <SPLIT distance="900" swimtime="00:10:38.13" />
                    <SPLIT distance="1000" swimtime="00:11:50.14" />
                    <SPLIT distance="1100" swimtime="00:13:01.93" />
                    <SPLIT distance="1200" swimtime="00:14:14.59" />
                    <SPLIT distance="1300" swimtime="00:15:26.93" />
                    <SPLIT distance="1400" swimtime="00:16:38.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="457" swimtime="00:00:27.13" resultid="3526" heatid="4417" lane="3" entrytime="00:00:27.39" entrycourse="LCM" />
                <RESULT eventid="1290" points="502" swimtime="00:02:08.27" resultid="3527" heatid="4466" lane="5" entrytime="00:02:12.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="437" swimtime="00:01:07.95" resultid="3528" heatid="4531" lane="2" entrytime="00:01:08.28" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kethelyn" lastname="Ribeiro Rodrigues" birthdate="2009-04-24" gender="F" nation="BRA" license="367052" swrid="5600244" athleteid="3564" externalid="367052">
              <RESULTS>
                <RESULT eventid="1096" points="258" swimtime="00:00:38.36" resultid="3565" heatid="4291" lane="7" />
                <RESULT eventid="1148" points="447" swimtime="00:01:07.61" resultid="3566" heatid="4326" lane="3" entrytime="00:01:09.30" entrycourse="LCM" />
                <RESULT eventid="1228" points="397" swimtime="00:00:32.10" resultid="3567" heatid="4402" lane="1" entrytime="00:00:31.73" entrycourse="LCM" />
                <RESULT eventid="1282" points="432" swimtime="00:02:29.19" resultid="3568" heatid="4454" lane="6" entrytime="00:02:31.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="310" swimtime="00:01:24.68" resultid="3569" heatid="4520" lane="2" entrytime="00:01:26.29" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Novakoski" birthdate="2009-03-05" gender="F" nation="BRA" license="339136" swrid="5600225" athleteid="3529" externalid="339136">
              <RESULTS>
                <RESULT eventid="1148" points="499" swimtime="00:01:05.19" resultid="3530" heatid="4328" lane="2" entrytime="00:01:06.28" entrycourse="LCM" />
                <RESULT eventid="1180" points="278" swimtime="00:00:44.64" resultid="3531" heatid="4355" lane="4" />
                <RESULT eventid="1228" points="472" swimtime="00:00:30.31" resultid="3532" heatid="4403" lane="2" entrytime="00:00:30.68" entrycourse="LCM" />
                <RESULT eventid="1250" points="321" swimtime="00:11:47.42" resultid="3533" heatid="4426" lane="4" entrytime="00:11:16.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.88" />
                    <SPLIT distance="200" swimtime="00:02:50.22" />
                    <SPLIT distance="300" swimtime="00:04:19.94" />
                    <SPLIT distance="400" swimtime="00:05:50.02" />
                    <SPLIT distance="500" swimtime="00:07:20.19" />
                    <SPLIT distance="600" swimtime="00:08:52.06" />
                    <SPLIT distance="700" swimtime="00:10:23.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="419" swimtime="00:02:30.74" resultid="3534" heatid="4455" lane="8" entrytime="00:02:31.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cardim Martins" birthdate="2010-09-01" gender="F" nation="BRA" license="390920" swrid="5600130" athleteid="3722" externalid="390920">
              <RESULTS>
                <RESULT eventid="1064" points="289" swimtime="00:03:06.22" resultid="3723" heatid="4268" lane="7" entrytime="00:03:10.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="294" swimtime="00:01:17.71" resultid="3724" heatid="4321" lane="4" entrytime="00:01:22.86" entrycourse="LCM" />
                <RESULT eventid="1282" points="290" swimtime="00:02:50.44" resultid="3725" heatid="4451" lane="5" entrytime="00:02:52.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="284" swimtime="00:00:40.84" resultid="3726" heatid="4472" lane="6" entrytime="00:00:42.89" entrycourse="LCM" />
                <RESULT eventid="1366" points="277" swimtime="00:01:27.89" resultid="3727" heatid="4519" lane="4" entrytime="00:01:28.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Lopes Rempel" birthdate="2010-09-25" gender="M" nation="BRA" license="399739" swrid="5653294" athleteid="3676" externalid="399739">
              <RESULTS>
                <RESULT eventid="1072" points="248" swimtime="00:02:57.91" resultid="3677" heatid="4273" lane="5" entrytime="00:02:57.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="289" swimtime="00:01:10.80" resultid="3678" heatid="4334" lane="5" entrytime="00:01:21.79" entrycourse="LCM" />
                <RESULT eventid="1236" points="302" swimtime="00:00:31.14" resultid="3679" heatid="4411" lane="6" entrytime="00:00:34.69" entrycourse="LCM" />
                <RESULT eventid="1290" points="266" swimtime="00:02:38.46" resultid="3680" heatid="4461" lane="8" entrytime="00:02:41.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="235" swimtime="00:01:23.52" resultid="3681" heatid="4527" lane="7" entrytime="00:01:25.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Gelenski Pelaio" birthdate="2005-10-10" gender="M" nation="BRA" license="281473" swrid="5600173" athleteid="3622" externalid="281473">
              <RESULTS>
                <RESULT eventid="1104" points="573" swimtime="00:00:26.80" resultid="3623" heatid="4304" lane="2" entrytime="00:00:26.69" entrycourse="LCM" />
                <RESULT eventid="1188" points="461" swimtime="00:00:33.59" resultid="3624" heatid="4362" lane="2" />
                <RESULT eventid="1236" points="590" swimtime="00:00:24.92" resultid="3625" heatid="4421" lane="7" entrytime="00:00:25.01" entrycourse="LCM" />
                <RESULT eventid="1290" points="546" swimtime="00:02:04.76" resultid="3626" heatid="4467" lane="5" entrytime="00:02:07.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="555" swimtime="00:01:00.14" resultid="3627" heatid="4505" lane="1" entrytime="00:01:00.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Nalle Bejes" birthdate="2010-04-20" gender="F" nation="BRA" license="377323" swrid="5588826" athleteid="3658" externalid="377323">
              <RESULTS>
                <RESULT eventid="1080" points="364" swimtime="00:03:12.56" resultid="3659" heatid="4280" lane="3" entrytime="00:03:09.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="389" swimtime="00:01:10.83" resultid="3660" heatid="4322" lane="5" entrytime="00:01:15.58" entrycourse="LCM" />
                <RESULT eventid="1212" points="371" swimtime="00:01:29.24" resultid="3661" heatid="4382" lane="7" entrytime="00:01:29.05" entrycourse="LCM" />
                <RESULT eventid="1282" points="392" swimtime="00:02:34.09" resultid="3662" heatid="4451" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="264" swimtime="00:01:29.27" resultid="3663" heatid="4519" lane="7" entrytime="00:01:31.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Bello Costa Lange" birthdate="2010-09-13" gender="M" nation="BRA" license="367152" swrid="5588547" athleteid="3604" externalid="367152">
              <RESULTS>
                <RESULT eventid="1104" points="338" swimtime="00:00:31.96" resultid="3605" heatid="4300" lane="8" entrytime="00:00:32.42" entrycourse="LCM" />
                <RESULT eventid="1140" status="DSQ" swimtime="00:05:47.51" resultid="3606" heatid="4317" lane="8" entrytime="00:06:03.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.33" />
                    <SPLIT distance="200" swimtime="00:02:49.30" />
                    <SPLIT distance="300" swimtime="00:04:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="392" swimtime="00:19:49.88" resultid="3607" heatid="4431" lane="5" entrytime="00:20:08.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.44" />
                    <SPLIT distance="200" swimtime="00:02:30.66" />
                    <SPLIT distance="300" swimtime="00:03:49.87" />
                    <SPLIT distance="400" swimtime="00:05:10.77" />
                    <SPLIT distance="500" swimtime="00:06:32.22" />
                    <SPLIT distance="600" swimtime="00:07:52.48" />
                    <SPLIT distance="700" swimtime="00:09:13.77" />
                    <SPLIT distance="800" swimtime="00:10:34.44" />
                    <SPLIT distance="900" swimtime="00:11:54.20" />
                    <SPLIT distance="1000" swimtime="00:13:14.07" />
                    <SPLIT distance="1100" swimtime="00:14:33.67" />
                    <SPLIT distance="1200" swimtime="00:15:53.62" />
                    <SPLIT distance="1300" swimtime="00:17:14.17" />
                    <SPLIT distance="1400" swimtime="00:18:33.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="351" swimtime="00:02:24.48" resultid="3608" heatid="4464" lane="8" entrytime="00:02:24.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="300" swimtime="00:01:13.79" resultid="3609" heatid="4501" lane="6" entrytime="00:01:14.27" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wagner" lastname="Junior Cabral Gama" birthdate="2007-07-22" gender="M" nation="BRA" license="345334" swrid="5723027" athleteid="3737" externalid="345334">
              <RESULTS>
                <RESULT eventid="1104" points="405" swimtime="00:00:30.09" resultid="3738" heatid="4296" lane="6" />
                <RESULT eventid="1156" points="466" swimtime="00:01:00.43" resultid="3739" heatid="4343" lane="8" entrytime="00:01:01.90" entrycourse="LCM" />
                <RESULT eventid="1236" points="452" swimtime="00:00:27.23" resultid="3740" heatid="4406" lane="4" />
                <RESULT eventid="1290" points="406" swimtime="00:02:17.72" resultid="3741" heatid="4458" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="380" swimtime="00:01:11.19" resultid="3742" heatid="4530" lane="2" entrytime="00:01:10.44" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Murara" birthdate="1991-04-12" gender="M" nation="BRA" license="386866" swrid="5622296" athleteid="3743" externalid="386866">
              <RESULTS>
                <RESULT eventid="1104" points="612" swimtime="00:00:26.22" resultid="3744" heatid="4304" lane="6" entrytime="00:00:26.41" entrycourse="LCM" />
                <RESULT eventid="1236" points="576" swimtime="00:00:25.12" resultid="3745" heatid="4421" lane="4" entrytime="00:00:24.63" entrycourse="LCM" />
                <RESULT eventid="1306" points="559" swimtime="00:00:28.58" resultid="3746" heatid="4482" lane="5" entrytime="00:00:28.42" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Leticia Durat" birthdate="2008-02-09" gender="F" nation="BRA" license="331636" swrid="5600200" athleteid="3511" externalid="331636">
              <RESULTS>
                <RESULT eventid="1080" points="310" swimtime="00:03:23.23" resultid="3512" heatid="4280" lane="6" entrytime="00:03:10.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="428" swimtime="00:01:08.60" resultid="3513" heatid="4327" lane="8" entrytime="00:01:08.25" entrycourse="LCM" />
                <RESULT eventid="1180" points="371" swimtime="00:00:40.57" resultid="3514" heatid="4359" lane="8" entrytime="00:00:38.23" entrycourse="LCM" />
                <RESULT eventid="1228" points="457" swimtime="00:00:30.64" resultid="3515" heatid="4403" lane="3" entrytime="00:00:30.43" entrycourse="LCM" />
                <RESULT eventid="1212" points="338" swimtime="00:01:32.00" resultid="3516" heatid="4382" lane="5" entrytime="00:01:27.33" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabrizio" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="M" nation="BRA" license="344303" swrid="5559846" athleteid="3517" externalid="344303">
              <RESULTS>
                <RESULT eventid="1104" points="525" swimtime="00:00:27.60" resultid="3518" heatid="4302" lane="4" entrytime="00:00:28.22" entrycourse="LCM" />
                <RESULT eventid="1156" points="471" swimtime="00:01:00.19" resultid="3519" heatid="4344" lane="5" entrytime="00:00:59.78" entrycourse="LCM" />
                <RESULT eventid="1236" points="450" swimtime="00:00:27.28" resultid="3520" heatid="4419" lane="6" entrytime="00:00:26.44" entrycourse="LCM" />
                <RESULT eventid="1306" points="431" swimtime="00:00:31.16" resultid="3521" heatid="4481" lane="2" entrytime="00:00:31.45" entrycourse="LCM" />
                <RESULT eventid="1342" points="490" swimtime="00:01:02.69" resultid="3522" heatid="4503" lane="7" entrytime="00:01:04.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Ieger" birthdate="2009-02-20" gender="M" nation="BRA" license="356888" swrid="5600180" athleteid="3547" externalid="356888">
              <RESULTS>
                <RESULT eventid="1156" points="465" swimtime="00:01:00.45" resultid="3548" heatid="4344" lane="8" entrytime="00:01:00.53" entrycourse="LCM" />
                <RESULT eventid="1188" points="418" swimtime="00:00:34.68" resultid="3549" heatid="4367" lane="6" entrytime="00:00:34.80" entrycourse="LCM" />
                <RESULT eventid="1220" points="364" swimtime="00:01:19.62" resultid="3550" heatid="4391" lane="4" entrytime="00:01:20.41" entrycourse="LCM" />
                <RESULT eventid="1236" points="431" swimtime="00:00:27.67" resultid="3551" heatid="4417" lane="5" entrytime="00:00:27.39" entrycourse="LCM" />
                <RESULT eventid="1290" points="408" swimtime="00:02:17.42" resultid="3552" heatid="4465" lane="2" entrytime="00:02:18.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Zanatta Flizikowski" birthdate="2010-01-08" gender="F" nation="BRA" license="367051" swrid="5588969" athleteid="3704" externalid="367051">
              <RESULTS>
                <RESULT eventid="1096" points="362" swimtime="00:00:34.27" resultid="3705" heatid="4291" lane="1" />
                <RESULT eventid="1148" points="462" swimtime="00:01:06.87" resultid="3706" heatid="4328" lane="6" entrytime="00:01:06.16" entrycourse="LCM" />
                <RESULT eventid="1228" points="423" swimtime="00:00:31.43" resultid="3707" heatid="4402" lane="6" entrytime="00:00:31.16" entrycourse="LCM" />
                <RESULT eventid="1282" points="408" swimtime="00:02:32.14" resultid="3708" heatid="4456" lane="1" entrytime="00:02:24.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="290" swimtime="00:01:23.79" resultid="3709" heatid="4496" lane="7" entrytime="00:01:18.96" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Schlickmann Assis" birthdate="2003-07-24" gender="F" nation="BRA" license="303874" swrid="5600257" athleteid="3553" externalid="303874">
              <RESULTS>
                <RESULT eventid="1148" points="494" swimtime="00:01:05.40" resultid="3554" heatid="4320" lane="1" />
                <RESULT eventid="1180" points="488" swimtime="00:00:37.02" resultid="3555" heatid="4359" lane="5" entrytime="00:00:35.38" entrycourse="LCM" />
                <RESULT eventid="1228" points="456" swimtime="00:00:30.67" resultid="3556" heatid="4405" lane="1" entrytime="00:00:29.24" entrycourse="LCM" />
                <RESULT eventid="1212" points="492" swimtime="00:01:21.19" resultid="3557" heatid="4384" lane="6" entrytime="00:01:17.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Helena Vieira Jussen" birthdate="2011-12-29" gender="F" nation="BRA" license="372282" swrid="5588740" athleteid="3640" externalid="372282">
              <RESULTS>
                <RESULT eventid="1080" points="326" swimtime="00:03:19.81" resultid="3641" heatid="4279" lane="7" entrytime="00:03:26.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="155" swimtime="00:00:45.47" resultid="3642" heatid="4291" lane="5" entrytime="00:00:53.05" entrycourse="LCM" />
                <RESULT eventid="1212" points="294" swimtime="00:01:36.40" resultid="3643" heatid="4381" lane="1" entrytime="00:01:33.96" entrycourse="LCM" />
                <RESULT eventid="1282" points="288" swimtime="00:02:50.88" resultid="3644" heatid="4451" lane="3" entrytime="00:02:53.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="227" swimtime="00:00:44.03" resultid="3645" heatid="4471" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Blansky Hagebock" birthdate="2008-08-15" gender="M" nation="BRA" license="339123" swrid="5455418" athleteid="3535" externalid="339123">
              <RESULTS>
                <RESULT eventid="1104" points="462" swimtime="00:00:28.79" resultid="3536" heatid="4301" lane="4" entrytime="00:00:29.45" entrycourse="LCM" />
                <RESULT eventid="1156" points="549" swimtime="00:00:57.22" resultid="3537" heatid="4346" lane="3" entrytime="00:00:57.25" entrycourse="LCM" />
                <RESULT eventid="1236" points="511" swimtime="00:00:26.15" resultid="3538" heatid="4420" lane="7" entrytime="00:00:25.64" entrycourse="LCM" />
                <RESULT eventid="1290" points="490" swimtime="00:02:09.30" resultid="3539" heatid="4467" lane="7" entrytime="00:02:10.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="470" swimtime="00:04:42.98" resultid="3540" heatid="4511" lane="3" entrytime="00:05:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.56" />
                    <SPLIT distance="200" swimtime="00:02:18.43" />
                    <SPLIT distance="300" swimtime="00:03:32.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Breno" lastname="Borges Piekarzievicz" birthdate="2011-11-11" gender="M" nation="BRA" license="403144" swrid="5676295" athleteid="3694" externalid="403144">
              <RESULTS>
                <RESULT eventid="1156" points="138" swimtime="00:01:30.66" resultid="3695" heatid="4334" lane="8" entrytime="00:01:45.09" entrycourse="LCM" />
                <RESULT eventid="1188" points="125" swimtime="00:00:51.77" resultid="3696" heatid="4363" lane="4" entrytime="00:00:58.95" entrycourse="LCM" />
                <RESULT eventid="1220" points="124" swimtime="00:01:53.99" resultid="3697" heatid="4387" lane="7" entrytime="00:01:55.85" entrycourse="LCM" />
                <RESULT eventid="1236" points="125" swimtime="00:00:41.79" resultid="3698" heatid="4410" lane="3" entrytime="00:00:47.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Garcia Reschetti Rubbo" birthdate="2011-08-06" gender="F" nation="BRA" license="367053" swrid="5588720" athleteid="3570" externalid="367053">
              <RESULTS>
                <RESULT eventid="1080" points="318" swimtime="00:03:21.40" resultid="3571" heatid="4279" lane="1" entrytime="00:03:31.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="203" swimtime="00:00:41.52" resultid="3572" heatid="4290" lane="3" />
                <RESULT eventid="1180" points="274" swimtime="00:00:44.88" resultid="3573" heatid="4357" lane="1" entrytime="00:00:45.84" entrycourse="LCM" />
                <RESULT eventid="1228" points="345" swimtime="00:00:33.65" resultid="3574" heatid="4398" lane="4" entrytime="00:00:36.05" entrycourse="LCM" />
                <RESULT eventid="1212" points="291" swimtime="00:01:36.67" resultid="3575" heatid="4380" lane="3" entrytime="00:01:38.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Marques" birthdate="2007-06-29" gender="M" nation="BRA" license="367257" swrid="5600213" athleteid="3728" externalid="367257">
              <RESULTS>
                <RESULT eventid="1124" points="339" swimtime="00:10:48.22" resultid="3729" heatid="4310" lane="7" entrytime="00:11:24.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.52" />
                    <SPLIT distance="200" swimtime="00:02:30.35" />
                    <SPLIT distance="300" swimtime="00:03:51.44" />
                    <SPLIT distance="400" swimtime="00:05:14.46" />
                    <SPLIT distance="500" swimtime="00:06:38.43" />
                    <SPLIT distance="600" swimtime="00:08:02.99" />
                    <SPLIT distance="700" swimtime="00:09:27.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="398" swimtime="00:01:03.70" resultid="3730" heatid="4343" lane="1" entrytime="00:01:01.85" entrycourse="LCM" />
                <RESULT eventid="1258" points="363" swimtime="00:20:20.89" resultid="3731" heatid="4430" lane="8" entrytime="00:21:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.63" />
                    <SPLIT distance="200" swimtime="00:02:34.80" />
                    <SPLIT distance="300" swimtime="00:03:57.38" />
                    <SPLIT distance="400" swimtime="00:05:19.85" />
                    <SPLIT distance="500" swimtime="00:06:43.52" />
                    <SPLIT distance="600" swimtime="00:08:06.20" />
                    <SPLIT distance="700" swimtime="00:09:30.01" />
                    <SPLIT distance="800" swimtime="00:10:52.04" />
                    <SPLIT distance="900" swimtime="00:12:14.50" />
                    <SPLIT distance="1000" swimtime="00:13:37.66" />
                    <SPLIT distance="1100" swimtime="00:15:00.32" />
                    <SPLIT distance="1200" swimtime="00:16:22.91" />
                    <SPLIT distance="1300" swimtime="00:17:44.87" />
                    <SPLIT distance="1400" swimtime="00:19:05.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="375" swimtime="00:02:21.39" resultid="3732" heatid="4465" lane="7" entrytime="00:02:19.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="370" swimtime="00:05:06.30" resultid="3733" heatid="4514" lane="3" entrytime="00:04:57.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.87" />
                    <SPLIT distance="200" swimtime="00:02:27.16" />
                    <SPLIT distance="300" swimtime="00:03:46.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="F" nation="BRA" license="344301" swrid="5569976" athleteid="3481" externalid="344301">
              <RESULTS>
                <RESULT eventid="1096" points="551" swimtime="00:00:29.79" resultid="3482" heatid="4294" lane="5" entrytime="00:00:30.16" entrycourse="LCM" />
                <RESULT eventid="1164" points="564" swimtime="00:02:27.40" resultid="3483" heatid="4350" lane="5" entrytime="00:02:30.90" entrycourse="LCM" />
                <RESULT eventid="1228" points="569" swimtime="00:00:28.49" resultid="3484" heatid="4405" lane="2" entrytime="00:00:28.43" entrycourse="LCM" />
                <RESULT eventid="1282" points="639" swimtime="00:02:10.99" resultid="3485" heatid="4457" lane="8" entrytime="00:02:17.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="598" swimtime="00:01:05.83" resultid="3486" heatid="4497" lane="5" entrytime="00:01:04.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Vianna" birthdate="2011-01-31" gender="M" nation="BRA" license="371380" swrid="5588947" athleteid="3628" externalid="371380">
              <RESULTS>
                <RESULT eventid="1104" points="332" swimtime="00:00:32.14" resultid="3629" heatid="4299" lane="2" entrytime="00:00:34.31" entrycourse="LCM" />
                <RESULT eventid="1156" points="368" swimtime="00:01:05.38" resultid="3630" heatid="4340" lane="1" entrytime="00:01:06.52" entrycourse="LCM" />
                <RESULT eventid="1236" points="345" swimtime="00:00:29.80" resultid="3631" heatid="4413" lane="4" entrytime="00:00:30.48" entrycourse="LCM" />
                <RESULT eventid="1290" points="354" swimtime="00:02:24.10" resultid="3632" heatid="4462" lane="5" entrytime="00:02:30.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="309" swimtime="00:01:13.11" resultid="3633" heatid="4501" lane="1" entrytime="00:01:15.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Marques Machado" birthdate="2010-02-17" gender="M" nation="BRA" license="390918" swrid="5600212" athleteid="3664" externalid="390918">
              <RESULTS>
                <RESULT eventid="1124" points="339" swimtime="00:10:48.17" resultid="3665" heatid="4311" lane="1" entrytime="00:10:54.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.52" />
                    <SPLIT distance="200" swimtime="00:02:34.99" />
                    <SPLIT distance="300" swimtime="00:03:56.39" />
                    <SPLIT distance="400" swimtime="00:05:19.96" />
                    <SPLIT distance="500" swimtime="00:06:44.02" />
                    <SPLIT distance="600" swimtime="00:08:07.56" />
                    <SPLIT distance="700" swimtime="00:09:29.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="311" swimtime="00:00:32.85" resultid="3666" heatid="4298" lane="6" entrytime="00:00:38.21" entrycourse="LCM" />
                <RESULT eventid="1258" points="342" swimtime="00:20:44.62" resultid="3667" heatid="4431" lane="6" entrytime="00:20:49.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.32" />
                    <SPLIT distance="200" swimtime="00:02:31.23" />
                    <SPLIT distance="300" swimtime="00:03:55.35" />
                    <SPLIT distance="400" swimtime="00:05:24.01" />
                    <SPLIT distance="500" swimtime="00:06:47.82" />
                    <SPLIT distance="600" swimtime="00:08:12.26" />
                    <SPLIT distance="700" swimtime="00:09:35.21" />
                    <SPLIT distance="800" swimtime="00:10:57.57" />
                    <SPLIT distance="900" swimtime="00:12:20.54" />
                    <SPLIT distance="1000" swimtime="00:13:45.19" />
                    <SPLIT distance="1100" swimtime="00:15:09.03" />
                    <SPLIT distance="1200" swimtime="00:16:33.47" />
                    <SPLIT distance="1300" swimtime="00:18:00.25" />
                    <SPLIT distance="1400" swimtime="00:19:24.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="360" swimtime="00:02:23.31" resultid="3668" heatid="4464" lane="2" entrytime="00:02:22.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="256" swimtime="00:01:17.83" resultid="3669" heatid="4500" lane="3" entrytime="00:01:17.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Pinterich Almeida" birthdate="2005-03-13" gender="M" nation="BRA" license="330749" swrid="5600235" athleteid="3558" externalid="330749">
              <RESULTS>
                <RESULT eventid="1072" points="487" swimtime="00:02:22.24" resultid="3559" heatid="4276" lane="4" entrytime="00:02:20.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="654" swimtime="00:00:53.98" resultid="3560" heatid="4348" lane="1" entrytime="00:00:53.65" entrycourse="LCM" />
                <RESULT eventid="1290" points="663" swimtime="00:01:56.94" resultid="3561" heatid="4469" lane="6" entrytime="00:01:56.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1306" points="520" swimtime="00:00:29.27" resultid="3562" heatid="4482" lane="7" entrytime="00:00:28.82" entrycourse="LCM" />
                <RESULT eventid="1374" points="552" swimtime="00:01:02.87" resultid="3563" heatid="4533" lane="1" entrytime="00:01:01.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emily" lastname="Sayuri Tangueria De Lima" birthdate="2010-06-11" gender="F" nation="BRA" license="367215" swrid="5588901" athleteid="3610" externalid="367215">
              <RESULTS>
                <RESULT eventid="1096" points="406" swimtime="00:00:32.97" resultid="3611" heatid="4293" lane="6" entrytime="00:00:36.02" entrycourse="LCM" />
                <RESULT eventid="1164" points="318" swimtime="00:02:58.39" resultid="3612" heatid="4350" lane="1" entrytime="00:02:58.43" entrycourse="LCM" />
                <RESULT eventid="1250" points="390" swimtime="00:11:03.13" resultid="3613" heatid="4427" lane="7" entrytime="00:10:54.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.37" />
                    <SPLIT distance="200" swimtime="00:02:39.42" />
                    <SPLIT distance="300" swimtime="00:04:03.29" />
                    <SPLIT distance="400" swimtime="00:05:28.45" />
                    <SPLIT distance="500" swimtime="00:06:53.26" />
                    <SPLIT distance="600" swimtime="00:08:18.23" />
                    <SPLIT distance="700" swimtime="00:09:41.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="460" swimtime="00:02:26.14" resultid="3614" heatid="4449" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="374" swimtime="00:01:16.94" resultid="3615" heatid="4496" lane="5" entrytime="00:01:16.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="19" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1208" points="598" swimtime="00:08:16.53" resultid="3752" heatid="4375" lane="5" entrytime="00:08:17.90">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.43" />
                    <SPLIT distance="200" swimtime="00:02:09.60" />
                    <SPLIT distance="300" swimtime="00:03:07.57" />
                    <SPLIT distance="400" swimtime="00:04:09.86" />
                    <SPLIT distance="500" swimtime="00:05:09.84" />
                    <SPLIT distance="600" swimtime="00:06:16.76" />
                    <SPLIT distance="700" swimtime="00:07:14.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3616" number="1" />
                    <RELAYPOSITION athleteid="3558" number="2" />
                    <RELAYPOSITION athleteid="3622" number="3" />
                    <RELAYPOSITION athleteid="3493" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1206" points="503" swimtime="00:08:46.17" resultid="3753" heatid="4374" lane="8" entrytime="00:08:17.83">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.51" />
                    <SPLIT distance="200" swimtime="00:02:07.17" />
                    <SPLIT distance="300" swimtime="00:03:10.94" />
                    <SPLIT distance="400" swimtime="00:04:20.70" />
                    <SPLIT distance="500" swimtime="00:05:25.53" />
                    <SPLIT distance="600" swimtime="00:06:36.12" />
                    <SPLIT distance="700" swimtime="00:07:38.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3523" number="1" />
                    <RELAYPOSITION athleteid="3517" number="2" />
                    <RELAYPOSITION athleteid="3670" number="3" />
                    <RELAYPOSITION athleteid="3535" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1328" points="470" swimtime="00:04:25.95" resultid="3754" heatid="4490" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.14" />
                    <SPLIT distance="200" swimtime="00:02:22.68" />
                    <SPLIT distance="300" swimtime="00:03:25.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3523" number="1" />
                    <RELAYPOSITION athleteid="3670" number="2" />
                    <RELAYPOSITION athleteid="3517" number="3" />
                    <RELAYPOSITION athleteid="3547" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1396" points="483" swimtime="00:03:59.86" resultid="3757" heatid="4541" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.06" />
                    <SPLIT distance="200" swimtime="00:02:00.70" />
                    <SPLIT distance="300" swimtime="00:03:01.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3517" number="1" />
                    <RELAYPOSITION athleteid="3547" number="2" />
                    <RELAYPOSITION athleteid="3670" number="3" />
                    <RELAYPOSITION athleteid="3523" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1332" points="533" swimtime="00:04:14.96" resultid="3755" heatid="4492" lane="3" entrytime="00:04:15.67">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.73" />
                    <SPLIT distance="200" swimtime="00:02:18.49" />
                    <SPLIT distance="300" swimtime="00:03:20.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3558" number="1" />
                    <RELAYPOSITION athleteid="3616" number="2" />
                    <RELAYPOSITION athleteid="3622" number="3" />
                    <RELAYPOSITION athleteid="3493" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1400" points="610" swimtime="00:03:41.95" resultid="3756" heatid="4543" lane="5" entrytime="00:03:42.13">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.29" />
                    <SPLIT distance="200" swimtime="00:01:53.98" />
                    <SPLIT distance="300" swimtime="00:02:47.61" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3622" number="1" />
                    <RELAYPOSITION athleteid="3616" number="2" />
                    <RELAYPOSITION athleteid="3558" number="3" />
                    <RELAYPOSITION athleteid="3493" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1204" points="380" swimtime="00:09:37.85" resultid="3771" heatid="4373" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.25" />
                    <SPLIT distance="200" swimtime="00:02:19.05" />
                    <SPLIT distance="300" swimtime="00:03:30.45" />
                    <SPLIT distance="500" swimtime="00:05:53.07" />
                    <SPLIT distance="600" swimtime="00:07:06.60" />
                    <SPLIT distance="700" swimtime="00:08:18.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3582" number="1" />
                    <RELAYPOSITION athleteid="3664" number="2" />
                    <RELAYPOSITION athleteid="3604" number="3" />
                    <RELAYPOSITION athleteid="3598" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1324" points="322" swimtime="00:05:01.68" resultid="3772" heatid="4488" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.60" />
                    <SPLIT distance="200" swimtime="00:02:43.15" />
                    <SPLIT distance="300" swimtime="00:03:55.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3576" number="1" />
                    <RELAYPOSITION athleteid="3592" number="2" />
                    <RELAYPOSITION athleteid="3628" number="3" />
                    <RELAYPOSITION athleteid="3598" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1392" points="330" swimtime="00:04:32.37" resultid="3774" heatid="4539" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.74" />
                    <SPLIT distance="200" swimtime="00:02:13.32" />
                    <SPLIT distance="300" swimtime="00:03:20.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3628" number="1" />
                    <RELAYPOSITION athleteid="3598" number="2" />
                    <RELAYPOSITION athleteid="3576" number="3" />
                    <RELAYPOSITION athleteid="3592" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1326" points="298" swimtime="00:05:09.31" resultid="3773" heatid="4489" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.92" />
                    <SPLIT distance="200" swimtime="00:02:53.50" />
                    <SPLIT distance="300" swimtime="00:04:02.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3676" number="1" />
                    <RELAYPOSITION athleteid="3604" number="2" />
                    <RELAYPOSITION athleteid="3582" number="3" />
                    <RELAYPOSITION athleteid="3664" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1394" points="361" swimtime="00:04:24.27" resultid="3775" heatid="4540" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.76" />
                    <SPLIT distance="200" swimtime="00:02:08.28" />
                    <SPLIT distance="300" swimtime="00:03:14.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3582" number="1" />
                    <RELAYPOSITION athleteid="3664" number="2" />
                    <RELAYPOSITION athleteid="3604" number="3" />
                    <RELAYPOSITION athleteid="3676" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1324" points="177" swimtime="00:06:08.05" resultid="3761" heatid="4488" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3646" number="1" />
                    <RELAYPOSITION athleteid="3588" number="2" />
                    <RELAYPOSITION athleteid="3682" number="3" />
                    <RELAYPOSITION athleteid="3694" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1392" points="218" swimtime="00:05:12.38" resultid="3762" heatid="4539" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.28" />
                    <SPLIT distance="200" swimtime="00:02:23.41" />
                    <SPLIT distance="300" swimtime="00:03:43.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3682" number="1" />
                    <RELAYPOSITION athleteid="3646" number="2" />
                    <RELAYPOSITION athleteid="3588" number="3" />
                    <RELAYPOSITION athleteid="3694" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1198" points="496" swimtime="00:09:37.59" resultid="3747" heatid="4371" lane="7" entrytime="00:09:15.23">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.18" />
                    <SPLIT distance="200" swimtime="00:02:20.98" />
                    <SPLIT distance="300" swimtime="00:03:31.94" />
                    <SPLIT distance="400" swimtime="00:04:49.37" />
                    <SPLIT distance="500" swimtime="00:06:01.83" />
                    <SPLIT distance="700" swimtime="00:08:25.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3634" number="1" />
                    <RELAYPOSITION athleteid="3529" number="2" />
                    <RELAYPOSITION athleteid="3541" number="3" />
                    <RELAYPOSITION athleteid="3481" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1318" points="409" swimtime="00:05:10.14" resultid="3748" heatid="4485" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.46" />
                    <SPLIT distance="200" swimtime="00:02:58.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3541" number="1" />
                    <RELAYPOSITION athleteid="3529" number="2" />
                    <RELAYPOSITION athleteid="3481" number="3" />
                    <RELAYPOSITION athleteid="3634" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1386" points="534" swimtime="00:04:16.25" resultid="3751" heatid="4536" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.38" />
                    <SPLIT distance="200" swimtime="00:02:04.09" />
                    <SPLIT distance="300" swimtime="00:03:10.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3481" number="1" />
                    <RELAYPOSITION athleteid="3634" number="2" />
                    <RELAYPOSITION athleteid="3541" number="3" />
                    <RELAYPOSITION athleteid="3529" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1322" status="WDR" swimtime="00:00:00.00" resultid="3749" heatid="4487" lane="6" entrytime="00:04:44.99" />
                <RESULT eventid="1390" points="459" swimtime="00:04:29.51" resultid="3750" heatid="4538" lane="7" entrytime="00:04:07.12">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.15" />
                    <SPLIT distance="200" swimtime="00:02:08.68" />
                    <SPLIT distance="300" swimtime="00:03:20.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3553" number="1" />
                    <RELAYPOSITION athleteid="3499" number="2" />
                    <RELAYPOSITION athleteid="3734" number="3" />
                    <RELAYPOSITION athleteid="3487" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1196" points="441" swimtime="00:10:00.63" resultid="3766" heatid="4370" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.35" />
                    <SPLIT distance="200" swimtime="00:02:29.29" />
                    <SPLIT distance="300" swimtime="00:03:39.80" />
                    <SPLIT distance="400" swimtime="00:04:57.04" />
                    <SPLIT distance="500" swimtime="00:06:09.78" />
                    <SPLIT distance="600" swimtime="00:07:26.90" />
                    <SPLIT distance="700" swimtime="00:08:41.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3610" number="1" />
                    <RELAYPOSITION athleteid="3704" number="2" />
                    <RELAYPOSITION athleteid="3652" number="3" />
                    <RELAYPOSITION athleteid="3658" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1314" status="DSQ" swimtime="00:06:59.02" resultid="3767" heatid="4483" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.49" />
                    <SPLIT distance="200" swimtime="00:03:28.51" />
                    <SPLIT distance="300" swimtime="00:05:25.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3699" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="3570" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="3640" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="3688" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1382" points="248" swimtime="00:05:30.94" resultid="3770" heatid="4534" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.17" />
                    <SPLIT distance="200" swimtime="00:02:37.34" />
                    <SPLIT distance="300" swimtime="00:03:59.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3570" number="1" />
                    <RELAYPOSITION athleteid="3640" number="2" />
                    <RELAYPOSITION athleteid="3699" number="3" />
                    <RELAYPOSITION athleteid="3688" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1316" points="344" swimtime="00:05:28.57" resultid="3768" heatid="4484" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.74" />
                    <SPLIT distance="200" swimtime="00:02:56.98" />
                    <SPLIT distance="300" swimtime="00:04:17.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3658" number="1" />
                    <RELAYPOSITION athleteid="3652" number="2" />
                    <RELAYPOSITION athleteid="3610" number="3" />
                    <RELAYPOSITION athleteid="3704" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1384" points="435" swimtime="00:04:34.44" resultid="3769" heatid="4535" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.53" />
                    <SPLIT distance="200" swimtime="00:02:15.76" />
                    <SPLIT distance="300" swimtime="00:03:24.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3704" number="1" />
                    <RELAYPOSITION athleteid="3610" number="2" />
                    <RELAYPOSITION athleteid="3652" number="3" />
                    <RELAYPOSITION athleteid="3658" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1248" points="505" swimtime="00:04:33.16" resultid="3758" heatid="4425" lane="5" entrytime="00:04:25.46">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.79" />
                    <SPLIT distance="200" swimtime="00:02:29.19" />
                    <SPLIT distance="300" swimtime="00:03:30.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3487" number="1" />
                    <RELAYPOSITION athleteid="3616" number="2" />
                    <RELAYPOSITION athleteid="3622" number="3" />
                    <RELAYPOSITION athleteid="3499" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1246" points="366" swimtime="00:05:03.92" resultid="3759" heatid="4424" lane="5" entrytime="00:04:28.71">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3564" number="1" />
                    <RELAYPOSITION athleteid="3511" number="2" />
                    <RELAYPOSITION athleteid="3505" number="3" />
                    <RELAYPOSITION athleteid="3535" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1244" points="365" swimtime="00:05:04.38" resultid="3760" heatid="4423" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.37" />
                    <SPLIT distance="200" swimtime="00:02:53.40" />
                    <SPLIT distance="300" swimtime="00:03:55.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3670" number="1" />
                    <RELAYPOSITION athleteid="3529" number="2" />
                    <RELAYPOSITION athleteid="3517" number="3" />
                    <RELAYPOSITION athleteid="3541" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1112" points="329" swimtime="00:05:15.04" resultid="3776" heatid="4305" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.81" />
                    <SPLIT distance="200" swimtime="00:02:48.87" />
                    <SPLIT distance="300" swimtime="00:04:00.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3576" number="1" />
                    <RELAYPOSITION athleteid="3640" number="2" />
                    <RELAYPOSITION athleteid="3628" number="3" />
                    <RELAYPOSITION athleteid="3570" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1114" status="DSQ" swimtime="00:04:56.32" resultid="3777" heatid="4307" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.19" />
                    <SPLIT distance="200" swimtime="00:02:41.05" />
                    <SPLIT distance="300" swimtime="00:03:49.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3604" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="3652" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="3582" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="3704" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1112" status="DSQ" swimtime="00:06:27.99" resultid="3763" heatid="4306" lane="2" entrytime="00:05:50.63">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:03:55.30" />
                    <SPLIT distance="300" swimtime="00:05:21.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3699" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="3688" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="3592" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="3598" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1114" points="328" swimtime="00:05:15.23" resultid="3764" heatid="4307" lane="6" entrytime="00:04:55.25">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.74" />
                    <SPLIT distance="200" swimtime="00:02:51.18" />
                    <SPLIT distance="300" swimtime="00:04:10.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3676" number="1" />
                    <RELAYPOSITION athleteid="3658" number="2" />
                    <RELAYPOSITION athleteid="3610" number="3" />
                    <RELAYPOSITION athleteid="3664" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1244" points="493" swimtime="00:04:35.37" resultid="3765" heatid="4423" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.30" />
                    <SPLIT distance="200" swimtime="00:02:26.39" />
                    <SPLIT distance="300" swimtime="00:03:32.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3523" number="1" />
                    <RELAYPOSITION athleteid="3547" number="2" />
                    <RELAYPOSITION athleteid="3481" number="3" />
                    <RELAYPOSITION athleteid="3634" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="16830" nation="BRA" region="PR" clubid="1864" swrid="94883" name="Arenna Carvalho Ltda" shortname="Arenna Carvalho">
          <ATHLETES>
            <ATHLETE firstname="Pietro" lastname="Lobo Mussoi" birthdate="2008-07-05" gender="M" nation="BRA" license="398573" swrid="5658061" athleteid="1865" externalid="398573">
              <RESULTS>
                <RESULT eventid="1236" points="464" swimtime="00:00:27.00" resultid="1866" heatid="4417" lane="8" entrytime="00:00:27.57" entrycourse="LCM" />
                <RESULT eventid="1306" points="361" swimtime="00:00:33.05" resultid="1867" heatid="4480" lane="1" entrytime="00:00:33.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="3122" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Helena" lastname="Magalhães Rezende" birthdate="2010-05-29" gender="F" nation="BRA" license="366960" swrid="5588793" athleteid="3135" externalid="366960">
              <RESULTS>
                <RESULT eventid="1080" points="302" swimtime="00:03:25.00" resultid="3136" heatid="4279" lane="5" entrytime="00:03:21.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="329" swimtime="00:00:42.22" resultid="3137" heatid="4357" lane="5" entrytime="00:00:41.84" entrycourse="LCM" />
                <RESULT eventid="1212" points="296" swimtime="00:01:36.15" resultid="3138" heatid="4381" lane="4" entrytime="00:01:30.42" entrycourse="LCM" />
                <RESULT eventid="1250" points="301" swimtime="00:12:03.27" resultid="3139" heatid="4426" lane="3" entrytime="00:11:31.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.98" />
                    <SPLIT distance="200" swimtime="00:02:50.69" />
                    <SPLIT distance="300" swimtime="00:04:22.48" />
                    <SPLIT distance="400" swimtime="00:05:54.57" />
                    <SPLIT distance="500" swimtime="00:07:27.11" />
                    <SPLIT distance="600" swimtime="00:08:59.52" />
                    <SPLIT distance="700" swimtime="00:10:32.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="297" swimtime="00:05:52.42" resultid="3140" heatid="4506" lane="3" entrytime="00:05:46.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.68" />
                    <SPLIT distance="200" swimtime="00:02:47.00" />
                    <SPLIT distance="300" swimtime="00:04:20.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Jacobsen Donati" birthdate="2011-07-14" gender="M" nation="BRA" license="391851" swrid="5615735" athleteid="3189" externalid="391851">
              <RESULTS>
                <RESULT eventid="1072" status="DNS" swimtime="00:00:00.00" resultid="3190" heatid="4273" lane="6" entrytime="00:03:02.40" entrycourse="LCM" />
                <RESULT eventid="1156" points="339" swimtime="00:01:07.16" resultid="3191" heatid="4338" lane="8" entrytime="00:01:08.71" entrycourse="LCM" />
                <RESULT eventid="1236" points="385" swimtime="00:00:28.72" resultid="3192" heatid="4413" lane="5" entrytime="00:00:30.69" entrycourse="LCM" />
                <RESULT eventid="1290" points="271" swimtime="00:02:37.46" resultid="3193" heatid="4460" lane="6" entrytime="00:02:46.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" status="DNS" swimtime="00:00:00.00" resultid="3194" heatid="4528" lane="7" entrytime="00:01:18.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Henrique Ramos" birthdate="2010-02-25" gender="M" nation="BRA" license="406916" swrid="5723024" athleteid="3219" externalid="406916">
              <RESULTS>
                <RESULT eventid="1156" points="269" swimtime="00:01:12.53" resultid="3220" heatid="4336" lane="7" entrytime="00:01:13.74" entrycourse="LCM" />
                <RESULT eventid="1236" points="280" swimtime="00:00:31.96" resultid="3221" heatid="4409" lane="7" />
                <RESULT eventid="1290" points="259" swimtime="00:02:39.99" resultid="3222" heatid="4460" lane="5" entrytime="00:02:43.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1306" points="193" swimtime="00:00:40.69" resultid="3223" heatid="4477" lane="7" />
                <RESULT eventid="1374" status="DSQ" swimtime="00:01:29.08" resultid="3224" heatid="4527" lane="8" entrytime="00:01:29.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rodrigo" lastname="Zanatta Duda" birthdate="2011-09-12" gender="M" nation="BRA" license="406917" swrid="5717307" athleteid="3225" externalid="406917">
              <RESULTS>
                <RESULT eventid="1072" points="196" swimtime="00:03:12.59" resultid="3226" heatid="4273" lane="7" entrytime="00:03:10.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="179" swimtime="00:01:23.08" resultid="3227" heatid="4334" lane="7" entrytime="00:01:29.58" entrycourse="LCM" />
                <RESULT eventid="1188" points="167" swimtime="00:00:47.12" resultid="3228" heatid="4363" lane="8" />
                <RESULT eventid="1306" points="189" swimtime="00:00:41.02" resultid="3229" heatid="4477" lane="5" />
                <RESULT eventid="1374" points="188" swimtime="00:01:29.93" resultid="3230" heatid="4527" lane="1" entrytime="00:01:29.57" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Ribeiro Melo" birthdate="2011-07-01" gender="F" nation="BRA" license="390923" swrid="5602577" athleteid="3207" externalid="390923">
              <RESULTS>
                <RESULT eventid="1148" points="367" swimtime="00:01:12.20" resultid="3208" heatid="4325" lane="8" entrytime="00:01:11.49" entrycourse="LCM" />
                <RESULT eventid="1228" points="429" swimtime="00:00:31.29" resultid="3209" heatid="4401" lane="2" entrytime="00:00:32.42" entrycourse="LCM" />
                <RESULT eventid="1212" points="272" swimtime="00:01:38.88" resultid="3210" heatid="4379" lane="4" entrytime="00:01:49.17" entrycourse="LCM" />
                <RESULT eventid="1282" points="343" swimtime="00:02:41.08" resultid="3211" heatid="4454" lane="1" entrytime="00:02:34.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="285" swimtime="00:01:27.04" resultid="3212" heatid="4520" lane="7" entrytime="00:01:26.41" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aline" lastname="Hirano" birthdate="2007-11-13" gender="F" nation="BRA" license="358898" swrid="5622283" athleteid="3213" externalid="358898">
              <RESULTS>
                <RESULT eventid="1116" points="379" swimtime="00:21:10.98" resultid="3214" heatid="4308" lane="7" entrytime="00:22:41.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                    <SPLIT distance="200" swimtime="00:02:36.59" />
                    <SPLIT distance="300" swimtime="00:04:00.56" />
                    <SPLIT distance="400" swimtime="00:05:26.04" />
                    <SPLIT distance="500" swimtime="00:06:51.79" />
                    <SPLIT distance="600" swimtime="00:08:16.66" />
                    <SPLIT distance="700" swimtime="00:09:43.59" />
                    <SPLIT distance="800" swimtime="00:11:11.65" />
                    <SPLIT distance="900" swimtime="00:12:40.19" />
                    <SPLIT distance="1000" swimtime="00:14:10.71" />
                    <SPLIT distance="1100" swimtime="00:15:35.48" />
                    <SPLIT distance="1200" swimtime="00:16:59.84" />
                    <SPLIT distance="1300" swimtime="00:18:24.81" />
                    <SPLIT distance="1400" swimtime="00:19:51.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="283" swimtime="00:01:37.64" resultid="3215" heatid="4377" lane="5" />
                <RESULT eventid="1250" points="406" swimtime="00:10:54.24" resultid="3216" heatid="4427" lane="1" entrytime="00:11:03.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.26" />
                    <SPLIT distance="200" swimtime="00:02:37.84" />
                    <SPLIT distance="300" swimtime="00:04:01.13" />
                    <SPLIT distance="400" swimtime="00:05:23.95" />
                    <SPLIT distance="500" swimtime="00:06:47.40" />
                    <SPLIT distance="600" swimtime="00:08:11.69" />
                    <SPLIT distance="700" swimtime="00:09:35.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" points="369" swimtime="00:02:55.73" resultid="3217" heatid="4436" lane="4" entrytime="00:03:02.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="369" swimtime="00:01:19.89" resultid="3218" heatid="4521" lane="6" entrytime="00:01:22.87" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Berto" birthdate="2008-10-22" gender="M" nation="BRA" license="378342" swrid="5312223" athleteid="3141" externalid="378342">
              <RESULTS>
                <RESULT eventid="1088" points="398" swimtime="00:02:50.55" resultid="3142" heatid="4286" lane="4" entrytime="00:02:52.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="335" swimtime="00:01:07.46" resultid="3143" heatid="4337" lane="8" entrytime="00:01:11.13" entrycourse="LCM" />
                <RESULT eventid="1188" points="346" swimtime="00:00:36.95" resultid="3144" heatid="4366" lane="1" entrytime="00:00:36.67" entrycourse="LCM" />
                <RESULT eventid="1220" points="369" swimtime="00:01:19.30" resultid="3145" heatid="4391" lane="3" entrytime="00:01:20.81" entrycourse="LCM" />
                <RESULT eventid="1274" points="328" swimtime="00:02:45.24" resultid="3146" heatid="4441" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Traci Rodrigues" birthdate="2011-03-06" gender="M" nation="BRA" license="406927" swrid="5718893" athleteid="3231" externalid="406927">
              <RESULTS>
                <RESULT eventid="1156" points="176" swimtime="00:01:23.49" resultid="3232" heatid="4331" lane="3" />
                <RESULT eventid="1188" points="168" swimtime="00:00:46.94" resultid="3233" heatid="4361" lane="2" />
                <RESULT eventid="1220" points="135" swimtime="00:01:50.82" resultid="3234" heatid="4385" lane="5" />
                <RESULT eventid="1236" points="191" swimtime="00:00:36.29" resultid="3235" heatid="4410" lane="6" />
                <RESULT eventid="1306" points="131" swimtime="00:00:46.27" resultid="3236" heatid="4478" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Pazinato" birthdate="2011-01-05" gender="M" nation="BRA" license="368149" swrid="5603889" athleteid="3171" externalid="368149">
              <RESULTS>
                <RESULT eventid="1072" points="252" swimtime="00:02:57.14" resultid="3172" heatid="4272" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="337" swimtime="00:01:07.28" resultid="3173" heatid="4337" lane="7" entrytime="00:01:10.36" entrycourse="LCM" />
                <RESULT eventid="1236" points="308" swimtime="00:00:30.94" resultid="3174" heatid="4412" lane="4" entrytime="00:00:31.43" entrycourse="LCM" />
                <RESULT eventid="1290" points="287" swimtime="00:02:34.46" resultid="3175" heatid="4461" lane="4" entrytime="00:02:36.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="265" swimtime="00:01:20.33" resultid="3176" heatid="4526" lane="4" entrytime="00:01:29.89" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theodoro" lastname="Marques Serra" birthdate="2009-11-24" gender="M" nation="BRA" license="370661" swrid="5603870" athleteid="3177" externalid="370661">
              <RESULTS>
                <RESULT eventid="1072" points="339" swimtime="00:02:40.45" resultid="3178" heatid="4274" lane="1" entrytime="00:02:47.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="426" swimtime="00:01:02.25" resultid="3179" heatid="4333" lane="7" />
                <RESULT eventid="1290" points="390" swimtime="00:02:19.59" resultid="3180" heatid="4463" lane="8" entrytime="00:02:27.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1306" points="353" swimtime="00:00:33.32" resultid="3181" heatid="4479" lane="5" entrytime="00:00:34.13" entrycourse="LCM" />
                <RESULT eventid="1374" points="373" swimtime="00:01:11.65" resultid="3182" heatid="4528" lane="4" entrytime="00:01:14.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Braga" birthdate="2010-05-07" gender="M" nation="BRA" license="378345" swrid="5343953" athleteid="3159" externalid="378345">
              <RESULTS>
                <RESULT eventid="1088" points="396" swimtime="00:02:50.77" resultid="3160" heatid="4286" lane="3" entrytime="00:02:53.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="378" swimtime="00:00:35.86" resultid="3161" heatid="4366" lane="7" entrytime="00:00:36.57" entrycourse="LCM" />
                <RESULT eventid="1220" points="409" swimtime="00:01:16.60" resultid="3162" heatid="4392" lane="8" entrytime="00:01:20.41" entrycourse="LCM" />
                <RESULT eventid="1274" points="326" swimtime="00:02:45.50" resultid="3163" heatid="4442" lane="4" entrytime="00:03:16.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="300" swimtime="00:05:28.60" resultid="3164" heatid="4511" lane="5" entrytime="00:05:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.98" />
                    <SPLIT distance="200" swimtime="00:02:38.47" />
                    <SPLIT distance="300" swimtime="00:04:04.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Sales" birthdate="2011-02-28" gender="F" nation="BRA" license="374103" swrid="5616410" athleteid="3165" externalid="374103">
              <RESULTS>
                <RESULT eventid="1080" points="321" swimtime="00:03:20.71" resultid="3166" heatid="4278" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="381" swimtime="00:01:11.28" resultid="3167" heatid="4322" lane="3" entrytime="00:01:15.99" entrycourse="LCM" />
                <RESULT eventid="1212" points="310" swimtime="00:01:34.71" resultid="3168" heatid="4912" lane="4" entrytime="00:01:33.07" entrycourse="LCM" />
                <RESULT eventid="1282" points="334" swimtime="00:02:42.61" resultid="3169" heatid="4977" lane="3" entrytime="00:02:42.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="373" swimtime="00:01:17.05" resultid="3170" heatid="4493" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Ferreira Rais" birthdate="2007-07-04" gender="M" nation="BRA" license="398656" swrid="5697227" athleteid="3201" externalid="398656">
              <RESULTS>
                <RESULT eventid="1104" points="268" swimtime="00:00:34.51" resultid="3202" heatid="4295" lane="7" />
                <RESULT eventid="1156" points="343" swimtime="00:01:06.94" resultid="3203" heatid="4339" lane="2" entrytime="00:01:06.94" entrycourse="LCM" />
                <RESULT eventid="1236" points="373" swimtime="00:00:29.03" resultid="3204" heatid="4406" lane="6" />
                <RESULT eventid="1290" points="219" swimtime="00:02:49.08" resultid="3205" heatid="4461" lane="1" entrytime="00:02:41.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1306" points="217" swimtime="00:00:39.16" resultid="3206" heatid="4478" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Guilherme Ballatka" birthdate="2007-06-24" gender="M" nation="BRA" license="398616" swrid="5697228" athleteid="3195" externalid="398616">
              <RESULTS>
                <RESULT eventid="1156" points="410" swimtime="00:01:03.07" resultid="3196" heatid="4341" lane="7" entrytime="00:01:05.35" entrycourse="LCM" />
                <RESULT eventid="1188" points="280" swimtime="00:00:39.62" resultid="3197" heatid="4363" lane="6" />
                <RESULT eventid="1236" points="443" swimtime="00:00:27.41" resultid="3198" heatid="4406" lane="8" />
                <RESULT eventid="1306" points="399" swimtime="00:00:31.97" resultid="3199" heatid="4476" lane="2" />
                <RESULT eventid="1374" points="303" swimtime="00:01:16.79" resultid="3200" heatid="4529" lane="7" entrytime="00:01:13.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Kenji Yamaguchi" birthdate="2011-08-25" gender="M" nation="BRA" license="385708" swrid="5603862" athleteid="3183" externalid="385708">
              <RESULTS>
                <RESULT eventid="1104" points="248" swimtime="00:00:35.41" resultid="3184" heatid="4298" lane="7" entrytime="00:00:39.20" entrycourse="LCM" />
                <RESULT eventid="1172" points="171" swimtime="00:03:18.70" resultid="3185" heatid="4352" lane="8" entrytime="00:03:55.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="224" swimtime="00:01:33.55" resultid="3186" heatid="4387" lane="8" />
                <RESULT eventid="1274" points="258" swimtime="00:02:58.88" resultid="3187" heatid="4442" lane="5" entrytime="00:03:18.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="210" swimtime="00:01:23.15" resultid="3188" heatid="4499" lane="7" entrytime="00:01:47.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benicio" lastname="Garcia" birthdate="2011-09-09" gender="M" nation="BRA" license="378347" swrid="5603842" athleteid="3123" externalid="378347">
              <RESULTS>
                <RESULT eventid="1072" points="234" swimtime="00:03:01.46" resultid="3124" heatid="4273" lane="2" entrytime="00:03:09.17" entrycourse="LCM" />
                <RESULT eventid="1156" points="268" swimtime="00:01:12.60" resultid="3125" heatid="4335" lane="4" entrytime="00:01:15.43" entrycourse="LCM" />
                <RESULT eventid="1306" points="242" swimtime="00:00:37.78" resultid="3126" heatid="4479" lane="1" entrytime="00:00:37.58" entrycourse="LCM" />
                <RESULT eventid="1274" points="210" swimtime="00:03:11.71" resultid="3127" heatid="4442" lane="6" entrytime="00:03:21.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="271" swimtime="00:01:19.68" resultid="3128" heatid="4527" lane="6" entrytime="00:01:23.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Camillo Sabim" birthdate="2010-08-02" gender="F" nation="BRA" license="406931" swrid="5723021" athleteid="3237" externalid="406931">
              <RESULTS>
                <RESULT eventid="1148" points="247" swimtime="00:01:22.40" resultid="3238" heatid="4321" lane="2" entrytime="00:01:25.08" entrycourse="LCM" />
                <RESULT eventid="1180" points="297" swimtime="00:00:43.67" resultid="3239" heatid="4355" lane="7" />
                <RESULT eventid="1228" points="296" swimtime="00:00:35.39" resultid="3240" heatid="4396" lane="3" />
                <RESULT eventid="1298" points="277" swimtime="00:00:41.20" resultid="3241" heatid="4470" lane="5" />
                <RESULT eventid="1366" points="245" swimtime="00:01:31.53" resultid="3242" heatid="4518" lane="6" entrytime="00:01:38.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Ortega" birthdate="1999-08-05" gender="M" nation="BRA" license="383118" swrid="5603852" athleteid="3129" externalid="383118">
              <RESULTS>
                <RESULT eventid="1072" points="363" swimtime="00:02:36.88" resultid="3130" heatid="4274" lane="4" entrytime="00:02:39.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="425" swimtime="00:00:27.79" resultid="3131" heatid="4406" lane="1" />
                <RESULT eventid="1290" points="315" swimtime="00:02:29.82" resultid="3132" heatid="4463" lane="3" entrytime="00:02:26.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1306" points="390" swimtime="00:00:32.22" resultid="3133" heatid="4480" lane="5" entrytime="00:00:32.13" entrycourse="LCM" />
                <RESULT eventid="1374" points="390" swimtime="00:01:10.61" resultid="3134" heatid="4530" lane="1" entrytime="00:01:11.59" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Silveira De Almeida" birthdate="2008-07-08" gender="M" nation="BRA" license="368152" swrid="5603912" athleteid="3147" externalid="368152">
              <RESULTS>
                <RESULT eventid="1104" points="516" swimtime="00:00:27.76" resultid="3148" heatid="4302" lane="2" entrytime="00:00:28.79" entrycourse="LCM" />
                <RESULT eventid="1172" points="378" swimtime="00:02:32.58" resultid="3149" heatid="4354" lane="8" entrytime="00:02:20.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="411" swimtime="00:00:28.12" resultid="3150" heatid="4417" lane="7" entrytime="00:00:27.49" entrycourse="LCM" />
                <RESULT eventid="1274" points="432" swimtime="00:02:30.72" resultid="3151" heatid="4445" lane="6" entrytime="00:02:41.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" status="DSQ" swimtime="00:01:01.70" resultid="3152" heatid="4504" lane="8" entrytime="00:01:02.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jennifer" lastname="De Abreu" birthdate="2009-11-07" gender="F" nation="BRA" license="356212" swrid="5600144" athleteid="3153" externalid="356212">
              <RESULTS>
                <RESULT eventid="1148" points="500" swimtime="00:01:05.15" resultid="3154" heatid="4329" lane="8" entrytime="00:01:05.23" entrycourse="LCM" />
                <RESULT eventid="1228" points="454" swimtime="00:00:30.71" resultid="3155" heatid="4404" lane="1" entrytime="00:00:30.20" entrycourse="LCM" />
                <RESULT eventid="1212" points="375" swimtime="00:01:28.91" resultid="3156" heatid="4382" lane="6" entrytime="00:01:28.23" entrycourse="LCM" />
                <RESULT eventid="1266" points="444" swimtime="00:02:45.28" resultid="3157" heatid="4438" lane="7" entrytime="00:02:53.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="396" swimtime="00:01:15.52" resultid="3158" heatid="4496" lane="3" entrytime="00:01:17.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1204" points="289" swimtime="00:10:32.54" resultid="3244" heatid="4373" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.24" />
                    <SPLIT distance="200" swimtime="00:02:37.98" />
                    <SPLIT distance="300" swimtime="00:03:51.15" />
                    <SPLIT distance="400" swimtime="00:05:10.85" />
                    <SPLIT distance="500" swimtime="00:06:28.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3171" number="1" />
                    <RELAYPOSITION athleteid="3159" number="2" />
                    <RELAYPOSITION athleteid="3123" number="3" />
                    <RELAYPOSITION athleteid="3189" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1324" points="210" swimtime="00:05:47.85" resultid="3245" heatid="4488" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.37" />
                    <SPLIT distance="200" swimtime="00:03:07.62" />
                    <SPLIT distance="300" swimtime="00:04:30.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3189" number="1" />
                    <RELAYPOSITION athleteid="3171" number="2" />
                    <RELAYPOSITION athleteid="3183" number="3" />
                    <RELAYPOSITION athleteid="3123" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1392" points="240" swimtime="00:05:02.73" resultid="3247" heatid="4539" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.69" />
                    <SPLIT distance="200" swimtime="00:02:31.39" />
                    <SPLIT distance="300" swimtime="00:03:48.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3171" number="1" />
                    <RELAYPOSITION athleteid="3225" number="2" />
                    <RELAYPOSITION athleteid="3123" number="3" />
                    <RELAYPOSITION athleteid="3183" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1326" points="210" swimtime="00:05:47.71" resultid="3246" heatid="4489" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.95" />
                    <SPLIT distance="300" swimtime="00:04:35.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3225" number="1" />
                    <RELAYPOSITION athleteid="3231" number="2" />
                    <RELAYPOSITION athleteid="3159" number="3" />
                    <RELAYPOSITION athleteid="3219" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1394" status="WDR" swimtime="00:00:00.00" resultid="3248" heatid="4540" lane="7" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1384" points="310" swimtime="00:05:07.10" resultid="3243" heatid="4535" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.19" />
                    <SPLIT distance="200" swimtime="00:02:38.54" />
                    <SPLIT distance="300" swimtime="00:03:54.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3165" number="1" />
                    <RELAYPOSITION athleteid="3237" number="2" />
                    <RELAYPOSITION athleteid="3135" number="3" />
                    <RELAYPOSITION athleteid="3207" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1112" points="288" swimtime="00:05:29.10" resultid="3249" heatid="4305" lane="4">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:02:51.70" />
                    <SPLIT distance="300" swimtime="00:04:15.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3189" number="1" />
                    <RELAYPOSITION athleteid="3165" number="2" />
                    <RELAYPOSITION athleteid="3183" number="3" />
                    <RELAYPOSITION athleteid="3207" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1114" points="248" swimtime="00:05:45.91" resultid="3250" heatid="4307" lane="1">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:03:05.98" />
                    <SPLIT distance="300" swimtime="00:04:23.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3219" number="1" />
                    <RELAYPOSITION athleteid="3135" number="2" />
                    <RELAYPOSITION athleteid="3159" number="3" />
                    <RELAYPOSITION athleteid="3237" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="15981" nation="BRA" region="PR" clubid="1403" swrid="93783" name="Quinto Nado" shortname="5º Nado">
          <ATHLETES>
            <ATHLETE firstname="Gabriela" lastname="Poletti Veiga" birthdate="2010-10-01" gender="F" nation="BRA" license="376951" swrid="5603895" athleteid="1427" externalid="376951">
              <RESULTS>
                <RESULT eventid="1064" points="403" swimtime="00:02:46.62" resultid="1428" heatid="4266" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="491" swimtime="00:01:05.51" resultid="1429" heatid="4327" lane="7" entrytime="00:01:08.14" entrycourse="LCM" />
                <RESULT eventid="1228" points="478" swimtime="00:00:30.19" resultid="1430" heatid="4402" lane="3" entrytime="00:00:31.10" entrycourse="LCM" />
                <RESULT eventid="1334" points="304" swimtime="00:01:22.45" resultid="1431" heatid="4493" lane="3" />
                <RESULT eventid="1366" points="402" swimtime="00:01:17.67" resultid="1432" heatid="4522" lane="6" entrytime="00:01:19.19" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Takemura Couto" birthdate="2010-02-08" gender="F" nation="BRA" license="376950" swrid="5603919" athleteid="1433" externalid="376950">
              <RESULTS>
                <RESULT eventid="1064" points="364" swimtime="00:02:52.38" resultid="1434" heatid="4269" lane="7" entrytime="00:02:58.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="503" swimtime="00:01:05.02" resultid="1435" heatid="4324" lane="6" entrytime="00:01:12.18" entrycourse="LCM" />
                <RESULT eventid="1228" points="506" swimtime="00:00:29.61" resultid="1436" heatid="4403" lane="7" entrytime="00:00:30.69" entrycourse="LCM" />
                <RESULT eventid="1282" points="384" swimtime="00:02:35.18" resultid="1437" heatid="4449" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" points="338" swimtime="00:03:00.98" resultid="1438" heatid="4437" lane="7" entrytime="00:03:01.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Bordini Zocco" birthdate="2008-08-04" gender="F" nation="BRA" license="385677" swrid="5332871" athleteid="1415" externalid="385677">
              <RESULTS>
                <RESULT eventid="1064" points="327" swimtime="00:02:58.68" resultid="1416" heatid="4266" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="401" swimtime="00:01:10.10" resultid="1417" heatid="4324" lane="7" entrytime="00:01:13.20" entrycourse="LCM" />
                <RESULT eventid="1212" points="319" swimtime="00:01:33.80" resultid="1418" heatid="4381" lane="8" entrytime="00:01:35.24" entrycourse="LCM" />
                <RESULT eventid="1266" points="344" swimtime="00:02:59.87" resultid="1419" heatid="4437" lane="5" entrytime="00:02:59.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="343" swimtime="00:01:21.83" resultid="1420" heatid="4521" lane="7" entrytime="00:01:22.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Kikuchi Fujii" birthdate="2007-01-04" gender="M" nation="BRA" license="297805" swrid="5603863" athleteid="1404" externalid="297805">
              <RESULTS>
                <RESULT eventid="1088" points="624" swimtime="00:02:26.84" resultid="1405" heatid="4289" lane="2" entrytime="00:02:24.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="438" swimtime="00:02:25.21" resultid="1406" heatid="4353" lane="6" entrytime="00:02:32.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="596" swimtime="00:01:07.58" resultid="1407" heatid="4395" lane="1" entrytime="00:01:06.44" entrycourse="LCM" />
                <RESULT eventid="1274" points="594" swimtime="00:02:15.59" resultid="1408" heatid="4448" lane="6" entrytime="00:02:14.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="606" swimtime="00:00:58.41" resultid="1409" heatid="4498" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Betina" lastname="Tramontini Queiroz" birthdate="2007-09-11" gender="F" nation="BRA" license="357155" swrid="5658063" athleteid="1421" externalid="357155">
              <RESULTS>
                <RESULT eventid="1116" points="491" swimtime="00:19:26.49" resultid="1422" heatid="4309" lane="6" entrytime="00:19:19.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.91" />
                    <SPLIT distance="200" swimtime="00:02:30.32" />
                    <SPLIT distance="300" swimtime="00:03:49.12" />
                    <SPLIT distance="400" swimtime="00:05:07.81" />
                    <SPLIT distance="500" swimtime="00:06:26.11" />
                    <SPLIT distance="600" swimtime="00:07:44.36" />
                    <SPLIT distance="700" swimtime="00:09:02.27" />
                    <SPLIT distance="800" swimtime="00:10:20.88" />
                    <SPLIT distance="900" swimtime="00:11:39.00" />
                    <SPLIT distance="1000" swimtime="00:12:57.62" />
                    <SPLIT distance="1100" swimtime="00:14:16.06" />
                    <SPLIT distance="1200" swimtime="00:15:34.00" />
                    <SPLIT distance="1300" swimtime="00:16:51.10" />
                    <SPLIT distance="1400" swimtime="00:18:09.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="559" swimtime="00:01:02.77" resultid="1423" heatid="4329" lane="2" entrytime="00:01:04.64" entrycourse="LCM" />
                <RESULT eventid="1250" points="479" swimtime="00:10:19.48" resultid="1424" heatid="4428" lane="2" entrytime="00:10:03.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.30" />
                    <SPLIT distance="200" swimtime="00:02:30.36" />
                    <SPLIT distance="300" swimtime="00:03:49.83" />
                    <SPLIT distance="400" swimtime="00:05:09.38" />
                    <SPLIT distance="500" swimtime="00:06:27.86" />
                    <SPLIT distance="600" swimtime="00:07:46.13" />
                    <SPLIT distance="700" swimtime="00:09:03.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="554" swimtime="00:02:17.39" resultid="1425" heatid="4456" lane="5" entrytime="00:02:18.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="482" swimtime="00:05:00.19" resultid="1426" heatid="4509" lane="4" entrytime="00:04:54.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.94" />
                    <SPLIT distance="200" swimtime="00:02:26.20" />
                    <SPLIT distance="300" swimtime="00:03:43.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Dequech Queiroz" birthdate="2004-05-20" gender="M" nation="BRA" license="318401" athleteid="1410" externalid="318401">
              <RESULTS>
                <RESULT eventid="1104" points="566" swimtime="00:00:26.92" resultid="1411" heatid="4303" lane="5" entrytime="00:00:27.62" entrycourse="LCM" />
                <RESULT eventid="1156" points="588" swimtime="00:00:55.92" resultid="1412" heatid="4331" lane="4" />
                <RESULT eventid="1236" points="606" swimtime="00:00:24.70" resultid="1413" heatid="4421" lane="3" entrytime="00:00:24.75" entrycourse="LCM" />
                <RESULT eventid="1342" points="490" swimtime="00:01:02.69" resultid="1414" heatid="4498" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Gomes" birthdate="2011-12-03" gender="F" nation="BRA" license="382051" swrid="5603846" athleteid="1439" externalid="382051">
              <RESULTS>
                <RESULT eventid="1228" points="214" swimtime="00:00:39.46" resultid="1440" heatid="4397" lane="8" />
                <RESULT eventid="1212" points="111" swimtime="00:02:13.32" resultid="1441" heatid="4378" lane="3" />
                <RESULT eventid="1282" points="240" swimtime="00:03:01.42" resultid="1442" heatid="4450" lane="2" />
                <RESULT eventid="1298" points="210" swimtime="00:00:45.14" resultid="1443" heatid="4471" lane="2" />
                <RESULT eventid="1366" status="DSQ" swimtime="00:01:40.14" resultid="1444" heatid="4517" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Fernanda Romero" birthdate="2007-04-18" gender="F" nation="BRA" license="404750" swrid="4828153" athleteid="1445" externalid="404750">
              <RESULTS>
                <RESULT eventid="1164" points="408" swimtime="00:02:44.23" resultid="1446" heatid="4350" lane="6" entrytime="00:02:48.88" entrycourse="LCM" />
                <RESULT eventid="1180" points="515" swimtime="00:00:36.37" resultid="1447" heatid="4355" lane="2" />
                <RESULT eventid="1212" status="DSQ" swimtime="00:01:23.80" resultid="1448" heatid="4383" lane="2" entrytime="00:01:24.36" entrycourse="LCM" />
                <RESULT eventid="1266" points="498" swimtime="00:02:39.07" resultid="1449" heatid="4439" lane="2" entrytime="00:02:38.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="414" swimtime="00:01:14.39" resultid="1450" heatid="4493" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="5º NADO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1248" points="535" swimtime="00:04:27.90" resultid="1451" heatid="4425" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.69" />
                    <SPLIT distance="200" swimtime="00:02:21.78" />
                    <SPLIT distance="300" swimtime="00:03:24.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1445" number="1" />
                    <RELAYPOSITION athleteid="1404" number="2" />
                    <RELAYPOSITION athleteid="1410" number="3" />
                    <RELAYPOSITION athleteid="1421" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="263" nation="BRA" region="PR" clubid="2444" swrid="75436" name="Clube Curitibano" shortname="Curitibano">
          <ATHLETES>
            <ATHLETE firstname="Alice" lastname="Jardim" birthdate="2010-03-23" gender="F" nation="BRA" license="368006" swrid="5600192" athleteid="2839" externalid="368006">
              <RESULTS>
                <RESULT eventid="1148" points="379" swimtime="00:01:11.40" resultid="2840" heatid="4326" lane="7" entrytime="00:01:09.93" entrycourse="LCM" />
                <RESULT eventid="1228" points="381" swimtime="00:00:32.55" resultid="2841" heatid="4401" lane="5" entrytime="00:00:31.90" entrycourse="LCM" />
                <RESULT eventid="1282" points="343" swimtime="00:02:41.08" resultid="2842" heatid="4454" lane="3" entrytime="00:02:31.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" points="320" swimtime="00:03:04.26" resultid="2843" heatid="4436" lane="3" entrytime="00:03:06.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="311" swimtime="00:05:47.40" resultid="2844" heatid="4508" lane="2" entrytime="00:05:32.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.94" />
                    <SPLIT distance="200" swimtime="00:02:49.58" />
                    <SPLIT distance="300" swimtime="00:04:21.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo" lastname="Gabriel Nascimento" birthdate="2008-11-14" gender="M" nation="BRA" license="348028" swrid="5600171" athleteid="2940" externalid="348028">
              <RESULTS>
                <RESULT eventid="1104" points="499" swimtime="00:00:28.07" resultid="2941" heatid="4302" lane="1" entrytime="00:00:29.09" entrycourse="LCM" />
                <RESULT eventid="1156" points="478" swimtime="00:00:59.91" resultid="2942" heatid="4344" lane="4" entrytime="00:00:59.61" entrycourse="LCM" />
                <RESULT eventid="1236" points="470" swimtime="00:00:26.89" resultid="2943" heatid="4419" lane="8" entrytime="00:00:26.68" entrycourse="LCM" />
                <RESULT eventid="1342" points="448" swimtime="00:01:04.62" resultid="2944" heatid="4503" lane="6" entrytime="00:01:04.11" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Fontes Bonardi" birthdate="2008-10-26" gender="M" nation="BRA" license="307662" swrid="5600164" athleteid="2478" externalid="307662">
              <RESULTS>
                <RESULT eventid="1088" points="537" swimtime="00:02:34.29" resultid="2479" heatid="4289" lane="8" entrytime="00:02:31.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="535" swimtime="00:04:58.65" resultid="2480" heatid="4318" lane="6" entrytime="00:04:54.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.74" />
                    <SPLIT distance="200" swimtime="00:02:27.13" />
                    <SPLIT distance="300" swimtime="00:03:51.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="506" swimtime="00:01:11.36" resultid="2481" heatid="4394" lane="2" entrytime="00:01:10.01" entrycourse="LCM" />
                <RESULT eventid="1274" points="565" swimtime="00:02:17.82" resultid="2482" heatid="4448" lane="8" entrytime="00:02:18.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="454" swimtime="00:01:07.09" resultid="2483" heatid="4531" lane="4" entrytime="00:01:07.89" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Rocha Silva" birthdate="2007-10-10" gender="M" nation="BRA" license="372280" swrid="5717294" athleteid="2547" externalid="372280">
              <RESULTS>
                <RESULT eventid="1104" points="605" swimtime="00:00:26.33" resultid="2548" heatid="4302" lane="8" entrytime="00:00:29.21" entrycourse="LCM" />
                <RESULT eventid="1156" points="774" swimtime="00:00:51.02" resultid="2549" heatid="4348" lane="4" entrytime="00:00:51.08" entrycourse="LCM" />
                <RESULT eventid="1236" points="678" swimtime="00:00:23.80" resultid="2550" heatid="4422" lane="4" entrytime="00:00:23.27" entrycourse="LCM" />
                <RESULT eventid="1290" points="753" swimtime="00:01:52.10" resultid="2551" heatid="4469" lane="3" entrytime="00:01:54.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" status="DNS" swimtime="00:00:00.00" resultid="2552" heatid="4516" lane="7" entrytime="00:04:31.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietra" lastname="Ruschel Carvalho" birthdate="2009-03-21" gender="F" nation="BRA" license="324999" swrid="5600250" athleteid="2460" externalid="324999">
              <RESULTS>
                <RESULT eventid="1096" points="452" swimtime="00:00:31.81" resultid="2461" heatid="4294" lane="6" entrytime="00:00:31.15" entrycourse="LCM" />
                <RESULT eventid="1148" points="616" swimtime="00:01:00.76" resultid="2462" heatid="4330" lane="2" entrytime="00:01:01.08" entrycourse="LCM" />
                <RESULT eventid="1228" points="626" swimtime="00:00:27.59" resultid="2463" heatid="4405" lane="4" entrytime="00:00:27.34" entrycourse="LCM" />
                <RESULT eventid="1282" points="597" swimtime="00:02:14.01" resultid="2464" heatid="4457" lane="7" entrytime="00:02:13.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo" lastname="De Hamerschmidt" birthdate="2009-04-15" gender="M" nation="BRA" license="339069" swrid="5600147" athleteid="2647" externalid="339069">
              <RESULTS>
                <RESULT eventid="1104" status="DNS" swimtime="00:00:00.00" resultid="2648" heatid="4301" lane="8" entrytime="00:00:30.30" entrycourse="LCM" />
                <RESULT eventid="1172" status="DNS" swimtime="00:00:00.00" resultid="2649" heatid="4353" lane="7" entrytime="00:02:37.19" entrycourse="LCM" />
                <RESULT eventid="1236" status="DNS" swimtime="00:00:00.00" resultid="2650" heatid="4416" lane="6" entrytime="00:00:28.00" entrycourse="LCM" />
                <RESULT eventid="1342" status="DNS" swimtime="00:00:00.00" resultid="2651" heatid="4502" lane="3" entrytime="00:01:06.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Fontana Moraes" birthdate="2006-08-17" gender="M" nation="BRA" license="296593" swrid="5600163" athleteid="2564" externalid="296593">
              <RESULTS>
                <RESULT eventid="1124" points="290" swimtime="00:11:22.32" resultid="2565" heatid="4310" lane="3" entrytime="00:11:20.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.31" />
                    <SPLIT distance="200" swimtime="00:02:45.20" />
                    <SPLIT distance="300" swimtime="00:04:13.08" />
                    <SPLIT distance="400" swimtime="00:05:40.80" />
                    <SPLIT distance="500" swimtime="00:07:08.55" />
                    <SPLIT distance="600" swimtime="00:08:35.69" />
                    <SPLIT distance="700" swimtime="00:10:00.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="294" swimtime="00:01:10.44" resultid="2566" heatid="4340" lane="8" entrytime="00:01:06.57" entrycourse="LCM" />
                <RESULT eventid="1236" points="323" swimtime="00:00:30.47" resultid="2567" heatid="4414" lane="3" entrytime="00:00:30.16" entrycourse="LCM" />
                <RESULT eventid="1290" points="275" swimtime="00:02:36.74" resultid="2568" heatid="4462" lane="3" entrytime="00:02:31.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="281" swimtime="00:05:35.90" resultid="2569" heatid="4513" lane="1" entrytime="00:05:23.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.79" />
                    <SPLIT distance="200" swimtime="00:02:44.18" />
                    <SPLIT distance="300" swimtime="00:04:11.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pablo" lastname="Souza Tavares" birthdate="2006-05-03" gender="M" nation="BRA" license="331982" swrid="5600261" athleteid="2465" externalid="331982">
              <RESULTS>
                <RESULT eventid="1072" points="608" swimtime="00:02:12.04" resultid="2466" heatid="4277" lane="5" entrytime="00:02:11.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="645" swimtime="00:00:59.72" resultid="2467" heatid="4533" lane="5" entrytime="00:00:59.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Correa Nascimento" birthdate="2009-01-19" gender="M" nation="BRA" license="342235" swrid="5600140" athleteid="2605" externalid="342235">
              <RESULTS>
                <RESULT eventid="1104" points="386" swimtime="00:00:30.57" resultid="2606" heatid="4297" lane="5" />
                <RESULT eventid="1156" points="485" swimtime="00:00:59.63" resultid="2607" heatid="4345" lane="5" entrytime="00:00:58.77" entrycourse="LCM" />
                <RESULT eventid="1220" points="370" swimtime="00:01:19.23" resultid="2608" heatid="4386" lane="2" />
                <RESULT eventid="1290" points="428" swimtime="00:02:15.28" resultid="2609" heatid="4465" lane="5" entrytime="00:02:15.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="De Krinski" birthdate="2007-07-20" gender="M" nation="BRA" license="334494" swrid="5600148" athleteid="2987" externalid="334494">
              <RESULTS>
                <RESULT eventid="1072" points="513" swimtime="00:02:19.75" resultid="2988" heatid="4277" lane="8" entrytime="00:02:19.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="575" swimtime="00:00:56.34" resultid="2989" heatid="4346" lane="5" entrytime="00:00:57.10" entrycourse="LCM" />
                <RESULT eventid="1306" points="543" swimtime="00:00:28.86" resultid="2990" heatid="4482" lane="3" entrytime="00:00:28.56" entrycourse="LCM" />
                <RESULT eventid="1374" points="531" swimtime="00:01:03.72" resultid="2991" heatid="4533" lane="2" entrytime="00:01:01.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Schiavon" birthdate="2010-05-03" gender="M" nation="BRA" license="356354" swrid="5600256" athleteid="2706" externalid="356354">
              <RESULTS>
                <RESULT eventid="1124" points="457" swimtime="00:09:46.82" resultid="2707" heatid="4312" lane="4" entrytime="00:09:37.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.96" />
                    <SPLIT distance="200" swimtime="00:02:18.86" />
                    <SPLIT distance="300" swimtime="00:03:32.03" />
                    <SPLIT distance="400" swimtime="00:04:46.85" />
                    <SPLIT distance="500" swimtime="00:06:02.11" />
                    <SPLIT distance="600" swimtime="00:07:17.56" />
                    <SPLIT distance="700" swimtime="00:08:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="430" swimtime="00:01:02.08" resultid="2708" heatid="4342" lane="7" entrytime="00:01:02.83" entrycourse="LCM" />
                <RESULT eventid="1258" points="474" swimtime="00:18:36.89" resultid="2709" heatid="4432" lane="0" entrytime="00:19:13.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.34" />
                    <SPLIT distance="200" swimtime="00:02:21.56" />
                    <SPLIT distance="300" swimtime="00:03:35.68" />
                    <SPLIT distance="400" swimtime="00:04:50.16" />
                    <SPLIT distance="500" swimtime="00:06:05.27" />
                    <SPLIT distance="600" swimtime="00:07:20.06" />
                    <SPLIT distance="700" swimtime="00:08:34.50" />
                    <SPLIT distance="800" swimtime="00:09:49.67" />
                    <SPLIT distance="900" swimtime="00:11:04.32" />
                    <SPLIT distance="1000" swimtime="00:12:19.22" />
                    <SPLIT distance="1100" swimtime="00:13:35.07" />
                    <SPLIT distance="1200" swimtime="00:14:50.46" />
                    <SPLIT distance="1300" swimtime="00:16:05.96" />
                    <SPLIT distance="1400" swimtime="00:17:22.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="442" swimtime="00:02:13.85" resultid="2710" heatid="4466" lane="8" entrytime="00:02:14.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="464" swimtime="00:04:44.06" resultid="2711" heatid="4515" lane="8" entrytime="00:04:48.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.95" />
                    <SPLIT distance="200" swimtime="00:02:17.98" />
                    <SPLIT distance="300" swimtime="00:03:31.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ferreira Motta" birthdate="2008-10-24" gender="M" nation="BRA" license="378068" swrid="5600160" athleteid="2902" externalid="378068">
              <RESULTS>
                <RESULT eventid="1088" points="418" swimtime="00:02:47.77" resultid="2903" heatid="4287" lane="5" entrytime="00:02:46.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="402" swimtime="00:00:35.14" resultid="2904" heatid="4367" lane="2" entrytime="00:00:35.20" entrycourse="LCM" />
                <RESULT eventid="1220" points="413" swimtime="00:01:16.35" resultid="2905" heatid="4393" lane="1" entrytime="00:01:15.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="CAUê" lastname="Glück" lastname.en="Gluck" birthdate="2006-07-16" gender="M" nation="BRA" license="296595" athleteid="2503" externalid="296595">
              <RESULTS>
                <RESULT eventid="1156" points="744" swimtime="00:00:51.70" resultid="2504" heatid="4348" lane="5" entrytime="00:00:51.46" entrycourse="LCM" />
                <RESULT eventid="1290" points="786" swimtime="00:01:50.51" resultid="2505" heatid="4469" lane="4" entrytime="00:01:51.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:53.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="783" swimtime="00:03:58.69" resultid="2506" heatid="4516" lane="4" entrytime="00:03:58.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.32" />
                    <SPLIT distance="200" swimtime="00:01:57.40" />
                    <SPLIT distance="300" swimtime="00:02:57.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Gustavo Souza" birthdate="2011-08-24" gender="M" nation="BRA" license="366901" swrid="5588733" athleteid="2793" externalid="366901">
              <RESULTS>
                <RESULT eventid="1172" points="291" swimtime="00:02:46.38" resultid="2794" heatid="4352" lane="4" entrytime="00:02:49.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="355" swimtime="00:20:29.27" resultid="2795" heatid="4430" lane="3" entrytime="00:21:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.73" />
                    <SPLIT distance="200" swimtime="00:02:44.32" />
                    <SPLIT distance="300" swimtime="00:04:08.96" />
                    <SPLIT distance="400" swimtime="00:05:32.49" />
                    <SPLIT distance="500" swimtime="00:06:57.82" />
                    <SPLIT distance="600" swimtime="00:08:21.33" />
                    <SPLIT distance="700" swimtime="00:09:44.19" />
                    <SPLIT distance="800" swimtime="00:11:06.61" />
                    <SPLIT distance="1100" swimtime="00:15:14.20" />
                    <SPLIT distance="1200" swimtime="00:16:34.07" />
                    <SPLIT distance="1300" swimtime="00:17:55.03" />
                    <SPLIT distance="1400" swimtime="00:19:15.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1274" points="294" swimtime="00:02:51.30" resultid="2796" heatid="4443" lane="6" entrytime="00:03:03.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="349" swimtime="00:05:12.50" resultid="2797" heatid="4513" lane="5" entrytime="00:05:15.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.26" />
                    <SPLIT distance="200" swimtime="00:02:39.01" />
                    <SPLIT distance="300" swimtime="00:03:58.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="292" swimtime="00:01:14.50" resultid="2798" heatid="4501" lane="8" entrytime="00:01:15.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Muxfeldt" birthdate="2011-05-13" gender="F" nation="BRA" license="366903" swrid="5602563" athleteid="2799" externalid="366903">
              <RESULTS>
                <RESULT eventid="1080" points="370" swimtime="00:03:11.59" resultid="2800" heatid="4280" lane="5" entrytime="00:03:08.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="444" swimtime="00:01:07.77" resultid="2801" heatid="4326" lane="8" entrytime="00:01:10.07" entrycourse="LCM" />
                <RESULT eventid="1228" points="411" swimtime="00:00:31.73" resultid="2802" heatid="4401" lane="1" entrytime="00:00:32.56" entrycourse="LCM" />
                <RESULT eventid="1212" points="352" swimtime="00:01:30.81" resultid="2803" heatid="4382" lane="2" entrytime="00:01:28.54" entrycourse="LCM" />
                <RESULT eventid="1282" points="418" swimtime="00:02:30.91" resultid="2804" heatid="4454" lane="4" entrytime="00:02:31.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Francisco Saldo" birthdate="2007-01-23" gender="M" nation="BRA" license="313537" swrid="5600169" athleteid="2507" externalid="313537">
              <RESULTS>
                <RESULT eventid="1104" points="519" swimtime="00:00:27.71" resultid="2508" heatid="4295" lane="5" />
                <RESULT eventid="1172" points="702" swimtime="00:02:04.15" resultid="2509" heatid="4354" lane="4" entrytime="00:02:02.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="499" swimtime="00:01:11.67" resultid="2510" heatid="4386" lane="5" />
                <RESULT eventid="1274" points="613" swimtime="00:02:14.15" resultid="2511" heatid="4448" lane="3" entrytime="00:02:13.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="661" swimtime="00:00:56.74" resultid="2512" heatid="4505" lane="4" entrytime="00:00:56.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Cabrera Cirino" birthdate="2011-01-28" gender="M" nation="BRA" license="369531" swrid="5588569" athleteid="2857" externalid="369531">
              <RESULTS>
                <RESULT eventid="1072" points="402" swimtime="00:02:31.54" resultid="2858" heatid="4275" lane="5" entrytime="00:02:31.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="460" swimtime="00:01:00.69" resultid="2859" heatid="4342" lane="5" entrytime="00:01:02.09" entrycourse="LCM" />
                <RESULT eventid="1236" points="431" swimtime="00:00:27.68" resultid="2860" heatid="4416" lane="7" entrytime="00:00:28.44" entrycourse="LCM" />
                <RESULT eventid="1290" points="426" swimtime="00:02:15.49" resultid="2861" heatid="4465" lane="6" entrytime="00:02:17.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="427" swimtime="00:04:52.14" resultid="2862" heatid="4514" lane="4" entrytime="00:04:56.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.48" />
                    <SPLIT distance="200" swimtime="00:02:25.10" />
                    <SPLIT distance="300" swimtime="00:03:40.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Fantin Dias De Andrade" birthdate="2010-11-06" gender="F" nation="BRA" license="339262" swrid="5588684" athleteid="2863" externalid="339262">
              <RESULTS>
                <RESULT eventid="1080" points="300" swimtime="00:03:25.46" resultid="2864" heatid="4279" lane="4" entrytime="00:03:20.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="334" swimtime="00:01:14.49" resultid="2865" heatid="4323" lane="2" entrytime="00:01:13.89" entrycourse="LCM" />
                <RESULT eventid="1228" points="361" swimtime="00:00:33.13" resultid="2866" heatid="4400" lane="4" entrytime="00:00:32.70" entrycourse="LCM" />
                <RESULT eventid="1212" points="289" swimtime="00:01:36.90" resultid="2867" heatid="4381" lane="2" entrytime="00:01:33.13" entrycourse="LCM" />
                <RESULT eventid="1266" points="314" swimtime="00:03:05.42" resultid="2868" heatid="4436" lane="5" entrytime="00:03:03.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabelly" lastname="Sinnott" birthdate="2009-03-14" gender="F" nation="BRA" license="367255" swrid="5600258" athleteid="2520" externalid="367255">
              <RESULTS>
                <RESULT eventid="1116" points="547" swimtime="00:18:44.92" resultid="2521" heatid="4309" lane="3" entrytime="00:18:45.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.10" />
                    <SPLIT distance="200" swimtime="00:02:25.04" />
                    <SPLIT distance="300" swimtime="00:03:40.42" />
                    <SPLIT distance="400" swimtime="00:04:56.11" />
                    <SPLIT distance="500" swimtime="00:06:11.85" />
                    <SPLIT distance="600" swimtime="00:07:26.95" />
                    <SPLIT distance="700" swimtime="00:08:42.12" />
                    <SPLIT distance="800" swimtime="00:09:57.38" />
                    <SPLIT distance="900" swimtime="00:11:13.14" />
                    <SPLIT distance="1000" swimtime="00:12:28.59" />
                    <SPLIT distance="1100" swimtime="00:13:44.25" />
                    <SPLIT distance="1200" swimtime="00:15:00.05" />
                    <SPLIT distance="1300" swimtime="00:16:16.04" />
                    <SPLIT distance="1400" swimtime="00:17:31.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="581" swimtime="00:01:01.95" resultid="2522" heatid="4330" lane="7" entrytime="00:01:01.98" entrycourse="LCM" />
                <RESULT eventid="1250" points="552" swimtime="00:09:50.70" resultid="2523" heatid="4428" lane="6" entrytime="00:09:47.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.93" />
                    <SPLIT distance="200" swimtime="00:02:24.17" />
                    <SPLIT distance="300" swimtime="00:03:39.99" />
                    <SPLIT distance="400" swimtime="00:04:55.31" />
                    <SPLIT distance="500" swimtime="00:06:10.16" />
                    <SPLIT distance="600" swimtime="00:07:24.81" />
                    <SPLIT distance="700" swimtime="00:08:38.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="618" swimtime="00:02:12.48" resultid="2524" heatid="4457" lane="2" entrytime="00:02:12.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="560" swimtime="00:04:45.49" resultid="2525" heatid="4510" lane="6" entrytime="00:04:38.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.15" />
                    <SPLIT distance="200" swimtime="00:02:20.02" />
                    <SPLIT distance="300" swimtime="00:03:32.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Magalhaes Dos Reis" birthdate="2010-05-05" gender="M" nation="BRA" license="356361" swrid="5600207" athleteid="2718" externalid="356361">
              <RESULTS>
                <RESULT eventid="1088" points="355" swimtime="00:02:57.17" resultid="2719" heatid="4286" lane="2" entrytime="00:02:56.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="468" swimtime="00:01:00.35" resultid="2720" heatid="4343" lane="4" entrytime="00:01:00.56" entrycourse="LCM" />
                <RESULT eventid="1220" points="344" swimtime="00:01:21.13" resultid="2721" heatid="4391" lane="6" entrytime="00:01:21.07" entrycourse="LCM" />
                <RESULT eventid="1274" points="339" swimtime="00:02:43.44" resultid="2722" heatid="4445" lane="1" entrytime="00:02:45.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Severo" lastname="Berger Leal" birthdate="2008-08-05" gender="M" nation="BRA" license="330073" swrid="5449277" athleteid="2586" externalid="330073">
              <RESULTS>
                <RESULT eventid="1088" status="DNS" swimtime="00:00:00.00" resultid="2587" heatid="4287" lane="7" entrytime="00:02:51.07" entrycourse="LCM" />
                <RESULT eventid="1188" points="377" swimtime="00:00:35.89" resultid="2588" heatid="4367" lane="8" entrytime="00:00:35.46" entrycourse="LCM" />
                <RESULT eventid="1220" points="348" swimtime="00:01:20.80" resultid="2589" heatid="4392" lane="6" entrytime="00:01:17.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Carneiro Silva" birthdate="2011-02-21" gender="F" nation="BRA" license="390924" swrid="5602522" athleteid="2945" externalid="390924">
              <RESULTS>
                <RESULT eventid="1064" points="337" swimtime="00:02:56.91" resultid="2946" heatid="4268" lane="3" entrytime="00:03:04.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="379" swimtime="00:01:11.45" resultid="2947" heatid="4323" lane="3" entrytime="00:01:13.76" entrycourse="LCM" />
                <RESULT eventid="1298" points="410" swimtime="00:00:36.15" resultid="2948" heatid="4473" lane="5" entrytime="00:00:37.83" entrycourse="LCM" />
                <RESULT eventid="1366" points="292" swimtime="00:01:26.40" resultid="2949" heatid="4521" lane="4" entrytime="00:01:21.20" entrycourse="LCM" />
                <RESULT eventid="1350" points="309" swimtime="00:05:47.86" resultid="2950" heatid="4507" lane="2" entrytime="00:05:46.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.51" />
                    <SPLIT distance="200" swimtime="00:02:47.68" />
                    <SPLIT distance="300" swimtime="00:04:17.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Fontoura" birthdate="2010-08-26" gender="M" nation="BRA" license="338922" swrid="5600167" athleteid="2729" externalid="338922">
              <RESULTS>
                <RESULT eventid="1156" points="378" swimtime="00:01:04.78" resultid="2730" heatid="4341" lane="1" entrytime="00:01:05.38" entrycourse="LCM" />
                <RESULT eventid="1140" status="DSQ" swimtime="00:05:56.66" resultid="2731" heatid="4317" lane="1" entrytime="00:05:59.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.08" />
                    <SPLIT distance="200" swimtime="00:02:52.30" />
                    <SPLIT distance="300" swimtime="00:04:36.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="353" swimtime="00:00:29.57" resultid="2732" heatid="4413" lane="1" entrytime="00:00:31.08" entrycourse="LCM" />
                <RESULT eventid="1274" points="318" swimtime="00:02:46.92" resultid="2733" heatid="4443" lane="3" entrytime="00:03:00.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="274" swimtime="00:01:16.10" resultid="2734" heatid="4500" lane="6" entrytime="00:01:17.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manoela" lastname="Andrade" birthdate="2010-03-10" gender="F" nation="BRA" license="339042" swrid="5363102" athleteid="2735" externalid="339042">
              <RESULTS>
                <RESULT eventid="1250" points="374" swimtime="00:11:12.34" resultid="2736" heatid="4427" lane="2" entrytime="00:10:49.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.62" />
                    <SPLIT distance="200" swimtime="00:02:42.26" />
                    <SPLIT distance="300" swimtime="00:04:06.22" />
                    <SPLIT distance="400" swimtime="00:05:32.18" />
                    <SPLIT distance="500" swimtime="00:06:58.51" />
                    <SPLIT distance="600" swimtime="00:08:24.57" />
                    <SPLIT distance="700" swimtime="00:09:48.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="359" swimtime="00:02:38.71" resultid="2737" heatid="4453" lane="5" entrytime="00:02:34.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="269" swimtime="00:01:25.85" resultid="2738" heatid="4496" lane="1" entrytime="00:01:19.51" entrycourse="LCM" />
                <RESULT eventid="1350" points="331" swimtime="00:05:39.94" resultid="2739" heatid="4508" lane="4" entrytime="00:05:25.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.37" />
                    <SPLIT distance="200" swimtime="00:02:46.55" />
                    <SPLIT distance="300" swimtime="00:04:14.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Rocha" birthdate="2011-08-25" gender="F" nation="BRA" license="366904" swrid="5602578" athleteid="2805" externalid="366904">
              <RESULTS>
                <RESULT eventid="1064" points="391" swimtime="00:02:48.33" resultid="2806" heatid="4269" lane="4" entrytime="00:02:52.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="464" swimtime="00:01:06.79" resultid="2807" heatid="4327" lane="5" entrytime="00:01:07.33" entrycourse="LCM" />
                <RESULT eventid="1228" points="473" swimtime="00:00:30.30" resultid="2808" heatid="4403" lane="1" entrytime="00:00:30.77" entrycourse="LCM" />
                <RESULT eventid="1282" points="461" swimtime="00:02:25.99" resultid="2809" heatid="4455" lane="5" entrytime="00:02:26.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="395" swimtime="00:01:18.07" resultid="2810" heatid="4522" lane="2" entrytime="00:01:19.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorena" lastname="Mascarenhas" birthdate="2011-08-31" gender="F" nation="BRA" license="370581" swrid="5602558" athleteid="2869" externalid="370581">
              <RESULTS>
                <RESULT eventid="1064" points="373" swimtime="00:02:50.97" resultid="2870" heatid="4270" lane="7" entrytime="00:02:49.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="411" swimtime="00:01:09.54" resultid="2871" heatid="4325" lane="4" entrytime="00:01:10.32" entrycourse="LCM" />
                <RESULT eventid="1212" points="307" swimtime="00:01:35.01" resultid="2872" heatid="4378" lane="2" />
                <RESULT eventid="1282" points="394" swimtime="00:02:33.91" resultid="2873" heatid="4453" lane="4" entrytime="00:02:34.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="384" swimtime="00:01:18.81" resultid="2874" heatid="4522" lane="8" entrytime="00:01:20.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Moreira Segadaes" birthdate="2008-05-15" gender="M" nation="BRA" license="331574" swrid="5600220" athleteid="2494" externalid="331574">
              <RESULTS>
                <RESULT eventid="1088" points="536" swimtime="00:02:34.44" resultid="2495" heatid="4288" lane="4" entrytime="00:02:33.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="578" swimtime="00:00:31.14" resultid="2496" heatid="4368" lane="5" entrytime="00:00:31.74" entrycourse="LCM" />
                <RESULT eventid="1220" points="529" swimtime="00:01:10.29" resultid="2497" heatid="4394" lane="5" entrytime="00:01:09.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Sabedotti" birthdate="2002-07-07" gender="M" nation="BRA" license="134704" swrid="5600252" athleteid="2652" externalid="134704">
              <RESULTS>
                <RESULT eventid="1156" points="696" swimtime="00:00:52.86" resultid="2653" heatid="4348" lane="2" entrytime="00:00:52.82" entrycourse="LCM" />
                <RESULT eventid="1188" points="657" swimtime="00:00:29.85" resultid="2654" heatid="4369" lane="3" entrytime="00:00:28.96" entrycourse="LCM" />
                <RESULT eventid="1220" points="616" swimtime="00:01:06.84" resultid="2655" heatid="4395" lane="6" entrytime="00:01:04.14" entrycourse="LCM" />
                <RESULT eventid="1236" points="634" swimtime="00:00:24.34" resultid="2656" heatid="4422" lane="2" entrytime="00:00:23.74" entrycourse="LCM" />
                <RESULT eventid="1274" points="660" swimtime="00:02:10.90" resultid="2657" heatid="4448" lane="4" entrytime="00:02:06.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="LIV" lastname="Carvalho" birthdate="2011-09-13" gender="F" nation="BRA" license="366899" swrid="5602524" athleteid="2787" externalid="366899">
              <RESULTS>
                <RESULT eventid="1080" points="303" swimtime="00:03:24.65" resultid="2788" heatid="4279" lane="6" entrytime="00:03:23.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="325" swimtime="00:01:15.19" resultid="2789" heatid="4321" lane="5" entrytime="00:01:23.25" entrycourse="LCM" />
                <RESULT eventid="1180" points="311" swimtime="00:00:43.03" resultid="2790" heatid="4356" lane="3" entrytime="00:00:49.61" entrycourse="LCM" />
                <RESULT eventid="1212" points="275" swimtime="00:01:38.54" resultid="2791" heatid="4380" lane="5" entrytime="00:01:37.48" entrycourse="LCM" />
                <RESULT eventid="1282" points="322" swimtime="00:02:44.61" resultid="2792" heatid="4451" lane="4" entrytime="00:02:52.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Cristina Ferreira" birthdate="2011-08-24" gender="F" nation="BRA" license="358334" swrid="5588611" athleteid="2881" externalid="358334">
              <RESULTS>
                <RESULT eventid="1080" points="549" swimtime="00:02:47.89" resultid="2882" heatid="4282" lane="6" entrytime="00:02:54.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="639" swimtime="00:02:21.40" resultid="2883" heatid="4350" lane="4" entrytime="00:02:27.98" entrycourse="LCM" />
                <RESULT eventid="1266" points="593" swimtime="00:02:30.04" resultid="2884" heatid="4435" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="625" swimtime="00:01:04.86" resultid="2885" heatid="4497" lane="3" entrytime="00:01:04.99" entrycourse="LCM" />
                <RESULT eventid="1350" points="588" swimtime="00:04:40.85" resultid="2886" heatid="4510" lane="2" entrytime="00:04:45.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.78" />
                    <SPLIT distance="200" swimtime="00:02:20.00" />
                    <SPLIT distance="300" swimtime="00:03:31.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="David Cella" birthdate="2008-02-17" gender="M" nation="BRA" license="341107" swrid="5634581" athleteid="2957" externalid="341107">
              <RESULTS>
                <RESULT eventid="1156" points="622" swimtime="00:00:54.88" resultid="2958" heatid="4347" lane="2" entrytime="00:00:55.13" entrycourse="LCM" />
                <RESULT eventid="1188" points="604" swimtime="00:00:30.69" resultid="2959" heatid="4369" lane="8" entrytime="00:00:31.31" entrycourse="LCM" />
                <RESULT eventid="1220" points="497" swimtime="00:01:11.80" resultid="2960" heatid="4394" lane="7" entrytime="00:01:11.28" entrycourse="LCM" />
                <RESULT eventid="1236" points="601" swimtime="00:00:24.77" resultid="2961" heatid="4421" lane="6" entrytime="00:00:24.79" entrycourse="LCM" />
                <RESULT eventid="1274" points="495" swimtime="00:02:24.07" resultid="2962" heatid="4447" lane="2" entrytime="00:02:27.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Araujo Barros" birthdate="2008-12-26" gender="M" nation="BRA" license="331713" swrid="5367497" athleteid="2851" externalid="331713">
              <RESULTS>
                <RESULT eventid="1124" points="558" swimtime="00:09:09.15" resultid="2852" heatid="4313" lane="3" entrytime="00:09:09.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.63" />
                    <SPLIT distance="200" swimtime="00:02:09.74" />
                    <SPLIT distance="300" swimtime="00:03:17.28" />
                    <SPLIT distance="400" swimtime="00:04:26.23" />
                    <SPLIT distance="500" swimtime="00:05:36.84" />
                    <SPLIT distance="600" swimtime="00:06:48.72" />
                    <SPLIT distance="700" swimtime="00:08:00.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="607" swimtime="00:00:55.32" resultid="2853" heatid="4347" lane="7" entrytime="00:00:55.89" entrycourse="LCM" />
                <RESULT eventid="1258" points="558" swimtime="00:17:37.66" resultid="2854" heatid="4432" lane="4" entrytime="00:17:57.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.51" />
                    <SPLIT distance="200" swimtime="00:02:15.26" />
                    <SPLIT distance="300" swimtime="00:03:25.56" />
                    <SPLIT distance="400" swimtime="00:04:35.51" />
                    <SPLIT distance="500" swimtime="00:05:46.31" />
                    <SPLIT distance="600" swimtime="00:06:57.01" />
                    <SPLIT distance="700" swimtime="00:08:07.40" />
                    <SPLIT distance="800" swimtime="00:09:19.25" />
                    <SPLIT distance="900" swimtime="00:10:30.64" />
                    <SPLIT distance="1000" swimtime="00:11:41.98" />
                    <SPLIT distance="1100" swimtime="00:12:53.31" />
                    <SPLIT distance="1200" swimtime="00:14:05.52" />
                    <SPLIT distance="1300" swimtime="00:15:17.42" />
                    <SPLIT distance="1400" swimtime="00:16:29.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="591" swimtime="00:02:01.52" resultid="2855" heatid="4468" lane="5" entrytime="00:02:01.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="581" swimtime="00:04:23.62" resultid="2856" heatid="4516" lane="2" entrytime="00:04:21.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.09" />
                    <SPLIT distance="200" swimtime="00:02:05.78" />
                    <SPLIT distance="300" swimtime="00:03:14.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Martinez Diniz" birthdate="2008-11-22" gender="M" nation="BRA" license="339400" swrid="5717283" athleteid="2590" externalid="339400">
              <RESULTS>
                <RESULT eventid="1124" points="433" swimtime="00:09:57.16" resultid="2591" heatid="4311" lane="3" entrytime="00:10:27.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.21" />
                    <SPLIT distance="200" swimtime="00:02:25.08" />
                    <SPLIT distance="300" swimtime="00:03:41.91" />
                    <SPLIT distance="400" swimtime="00:04:57.85" />
                    <SPLIT distance="500" swimtime="00:06:13.71" />
                    <SPLIT distance="600" swimtime="00:07:28.78" />
                    <SPLIT distance="700" swimtime="00:08:44.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="527" swimtime="00:00:58.01" resultid="2592" heatid="4332" lane="6" />
                <RESULT eventid="1236" points="468" swimtime="00:00:26.92" resultid="2593" heatid="4407" lane="7" />
                <RESULT eventid="1290" points="465" swimtime="00:02:11.64" resultid="2594" heatid="4466" lane="1" entrytime="00:02:14.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="451" swimtime="00:04:46.93" resultid="2595" heatid="4512" lane="8" entrytime="00:05:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.62" />
                    <SPLIT distance="200" swimtime="00:02:20.47" />
                    <SPLIT distance="300" swimtime="00:03:34.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Laurindo Netto" birthdate="2005-07-15" gender="M" nation="BRA" license="289995" swrid="5600198" athleteid="2468" externalid="289995">
              <RESULTS>
                <RESULT eventid="1072" points="493" swimtime="00:02:21.65" resultid="2469" heatid="4277" lane="2" entrytime="00:02:18.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="534" swimtime="00:04:58.73" resultid="2470" heatid="4318" lane="5" entrytime="00:04:44.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.47" />
                    <SPLIT distance="200" swimtime="00:02:22.36" />
                    <SPLIT distance="300" swimtime="00:03:48.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" status="DNS" swimtime="00:00:00.00" resultid="2471" heatid="4394" lane="3" entrytime="00:01:09.74" entrycourse="LCM" />
                <RESULT eventid="1274" status="DNS" swimtime="00:00:00.00" resultid="2472" heatid="4448" lane="5" entrytime="00:02:11.28" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Galvao" birthdate="2011-03-11" gender="M" nation="BRA" license="381989" swrid="5602541" athleteid="2906" externalid="381989">
              <RESULTS>
                <RESULT eventid="1124" points="305" swimtime="00:11:11.11" resultid="2907" heatid="4310" lane="4" entrytime="00:11:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.08" />
                    <SPLIT distance="200" swimtime="00:02:41.79" />
                    <SPLIT distance="300" swimtime="00:04:07.15" />
                    <SPLIT distance="400" swimtime="00:05:33.07" />
                    <SPLIT distance="500" swimtime="00:06:59.70" />
                    <SPLIT distance="600" swimtime="00:08:26.62" />
                    <SPLIT distance="700" swimtime="00:09:51.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="294" swimtime="00:01:10.42" resultid="2908" heatid="4338" lane="7" entrytime="00:01:08.37" entrycourse="LCM" />
                <RESULT eventid="1236" points="291" swimtime="00:00:31.52" resultid="2909" heatid="4412" lane="2" entrytime="00:00:32.44" entrycourse="LCM" />
                <RESULT eventid="1290" points="293" swimtime="00:02:33.48" resultid="2910" heatid="4462" lane="7" entrytime="00:02:33.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Bussmann" birthdate="2007-01-16" gender="F" nation="BRA" license="313781" swrid="5579983" athleteid="2498" externalid="313781">
              <RESULTS>
                <RESULT eventid="1080" points="628" swimtime="00:02:40.58" resultid="2499" heatid="4282" lane="4" entrytime="00:02:39.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="553" swimtime="00:00:35.51" resultid="2500" heatid="4359" lane="3" entrytime="00:00:35.65" entrycourse="LCM" />
                <RESULT eventid="1212" points="581" swimtime="00:01:16.85" resultid="2501" heatid="4384" lane="5" entrytime="00:01:15.11" entrycourse="LCM" />
                <RESULT eventid="1266" status="DNS" swimtime="00:00:00.00" resultid="2502" heatid="4439" lane="4" entrytime="00:02:33.27" entrycourse="LCM" />
                <RESULT eventid="4970" points="630" swimtime="00:01:14.79" resultid="4973" heatid="4972" lane="4" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinícius" lastname="Oliveira Cruz" birthdate="2005-07-02" gender="M" nation="BRA" license="298495" swrid="5653299" athleteid="2982" externalid="298495">
              <RESULTS>
                <RESULT eventid="1156" points="740" swimtime="00:00:51.79" resultid="2983" heatid="4348" lane="3" entrytime="00:00:51.56" entrycourse="LCM" />
                <RESULT eventid="1236" points="660" swimtime="00:00:24.01" resultid="2984" heatid="4422" lane="6" entrytime="00:00:23.64" entrycourse="LCM" />
                <RESULT eventid="1290" points="747" swimtime="00:01:52.41" resultid="2985" heatid="4469" lane="5" entrytime="00:01:51.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="701" swimtime="00:04:07.70" resultid="2986" heatid="4516" lane="5" entrytime="00:04:10.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.87" />
                    <SPLIT distance="200" swimtime="00:02:02.66" />
                    <SPLIT distance="300" swimtime="00:03:04.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Germer Munhoz" birthdate="2010-04-23" gender="F" nation="BRA" license="356632" swrid="5588722" athleteid="2723" externalid="356632">
              <RESULTS>
                <RESULT eventid="1164" points="368" swimtime="00:02:49.93" resultid="2724" heatid="4350" lane="7" entrytime="00:02:52.30" entrycourse="LCM" />
                <RESULT eventid="1250" points="475" swimtime="00:10:20.92" resultid="2725" heatid="4428" lane="8" entrytime="00:10:14.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.02" />
                    <SPLIT distance="200" swimtime="00:02:29.34" />
                    <SPLIT distance="300" swimtime="00:03:48.11" />
                    <SPLIT distance="400" swimtime="00:05:07.54" />
                    <SPLIT distance="500" swimtime="00:06:26.77" />
                    <SPLIT distance="600" swimtime="00:07:46.26" />
                    <SPLIT distance="700" swimtime="00:09:05.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" points="449" swimtime="00:02:44.66" resultid="2726" heatid="4438" lane="5" entrytime="00:02:49.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="397" swimtime="00:01:15.44" resultid="2727" heatid="4496" lane="4" entrytime="00:01:16.66" entrycourse="LCM" />
                <RESULT eventid="1350" points="459" swimtime="00:05:04.92" resultid="2728" heatid="4509" lane="3" entrytime="00:05:06.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.82" />
                    <SPLIT distance="200" swimtime="00:02:31.46" />
                    <SPLIT distance="300" swimtime="00:03:50.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rene" lastname="Osternack Erbe" birthdate="2011-04-03" gender="M" nation="BRA" license="366907" swrid="5588842" athleteid="2817" externalid="366907">
              <RESULTS>
                <RESULT eventid="1156" points="306" swimtime="00:01:09.51" resultid="2818" heatid="4336" lane="2" entrytime="00:01:13.02" entrycourse="LCM" />
                <RESULT eventid="1236" points="281" swimtime="00:00:31.89" resultid="2819" heatid="4412" lane="8" entrytime="00:00:33.09" entrycourse="LCM" />
                <RESULT eventid="1274" points="261" swimtime="00:02:58.28" resultid="2820" heatid="4441" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="322" swimtime="00:05:20.89" resultid="2821" heatid="4513" lane="8" entrytime="00:05:27.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.57" />
                    <SPLIT distance="200" swimtime="00:02:41.04" />
                    <SPLIT distance="300" swimtime="00:04:02.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="247" swimtime="00:01:22.19" resultid="2822" heatid="4527" lane="4" entrytime="00:01:21.28" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Brandt De Macedo" birthdate="2006-04-22" gender="M" nation="BRA" license="296648" swrid="5622265" athleteid="2518" externalid="296648">
              <RESULTS>
                <RESULT eventid="1290" points="667" swimtime="00:01:56.70" resultid="2519" heatid="4469" lane="1" entrytime="00:02:00.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Artigas Pinheiro" birthdate="2011-08-25" gender="M" nation="BRA" license="377040" swrid="5588535" athleteid="2896" externalid="377040">
              <RESULTS>
                <RESULT eventid="1088" points="297" swimtime="00:03:07.98" resultid="2897" heatid="4285" lane="2" entrytime="00:03:10.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="213" swimtime="00:03:04.70" resultid="2898" heatid="4352" lane="1" entrytime="00:03:06.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="277" swimtime="00:01:27.22" resultid="2899" heatid="4389" lane="8" entrytime="00:01:32.95" entrycourse="LCM" />
                <RESULT eventid="1274" points="274" swimtime="00:02:55.48" resultid="2900" heatid="4443" lane="7" entrytime="00:03:04.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="303" swimtime="00:05:27.64" resultid="2901" heatid="4512" lane="7" entrytime="00:05:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.27" />
                    <SPLIT distance="200" swimtime="00:02:43.39" />
                    <SPLIT distance="300" swimtime="00:04:07.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Perroni Ribeiro" birthdate="2004-11-06" gender="F" nation="BRA" license="310555" athleteid="2974" externalid="310555">
              <RESULTS>
                <RESULT eventid="1116" points="519" swimtime="00:19:04.84" resultid="2975" heatid="4308" lane="6" entrytime="00:22:41.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                    <SPLIT distance="200" swimtime="00:02:28.92" />
                    <SPLIT distance="300" swimtime="00:03:45.41" />
                    <SPLIT distance="400" swimtime="00:05:02.14" />
                    <SPLIT distance="500" swimtime="00:06:19.47" />
                    <SPLIT distance="600" swimtime="00:07:35.36" />
                    <SPLIT distance="700" swimtime="00:08:51.91" />
                    <SPLIT distance="800" swimtime="00:10:08.75" />
                    <SPLIT distance="900" swimtime="00:11:25.71" />
                    <SPLIT distance="1000" swimtime="00:12:42.87" />
                    <SPLIT distance="1100" swimtime="00:13:59.04" />
                    <SPLIT distance="1200" swimtime="00:15:15.75" />
                    <SPLIT distance="1300" swimtime="00:16:32.38" />
                    <SPLIT distance="1400" swimtime="00:17:49.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="535" swimtime="00:09:57.13" resultid="2976" heatid="4426" lane="9" entrytime="00:11:57.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.35" />
                    <SPLIT distance="200" swimtime="00:02:29.18" />
                    <SPLIT distance="300" swimtime="00:03:44.74" />
                    <SPLIT distance="400" swimtime="00:05:00.68" />
                    <SPLIT distance="500" swimtime="00:06:15.79" />
                    <SPLIT distance="600" swimtime="00:07:29.84" />
                    <SPLIT distance="700" swimtime="00:08:44.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" status="DNS" swimtime="00:00:00.00" resultid="2977" heatid="4506" lane="5" entrytime="00:05:46.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="De Czarnecki" birthdate="2008-06-24" gender="M" nation="BRA" license="329641" swrid="5600146" athleteid="2473" externalid="329641">
              <RESULTS>
                <RESULT eventid="1072" points="459" swimtime="00:02:25.00" resultid="2474" heatid="4277" lane="3" entrytime="00:02:13.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" status="DNS" swimtime="00:00:00.00" resultid="2475" heatid="4316" lane="6" entrytime="00:06:23.00" entrycourse="LCM" />
                <RESULT eventid="1306" points="539" swimtime="00:00:28.92" resultid="2476" heatid="4476" lane="3" />
                <RESULT eventid="1374" points="562" swimtime="00:01:02.51" resultid="2477" heatid="4533" lane="6" entrytime="00:01:01.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Lacerda" birthdate="2011-05-09" gender="M" nation="BRA" license="366909" swrid="5602550" athleteid="2829" externalid="366909">
              <RESULTS>
                <RESULT eventid="1088" status="DSQ" swimtime="00:00:00.00" resultid="2830" heatid="4285" lane="6" entrytime="00:03:09.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="272" swimtime="00:01:27.69" resultid="2831" heatid="4390" lane="1" entrytime="00:01:28.88" entrycourse="LCM" />
                <RESULT eventid="1274" points="328" swimtime="00:02:45.21" resultid="2832" heatid="4444" lane="5" entrytime="00:02:51.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="364" swimtime="00:05:07.96" resultid="2833" heatid="4512" lane="5" entrytime="00:05:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.49" />
                    <SPLIT distance="200" swimtime="00:02:33.80" />
                    <SPLIT distance="300" swimtime="00:03:53.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicole" lastname="Rosario Osternack" birthdate="2008-04-11" gender="F" nation="BRA" license="331584" swrid="5600248" athleteid="2454" externalid="331584">
              <RESULTS>
                <RESULT eventid="1096" points="535" swimtime="00:00:30.08" resultid="2455" heatid="4294" lane="3" entrytime="00:00:30.71" entrycourse="LCM" />
                <RESULT eventid="1164" points="385" swimtime="00:02:47.30" resultid="2456" heatid="4349" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" points="542" swimtime="00:02:34.63" resultid="2457" heatid="4439" lane="5" entrytime="00:02:36.67" entrycourse="LCM" />
                <RESULT eventid="1334" points="557" swimtime="00:01:07.42" resultid="2458" heatid="4497" lane="6" entrytime="00:01:07.15" entrycourse="LCM" />
                <RESULT eventid="1366" points="535" swimtime="00:01:10.62" resultid="2459" heatid="4524" lane="7" entrytime="00:01:10.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucca" lastname="Cruz Tonin" birthdate="2004-03-19" gender="M" nation="BRA" license="270821" swrid="5622272" athleteid="2834" externalid="270821">
              <RESULTS>
                <RESULT eventid="1072" points="723" swimtime="00:02:04.69" resultid="2835" heatid="4277" lane="4" entrytime="00:02:02.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="753" swimtime="00:00:51.50" resultid="2836" heatid="4333" lane="1" />
                <RESULT eventid="1306" points="701" swimtime="00:00:26.50" resultid="2837" heatid="4482" lane="4" entrytime="00:00:26.89" entrycourse="LCM" />
                <RESULT eventid="1374" points="741" swimtime="00:00:57.00" resultid="2838" heatid="4533" lane="4" entrytime="00:00:56.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Coelho" birthdate="2011-11-11" gender="M" nation="BRA" license="366889" swrid="5602527" athleteid="2757" externalid="366889">
              <RESULTS>
                <RESULT eventid="1124" points="375" swimtime="00:10:26.42" resultid="2758" heatid="4312" lane="8" entrytime="00:10:15.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.76" />
                    <SPLIT distance="200" swimtime="00:02:32.72" />
                    <SPLIT distance="300" swimtime="00:03:51.88" />
                    <SPLIT distance="400" swimtime="00:05:11.80" />
                    <SPLIT distance="500" swimtime="00:06:30.86" />
                    <SPLIT distance="600" swimtime="00:07:50.47" />
                    <SPLIT distance="700" swimtime="00:09:09.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="275" swimtime="00:02:49.67" resultid="2759" heatid="4352" lane="6" entrytime="00:02:54.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="366" swimtime="00:02:22.47" resultid="2760" heatid="4464" lane="7" entrytime="00:02:23.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="378" swimtime="00:05:04.31" resultid="2761" heatid="4513" lane="3" entrytime="00:05:16.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.10" />
                    <SPLIT distance="200" swimtime="00:02:29.31" />
                    <SPLIT distance="300" swimtime="00:03:47.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="312" swimtime="00:01:12.90" resultid="2762" heatid="4500" lane="4" entrytime="00:01:16.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Godino" birthdate="2010-04-27" gender="F" nation="BRA" license="356355" swrid="5600176" athleteid="2712" externalid="356355">
              <RESULTS>
                <RESULT eventid="1064" points="312" swimtime="00:03:01.52" resultid="2713" heatid="4268" lane="4" entrytime="00:03:02.54" entrycourse="LCM" />
                <RESULT eventid="1148" points="417" swimtime="00:01:09.21" resultid="2714" heatid="4325" lane="7" entrytime="00:01:11.24" entrycourse="LCM" />
                <RESULT eventid="1250" points="429" swimtime="00:10:42.33" resultid="2715" heatid="4427" lane="5" entrytime="00:10:40.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.67" />
                    <SPLIT distance="200" swimtime="00:02:33.59" />
                    <SPLIT distance="300" swimtime="00:03:54.85" />
                    <SPLIT distance="400" swimtime="00:05:16.65" />
                    <SPLIT distance="500" swimtime="00:06:38.27" />
                    <SPLIT distance="600" swimtime="00:08:00.42" />
                    <SPLIT distance="700" swimtime="00:09:22.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="422" swimtime="00:02:30.35" resultid="2716" heatid="4455" lane="7" entrytime="00:02:30.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="414" swimtime="00:05:15.68" resultid="2717" heatid="4509" lane="1" entrytime="00:05:17.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.11" />
                    <SPLIT distance="200" swimtime="00:02:34.95" />
                    <SPLIT distance="300" swimtime="00:03:55.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Vitoria Kuzmann Cercal" birthdate="2009-04-10" gender="F" nation="BRA" license="339082" swrid="5600274" athleteid="2625" externalid="339082">
              <RESULTS>
                <RESULT eventid="1064" points="401" swimtime="00:02:46.96" resultid="2626" heatid="4270" lane="6" entrytime="00:02:46.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="495" swimtime="00:01:05.33" resultid="2627" heatid="4328" lane="3" entrytime="00:01:05.90" entrycourse="LCM" />
                <RESULT eventid="1250" points="396" swimtime="00:10:59.75" resultid="2628" heatid="4427" lane="3" entrytime="00:10:40.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.78" />
                    <SPLIT distance="200" swimtime="00:02:33.05" />
                    <SPLIT distance="300" swimtime="00:03:56.20" />
                    <SPLIT distance="400" swimtime="00:05:21.12" />
                    <SPLIT distance="500" swimtime="00:06:47.19" />
                    <SPLIT distance="600" swimtime="00:08:13.47" />
                    <SPLIT distance="700" swimtime="00:09:39.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" status="DSQ" swimtime="00:02:46.43" resultid="2629" heatid="4438" lane="8" entrytime="00:02:56.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="433" swimtime="00:05:11.10" resultid="2630" heatid="4509" lane="5" entrytime="00:05:01.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.59" />
                    <SPLIT distance="200" swimtime="00:02:30.84" />
                    <SPLIT distance="300" swimtime="00:03:51.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelo" lastname="Vanhazebrouck" birthdate="2010-01-09" gender="M" nation="BRA" license="339043" swrid="5600269" athleteid="2658" externalid="339043">
              <RESULTS>
                <RESULT eventid="1088" points="306" swimtime="00:03:06.03" resultid="2659" heatid="4286" lane="1" entrytime="00:03:02.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="469" swimtime="00:01:00.30" resultid="2660" heatid="4343" lane="6" entrytime="00:01:00.98" entrycourse="LCM" />
                <RESULT eventid="1220" points="315" swimtime="00:01:23.53" resultid="2661" heatid="4391" lane="8" entrytime="00:01:23.11" entrycourse="LCM" />
                <RESULT eventid="1236" points="436" swimtime="00:00:27.57" resultid="2662" heatid="4415" lane="4" entrytime="00:00:28.62" entrycourse="LCM" />
                <RESULT eventid="1290" points="423" swimtime="00:02:15.87" resultid="2663" heatid="4465" lane="3" entrytime="00:02:16.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Iglesias Vargas" birthdate="2009-01-11" gender="M" nation="BRA" license="324792" swrid="5600189" athleteid="2536" externalid="324792">
              <RESULTS>
                <RESULT eventid="1124" points="463" swimtime="00:09:44.08" resultid="2537" heatid="4313" lane="7" entrytime="00:09:26.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.03" />
                    <SPLIT distance="200" swimtime="00:02:16.98" />
                    <SPLIT distance="300" swimtime="00:03:30.03" />
                    <SPLIT distance="400" swimtime="00:04:43.72" />
                    <SPLIT distance="500" swimtime="00:05:58.37" />
                    <SPLIT distance="600" swimtime="00:07:13.43" />
                    <SPLIT distance="700" swimtime="00:08:29.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="433" swimtime="00:05:20.37" resultid="2538" heatid="4316" lane="5" entrytime="00:06:23.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.22" />
                    <SPLIT distance="200" swimtime="00:02:30.56" />
                    <SPLIT distance="300" swimtime="00:04:06.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="476" swimtime="00:00:26.77" resultid="2539" heatid="4416" lane="4" entrytime="00:00:27.62" entrycourse="LCM" />
                <RESULT eventid="1274" points="477" swimtime="00:02:25.82" resultid="2540" heatid="4447" lane="7" entrytime="00:02:28.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="515" swimtime="00:04:34.54" resultid="2541" heatid="4516" lane="8" entrytime="00:04:34.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.71" />
                    <SPLIT distance="200" swimtime="00:02:11.09" />
                    <SPLIT distance="300" swimtime="00:03:22.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Leao" birthdate="2011-09-18" gender="M" nation="BRA" license="366880" swrid="5602553" athleteid="2751" externalid="366880">
              <RESULTS>
                <RESULT eventid="1124" points="391" swimtime="00:10:18.08" resultid="2752" heatid="4311" lane="5" entrytime="00:10:24.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.53" />
                    <SPLIT distance="200" swimtime="00:02:34.08" />
                    <SPLIT distance="300" swimtime="00:03:52.58" />
                    <SPLIT distance="400" swimtime="00:05:10.65" />
                    <SPLIT distance="500" swimtime="00:06:28.61" />
                    <SPLIT distance="600" swimtime="00:07:46.40" />
                    <SPLIT distance="700" swimtime="00:09:03.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="371" swimtime="00:01:05.18" resultid="2753" heatid="4340" lane="6" entrytime="00:01:06.02" entrycourse="LCM" />
                <RESULT eventid="1258" points="408" swimtime="00:19:34.15" resultid="2754" heatid="4430" lane="2" entrytime="00:21:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.40" />
                    <SPLIT distance="200" swimtime="00:02:32.00" />
                    <SPLIT distance="300" swimtime="00:03:50.46" />
                    <SPLIT distance="400" swimtime="00:05:07.91" />
                    <SPLIT distance="500" swimtime="00:06:26.14" />
                    <SPLIT distance="600" swimtime="00:07:43.99" />
                    <SPLIT distance="700" swimtime="00:09:02.81" />
                    <SPLIT distance="800" swimtime="00:10:22.01" />
                    <SPLIT distance="900" swimtime="00:11:41.83" />
                    <SPLIT distance="1000" swimtime="00:13:01.09" />
                    <SPLIT distance="1100" swimtime="00:14:20.65" />
                    <SPLIT distance="1200" swimtime="00:15:40.47" />
                    <SPLIT distance="1300" swimtime="00:16:59.64" />
                    <SPLIT distance="1400" swimtime="00:18:18.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="373" swimtime="00:02:21.60" resultid="2755" heatid="4463" lane="5" entrytime="00:02:25.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="400" swimtime="00:04:58.60" resultid="2756" heatid="4513" lane="4" entrytime="00:05:10.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.37" />
                    <SPLIT distance="200" swimtime="00:02:27.78" />
                    <SPLIT distance="300" swimtime="00:03:44.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolau" lastname="Neto" birthdate="2011-03-22" gender="M" nation="BRA" license="366906" swrid="5602565" athleteid="2811" externalid="366906">
              <RESULTS>
                <RESULT eventid="1088" points="321" swimtime="00:03:03.23" resultid="2812" heatid="4285" lane="5" entrytime="00:03:07.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="398" swimtime="00:01:03.67" resultid="2813" heatid="4341" lane="6" entrytime="00:01:04.66" entrycourse="LCM" />
                <RESULT eventid="1220" points="307" swimtime="00:01:24.23" resultid="2814" heatid="4390" lane="3" entrytime="00:01:24.42" entrycourse="LCM" />
                <RESULT eventid="1236" points="374" swimtime="00:00:29.00" resultid="2815" heatid="4413" lane="6" entrytime="00:00:30.80" entrycourse="LCM" />
                <RESULT eventid="1274" points="295" swimtime="00:02:51.14" resultid="2816" heatid="4444" lane="8" entrytime="00:02:58.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Yolanda Ferreira" birthdate="2008-03-17" gender="F" nation="BRA" license="358335" swrid="5600276" athleteid="2875" externalid="358335">
              <RESULTS>
                <RESULT eventid="1080" points="485" swimtime="00:02:54.96" resultid="2876" heatid="4282" lane="2" entrytime="00:02:55.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="517" swimtime="00:01:04.42" resultid="2877" heatid="4329" lane="1" entrytime="00:01:04.89" entrycourse="LCM" />
                <RESULT eventid="1180" points="472" swimtime="00:00:37.44" resultid="2878" heatid="4359" lane="2" entrytime="00:00:37.63" entrycourse="LCM" />
                <RESULT eventid="1228" points="492" swimtime="00:00:29.90" resultid="2879" heatid="4405" lane="8" entrytime="00:00:29.39" entrycourse="LCM" />
                <RESULT eventid="1212" points="486" swimtime="00:01:21.52" resultid="2880" heatid="4384" lane="2" entrytime="00:01:21.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="De Albuquerque" birthdate="2010-06-08" gender="F" nation="BRA" license="356249" swrid="5600145" athleteid="2670" externalid="356249">
              <RESULTS>
                <RESULT eventid="1064" points="398" swimtime="00:02:47.38" resultid="2671" heatid="4270" lane="5" entrytime="00:02:45.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="395" swimtime="00:01:10.44" resultid="2672" heatid="4325" lane="5" entrytime="00:01:10.55" entrycourse="LCM" />
                <RESULT eventid="1228" points="408" swimtime="00:00:31.83" resultid="2673" heatid="4401" lane="3" entrytime="00:00:31.99" entrycourse="LCM" />
                <RESULT eventid="1298" points="434" swimtime="00:00:35.45" resultid="2674" heatid="4474" lane="6" entrytime="00:00:36.96" entrycourse="LCM" />
                <RESULT eventid="1366" points="394" swimtime="00:01:18.15" resultid="2675" heatid="4523" lane="5" entrytime="00:01:16.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Pereira Galle" birthdate="2011-08-02" gender="F" nation="BRA" license="369465" swrid="5627330" athleteid="2951" externalid="369465">
              <RESULTS>
                <RESULT eventid="1080" points="358" swimtime="00:03:13.59" resultid="2952" heatid="4279" lane="3" entrytime="00:03:21.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="392" swimtime="00:01:27.57" resultid="2953" heatid="4382" lane="3" entrytime="00:01:28.00" entrycourse="LCM" />
                <RESULT eventid="1282" points="380" swimtime="00:02:35.68" resultid="2954" heatid="4454" lane="7" entrytime="00:02:33.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" points="351" swimtime="00:02:58.79" resultid="2955" heatid="4437" lane="1" entrytime="00:03:01.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="271" swimtime="00:01:25.69" resultid="2956" heatid="4495" lane="6" entrytime="00:01:30.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Henrique Pasqual" birthdate="2005-05-07" gender="M" nation="BRA" license="329284" swrid="5600185" athleteid="3011" externalid="329284">
              <RESULTS>
                <RESULT eventid="1104" points="678" swimtime="00:00:25.34" resultid="3012" heatid="4304" lane="5" entrytime="00:00:25.31" entrycourse="LCM" />
                <RESULT eventid="1156" points="652" swimtime="00:00:54.03" resultid="3013" heatid="4348" lane="7" entrytime="00:00:53.34" entrycourse="LCM" />
                <RESULT eventid="1236" points="658" swimtime="00:00:24.03" resultid="3014" heatid="4422" lane="7" entrytime="00:00:23.91" entrycourse="LCM" />
                <RESULT eventid="1290" points="608" swimtime="00:02:00.37" resultid="3015" heatid="4468" lane="4" entrytime="00:02:01.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="567" swimtime="00:00:59.74" resultid="3016" heatid="4505" lane="6" entrytime="00:00:58.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helen" lastname="Barato Bernardi" birthdate="2006-07-27" gender="F" nation="BRA" license="317031" swrid="5717244" athleteid="2978" externalid="317031">
              <RESULTS>
                <RESULT eventid="1080" points="619" swimtime="00:02:41.36" resultid="2979" heatid="4282" lane="5" entrytime="00:02:45.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="668" swimtime="00:00:33.35" resultid="2980" heatid="4359" lane="4" entrytime="00:00:33.44" entrycourse="LCM" />
                <RESULT eventid="1212" points="651" swimtime="00:01:13.97" resultid="2981" heatid="4384" lane="4" entrytime="00:01:14.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joshua" lastname="Gomide Capraro" birthdate="2009-01-18" gender="M" nation="BRA" license="339030" swrid="5600177" athleteid="2484" externalid="339030">
              <RESULTS>
                <RESULT eventid="1156" points="594" swimtime="00:00:55.71" resultid="2485" heatid="4347" lane="6" entrytime="00:00:55.09" entrycourse="LCM" />
                <RESULT eventid="1236" points="577" swimtime="00:00:25.11" resultid="2486" heatid="4421" lane="2" entrytime="00:00:24.96" entrycourse="LCM" />
                <RESULT eventid="1290" points="555" swimtime="00:02:04.10" resultid="2487" heatid="4468" lane="6" entrytime="00:02:03.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="431" swimtime="00:04:51.26" resultid="2488" heatid="4515" lane="4" entrytime="00:04:35.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.30" />
                    <SPLIT distance="200" swimtime="00:02:17.37" />
                    <SPLIT distance="300" swimtime="00:03:34.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Martynychen" birthdate="2011-12-19" gender="M" nation="BRA" license="366893" swrid="5602557" athleteid="2769" externalid="366893">
              <RESULTS>
                <RESULT eventid="1072" points="307" swimtime="00:02:45.77" resultid="2770" heatid="4274" lane="8" entrytime="00:02:49.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="382" swimtime="00:10:22.98" resultid="2771" heatid="4311" lane="2" entrytime="00:10:31.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.19" />
                    <SPLIT distance="200" swimtime="00:02:33.86" />
                    <SPLIT distance="300" swimtime="00:03:52.51" />
                    <SPLIT distance="400" swimtime="00:05:10.73" />
                    <SPLIT distance="500" swimtime="00:06:29.65" />
                    <SPLIT distance="600" swimtime="00:07:48.86" />
                    <SPLIT distance="700" swimtime="00:09:08.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="417" swimtime="00:19:25.33" resultid="2772" heatid="4430" lane="1" entrytime="00:21:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.49" />
                    <SPLIT distance="200" swimtime="00:02:32.73" />
                    <SPLIT distance="300" swimtime="00:03:51.41" />
                    <SPLIT distance="400" swimtime="00:05:08.91" />
                    <SPLIT distance="500" swimtime="00:06:26.35" />
                    <SPLIT distance="600" swimtime="00:07:43.17" />
                    <SPLIT distance="700" swimtime="00:08:59.63" />
                    <SPLIT distance="800" swimtime="00:10:17.77" />
                    <SPLIT distance="900" swimtime="00:11:35.97" />
                    <SPLIT distance="1000" swimtime="00:12:54.47" />
                    <SPLIT distance="1100" swimtime="00:14:12.78" />
                    <SPLIT distance="1200" swimtime="00:15:32.43" />
                    <SPLIT distance="1300" swimtime="00:16:50.46" />
                    <SPLIT distance="1400" swimtime="00:18:06.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="301" swimtime="00:02:32.06" resultid="2773" heatid="4463" lane="1" entrytime="00:02:27.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="369" swimtime="00:05:06.74" resultid="2774" heatid="4513" lane="6" entrytime="00:05:16.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.81" />
                    <SPLIT distance="200" swimtime="00:02:32.48" />
                    <SPLIT distance="300" swimtime="00:03:50.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Trevisan" birthdate="2000-11-28" gender="M" nation="BRA" license="346847" swrid="5600266" athleteid="2922" externalid="346847">
              <RESULTS>
                <RESULT eventid="1104" points="575" swimtime="00:00:26.77" resultid="2923" heatid="4304" lane="7" entrytime="00:00:26.98" entrycourse="LCM" />
                <RESULT eventid="1156" points="631" swimtime="00:00:54.62" resultid="2924" heatid="4347" lane="5" entrytime="00:00:54.74" entrycourse="LCM" />
                <RESULT eventid="1236" points="611" swimtime="00:00:24.63" resultid="2925" heatid="4422" lane="8" entrytime="00:00:24.46" entrycourse="LCM" />
                <RESULT eventid="1290" points="563" swimtime="00:02:03.48" resultid="2926" heatid="4468" lane="1" entrytime="00:02:05.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="521" swimtime="00:01:04.10" resultid="2927" heatid="4532" lane="5" entrytime="00:01:03.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Alves Franca Silva" birthdate="1987-05-14" gender="M" nation="BRA" license="059512" athleteid="2998" externalid="059512">
              <RESULTS>
                <RESULT eventid="1088" points="604" swimtime="00:02:28.40" resultid="2999" heatid="4289" lane="3" entrytime="00:02:17.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="676" swimtime="00:00:29.56" resultid="3000" heatid="4369" lane="4" entrytime="00:00:27.92" entrycourse="LCM" />
                <RESULT eventid="1220" status="DNS" swimtime="00:00:00.00" resultid="3001" heatid="4395" lane="5" entrytime="00:01:01.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Kirchgassner" birthdate="2007-02-10" gender="M" nation="BRA" license="313535" swrid="5600230" athleteid="2553" externalid="313535">
              <RESULTS>
                <RESULT eventid="1088" points="626" swimtime="00:02:26.63" resultid="2554" heatid="4289" lane="6" entrytime="00:02:21.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="578" swimtime="00:00:31.14" resultid="2555" heatid="4368" lane="4" entrytime="00:00:31.50" entrycourse="LCM" />
                <RESULT eventid="1220" points="623" swimtime="00:01:06.58" resultid="2556" heatid="4395" lane="7" entrytime="00:01:05.67" entrycourse="LCM" />
                <RESULT eventid="1274" points="554" swimtime="00:02:18.74" resultid="2557" heatid="4447" lane="4" entrytime="00:02:18.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="545" swimtime="00:01:00.51" resultid="2558" heatid="4504" lane="4" entrytime="00:01:01.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Cury" birthdate="2005-09-28" gender="M" nation="BRA" license="329251" swrid="5600270" athleteid="2746" externalid="329251">
              <RESULTS>
                <RESULT eventid="1104" points="616" swimtime="00:00:26.16" resultid="2747" heatid="4303" lane="4" entrytime="00:00:27.32" entrycourse="LCM" />
                <RESULT eventid="1172" points="626" swimtime="00:02:08.95" resultid="2748" heatid="4354" lane="5" entrytime="00:02:09.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="634" swimtime="00:01:58.70" resultid="2749" heatid="4469" lane="7" entrytime="00:01:59.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:57.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="638" swimtime="00:00:57.42" resultid="2750" heatid="4505" lane="3" entrytime="00:00:57.21" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thais" lastname="Mariany Bortolazzi" birthdate="2006-05-02" gender="F" nation="BRA" license="357048" swrid="5600210" athleteid="2887" externalid="357048">
              <RESULTS>
                <RESULT eventid="1116" points="636" swimtime="00:17:49.94" resultid="2888" heatid="4309" lane="5" entrytime="00:17:56.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.70" />
                    <SPLIT distance="200" swimtime="00:02:20.17" />
                    <SPLIT distance="300" swimtime="00:03:31.17" />
                    <SPLIT distance="400" swimtime="00:04:42.58" />
                    <SPLIT distance="500" swimtime="00:05:54.01" />
                    <SPLIT distance="600" swimtime="00:07:05.53" />
                    <SPLIT distance="700" swimtime="00:08:17.06" />
                    <SPLIT distance="800" swimtime="00:09:28.83" />
                    <SPLIT distance="900" swimtime="00:10:40.46" />
                    <SPLIT distance="1000" swimtime="00:11:51.98" />
                    <SPLIT distance="1100" swimtime="00:13:03.51" />
                    <SPLIT distance="1200" swimtime="00:14:15.34" />
                    <SPLIT distance="1300" swimtime="00:15:27.16" />
                    <SPLIT distance="1400" swimtime="00:16:38.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="607" swimtime="00:09:32.39" resultid="2889" heatid="4428" lane="5" entrytime="00:09:27.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.25" />
                    <SPLIT distance="200" swimtime="00:02:19.80" />
                    <SPLIT distance="300" swimtime="00:03:31.54" />
                    <SPLIT distance="400" swimtime="00:04:43.89" />
                    <SPLIT distance="500" swimtime="00:05:56.37" />
                    <SPLIT distance="600" swimtime="00:07:08.70" />
                    <SPLIT distance="700" swimtime="00:08:21.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="589" swimtime="00:04:40.66" resultid="2890" heatid="4510" lane="3" entrytime="00:04:38.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.10" />
                    <SPLIT distance="200" swimtime="00:02:19.28" />
                    <SPLIT distance="300" swimtime="00:03:30.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Pellanda" birthdate="2010-11-12" gender="M" nation="BRA" license="356352" swrid="5600233" athleteid="2694" externalid="356352">
              <RESULTS>
                <RESULT eventid="1124" points="554" swimtime="00:09:10.38" resultid="2695" heatid="4313" lane="6" entrytime="00:09:15.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.83" />
                    <SPLIT distance="200" swimtime="00:02:12.73" />
                    <SPLIT distance="300" swimtime="00:03:22.36" />
                    <SPLIT distance="400" swimtime="00:04:31.73" />
                    <SPLIT distance="500" swimtime="00:05:41.96" />
                    <SPLIT distance="600" swimtime="00:06:52.22" />
                    <SPLIT distance="700" swimtime="00:08:02.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="487" swimtime="00:00:59.56" resultid="2696" heatid="4344" lane="2" entrytime="00:00:59.88" entrycourse="LCM" />
                <RESULT eventid="1258" points="551" swimtime="00:17:41.93" resultid="2697" heatid="4432" lane="5" entrytime="00:18:12.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.90" />
                    <SPLIT distance="200" swimtime="00:02:15.98" />
                    <SPLIT distance="300" swimtime="00:03:26.66" />
                    <SPLIT distance="400" swimtime="00:04:37.61" />
                    <SPLIT distance="500" swimtime="00:05:48.99" />
                    <SPLIT distance="600" swimtime="00:07:00.27" />
                    <SPLIT distance="700" swimtime="00:08:11.99" />
                    <SPLIT distance="800" swimtime="00:09:23.05" />
                    <SPLIT distance="900" swimtime="00:10:34.45" />
                    <SPLIT distance="1000" swimtime="00:11:45.88" />
                    <SPLIT distance="1100" swimtime="00:12:56.62" />
                    <SPLIT distance="1200" swimtime="00:14:07.77" />
                    <SPLIT distance="1300" swimtime="00:15:18.93" />
                    <SPLIT distance="1400" swimtime="00:16:32.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1274" status="DSQ" swimtime="00:02:32.89" resultid="2698" heatid="4445" lane="7" entrytime="00:02:44.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="361" swimtime="00:01:12.43" resultid="2699" heatid="4529" lane="1" entrytime="00:01:13.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diego" lastname="Rafael Faria Vellozo" birthdate="2008-02-21" gender="M" nation="BRA" license="342231" swrid="5600239" athleteid="2596" externalid="342231">
              <RESULTS>
                <RESULT eventid="1072" points="374" swimtime="00:02:35.32" resultid="2597" heatid="4275" lane="4" entrytime="00:02:30.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1306" points="438" swimtime="00:00:31.00" resultid="2598" heatid="4480" lane="4" entrytime="00:00:32.06" entrycourse="LCM" />
                <RESULT eventid="1374" points="438" swimtime="00:01:07.93" resultid="2599" heatid="4531" lane="5" entrytime="00:01:07.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Albuquerque" birthdate="2008-03-14" gender="F" nation="BRA" license="324787" swrid="5315259" athleteid="2445" externalid="324787">
              <RESULTS>
                <RESULT eventid="1080" points="516" swimtime="00:02:51.39" resultid="2446" heatid="4282" lane="3" entrytime="00:02:48.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="523" swimtime="00:01:19.55" resultid="2447" heatid="4384" lane="3" entrytime="00:01:16.67" entrycourse="LCM" />
                <RESULT eventid="1266" points="494" swimtime="00:02:39.45" resultid="2448" heatid="4434" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Guimaraes E Souza" birthdate="2008-12-21" gender="M" nation="BRA" license="376972" swrid="5600182" athleteid="2891" externalid="376972">
              <RESULTS>
                <RESULT eventid="1088" points="441" swimtime="00:02:44.76" resultid="2892" heatid="4288" lane="2" entrytime="00:02:41.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="522" swimtime="00:00:32.22" resultid="2893" heatid="4368" lane="7" entrytime="00:00:33.70" entrycourse="LCM" />
                <RESULT eventid="1220" points="490" swimtime="00:01:12.11" resultid="2894" heatid="4393" lane="4" entrytime="00:01:12.45" entrycourse="LCM" />
                <RESULT eventid="1274" points="437" swimtime="00:02:30.16" resultid="2895" heatid="4446" lane="3" entrytime="00:02:32.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Kremer De Aguiar" birthdate="2009-12-22" gender="F" nation="BRA" license="338987" swrid="5600196" athleteid="2615" externalid="338987">
              <RESULTS>
                <RESULT eventid="1080" points="414" swimtime="00:03:04.47" resultid="2616" heatid="4281" lane="2" entrytime="00:03:03.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="412" swimtime="00:00:39.17" resultid="2617" heatid="4358" lane="7" entrytime="00:00:40.30" entrycourse="LCM" />
                <RESULT eventid="1212" points="412" swimtime="00:01:26.16" resultid="2618" heatid="4383" lane="1" entrytime="00:01:25.14" entrycourse="LCM" />
                <RESULT eventid="1266" points="428" swimtime="00:02:47.29" resultid="2619" heatid="4438" lane="3" entrytime="00:02:49.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Fontana" birthdate="2011-12-29" gender="M" nation="BRA" license="366897" swrid="5602539" athleteid="2781" externalid="366897">
              <RESULTS>
                <RESULT eventid="1088" points="184" swimtime="00:03:40.54" resultid="2782" heatid="4284" lane="3" entrytime="00:03:44.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="166" swimtime="00:01:43.47" resultid="2783" heatid="4387" lane="6" entrytime="00:01:46.55" entrycourse="LCM" />
                <RESULT eventid="1236" points="224" swimtime="00:00:34.38" resultid="2784" heatid="4411" lane="7" entrytime="00:00:35.48" entrycourse="LCM" />
                <RESULT eventid="1342" points="154" swimtime="00:01:32.09" resultid="2785" heatid="4498" lane="5" />
                <RESULT eventid="1374" points="175" swimtime="00:01:32.11" resultid="2786" heatid="4526" lane="5" entrytime="00:01:32.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia" lastname="Salesi Chicon" birthdate="2002-04-16" gender="F" nation="BRA" license="250865" swrid="5600255" athleteid="2934" externalid="250865">
              <RESULTS>
                <RESULT eventid="1116" points="678" swimtime="00:17:27.57" resultid="2935" heatid="4309" lane="4" entrytime="00:17:23.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.92" />
                    <SPLIT distance="200" swimtime="00:02:16.86" />
                    <SPLIT distance="300" swimtime="00:03:26.88" />
                    <SPLIT distance="400" swimtime="00:04:37.51" />
                    <SPLIT distance="500" swimtime="00:05:47.58" />
                    <SPLIT distance="600" swimtime="00:06:57.79" />
                    <SPLIT distance="700" swimtime="00:08:07.77" />
                    <SPLIT distance="800" swimtime="00:09:18.17" />
                    <SPLIT distance="900" swimtime="00:10:28.10" />
                    <SPLIT distance="1000" swimtime="00:11:38.10" />
                    <SPLIT distance="1100" swimtime="00:12:48.30" />
                    <SPLIT distance="1200" swimtime="00:13:58.37" />
                    <SPLIT distance="1300" swimtime="00:15:09.06" />
                    <SPLIT distance="1400" swimtime="00:16:19.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="609" swimtime="00:05:13.65" resultid="2936" heatid="4315" lane="4" entrytime="00:05:16.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.96" />
                    <SPLIT distance="200" swimtime="00:02:36.76" />
                    <SPLIT distance="300" swimtime="00:04:06.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="693" swimtime="00:09:07.74" resultid="2937" heatid="4428" lane="4" entrytime="00:09:04.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.74" />
                    <SPLIT distance="200" swimtime="00:02:13.17" />
                    <SPLIT distance="300" swimtime="00:03:22.45" />
                    <SPLIT distance="400" swimtime="00:04:31.31" />
                    <SPLIT distance="500" swimtime="00:05:40.92" />
                    <SPLIT distance="600" swimtime="00:06:50.51" />
                    <SPLIT distance="700" swimtime="00:08:00.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="755" swimtime="00:02:03.91" resultid="2938" heatid="4457" lane="4" entrytime="00:02:05.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="721" swimtime="00:04:22.46" resultid="2939" heatid="4510" lane="4" entrytime="00:04:20.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.88" />
                    <SPLIT distance="200" swimtime="00:02:09.38" />
                    <SPLIT distance="300" swimtime="00:03:16.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Zaroni" birthdate="2010-03-03" gender="F" nation="BRA" license="356345" swrid="5600282" athleteid="2526" externalid="356345">
              <RESULTS>
                <RESULT eventid="1080" points="452" swimtime="00:02:59.16" resultid="2527" heatid="4282" lane="7" entrytime="00:02:56.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="488" swimtime="00:01:05.65" resultid="2528" heatid="4327" lane="6" entrytime="00:01:07.86" entrycourse="LCM" />
                <RESULT eventid="1212" points="444" swimtime="00:01:24.05" resultid="2529" heatid="4384" lane="1" entrytime="00:01:21.40" entrycourse="LCM" />
                <RESULT eventid="1266" points="421" swimtime="00:02:48.24" resultid="2530" heatid="4438" lane="6" entrytime="00:02:52.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="4970" points="457" swimtime="00:01:23.24" resultid="4976" heatid="4972" lane="5" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Fontes Hoshina" birthdate="2008-02-15" gender="M" nation="BRA" license="369445" swrid="5600165" athleteid="2489" externalid="369445">
              <RESULTS>
                <RESULT eventid="1104" points="554" swimtime="00:00:27.10" resultid="2490" heatid="4304" lane="1" entrytime="00:00:27.16" entrycourse="LCM" />
                <RESULT eventid="1172" points="509" swimtime="00:02:18.18" resultid="2491" heatid="4351" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1274" points="562" swimtime="00:02:18.08" resultid="2492" heatid="4447" lane="5" entrytime="00:02:18.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="592" swimtime="00:00:58.87" resultid="2493" heatid="4505" lane="8" entrytime="00:01:00.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Clivatti" birthdate="2010-05-24" gender="M" nation="BRA" license="368007" swrid="5600139" athleteid="2845" externalid="368007">
              <RESULTS>
                <RESULT eventid="1124" points="482" swimtime="00:09:36.43" resultid="2846" heatid="4312" lane="5" entrytime="00:09:46.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.82" />
                    <SPLIT distance="200" swimtime="00:02:18.27" />
                    <SPLIT distance="300" swimtime="00:03:30.91" />
                    <SPLIT distance="400" swimtime="00:04:43.87" />
                    <SPLIT distance="500" swimtime="00:05:57.32" />
                    <SPLIT distance="600" swimtime="00:07:11.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="498" swimtime="00:00:59.09" resultid="2847" heatid="4344" lane="6" entrytime="00:00:59.82" entrycourse="LCM" />
                <RESULT eventid="1236" points="451" swimtime="00:00:27.25" resultid="2848" heatid="4417" lane="1" entrytime="00:00:27.57" entrycourse="LCM" />
                <RESULT eventid="1290" points="509" swimtime="00:02:07.68" resultid="2849" heatid="4467" lane="3" entrytime="00:02:09.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="501" swimtime="00:04:37.03" resultid="2850" heatid="4515" lane="3" entrytime="00:04:40.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.17" />
                    <SPLIT distance="200" swimtime="00:02:12.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Prosdocimo" birthdate="2010-11-23" gender="F" nation="BRA" license="356251" swrid="5600238" athleteid="2682" externalid="356251">
              <RESULTS>
                <RESULT eventid="1116" points="420" swimtime="00:20:28.62" resultid="2683" heatid="4309" lane="7" entrytime="00:20:44.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.37" />
                    <SPLIT distance="200" swimtime="00:02:37.98" />
                    <SPLIT distance="300" swimtime="00:03:59.01" />
                    <SPLIT distance="400" swimtime="00:05:20.87" />
                    <SPLIT distance="500" swimtime="00:06:42.55" />
                    <SPLIT distance="600" swimtime="00:08:03.86" />
                    <SPLIT distance="700" swimtime="00:09:25.82" />
                    <SPLIT distance="800" swimtime="00:10:48.07" />
                    <SPLIT distance="900" swimtime="00:12:10.90" />
                    <SPLIT distance="1000" swimtime="00:13:33.38" />
                    <SPLIT distance="1100" swimtime="00:14:57.80" />
                    <SPLIT distance="1200" swimtime="00:16:21.53" />
                    <SPLIT distance="1300" swimtime="00:17:45.49" />
                    <SPLIT distance="1400" swimtime="00:19:08.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="493" swimtime="00:01:05.45" resultid="2684" heatid="4328" lane="8" entrytime="00:01:06.84" entrycourse="LCM" />
                <RESULT eventid="1250" points="422" swimtime="00:10:46.21" resultid="2685" heatid="4428" lane="9" entrytime="00:10:34.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.11" />
                    <SPLIT distance="200" swimtime="00:02:37.52" />
                    <SPLIT distance="300" swimtime="00:04:00.24" />
                    <SPLIT distance="400" swimtime="00:05:22.38" />
                    <SPLIT distance="500" swimtime="00:06:44.94" />
                    <SPLIT distance="600" swimtime="00:08:07.21" />
                    <SPLIT distance="700" swimtime="00:09:28.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="416" swimtime="00:01:16.79" resultid="2686" heatid="4523" lane="3" entrytime="00:01:16.78" entrycourse="LCM" />
                <RESULT eventid="1350" points="427" swimtime="00:05:12.52" resultid="2687" heatid="4509" lane="2" entrytime="00:05:08.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.43" />
                    <SPLIT distance="200" swimtime="00:02:34.59" />
                    <SPLIT distance="300" swimtime="00:03:54.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Geremia" birthdate="2011-07-20" gender="F" nation="BRA" license="366908" swrid="5602543" athleteid="2823" externalid="366908">
              <RESULTS>
                <RESULT eventid="1064" points="463" swimtime="00:02:39.16" resultid="2824" heatid="4270" lane="2" entrytime="00:02:47.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="488" swimtime="00:01:05.65" resultid="2825" heatid="4328" lane="7" entrytime="00:01:06.33" entrycourse="LCM" />
                <RESULT eventid="1250" points="446" swimtime="00:10:34.48" resultid="2826" heatid="4428" lane="0" entrytime="00:10:28.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.76" />
                    <SPLIT distance="200" swimtime="00:02:33.79" />
                    <SPLIT distance="300" swimtime="00:03:54.46" />
                    <SPLIT distance="400" swimtime="00:05:15.26" />
                    <SPLIT distance="500" swimtime="00:06:35.95" />
                    <SPLIT distance="600" swimtime="00:07:56.70" />
                    <SPLIT distance="700" swimtime="00:09:16.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" points="438" swimtime="00:02:46.01" resultid="2827" heatid="4438" lane="1" entrytime="00:02:55.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="456" swimtime="00:05:05.72" resultid="2828" heatid="4509" lane="7" entrytime="00:05:09.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.89" />
                    <SPLIT distance="200" swimtime="00:02:33.01" />
                    <SPLIT distance="300" swimtime="00:03:50.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gael" lastname="Gluck" birthdate="2011-01-28" gender="M" nation="BRA" license="366891" swrid="5588726" athleteid="2763" externalid="366891">
              <RESULTS>
                <RESULT eventid="1088" points="331" swimtime="00:03:01.30" resultid="2764" heatid="4285" lane="4" entrytime="00:03:03.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="377" swimtime="00:01:04.84" resultid="2765" heatid="4339" lane="5" entrytime="00:01:06.61" entrycourse="LCM" />
                <RESULT eventid="1188" points="327" swimtime="00:00:37.64" resultid="2766" heatid="4365" lane="6" entrytime="00:00:39.86" entrycourse="LCM" />
                <RESULT eventid="1220" points="335" swimtime="00:01:21.82" resultid="2767" heatid="4390" lane="6" entrytime="00:01:24.43" entrycourse="LCM" />
                <RESULT eventid="1358" points="373" swimtime="00:05:05.57" resultid="2768" heatid="4514" lane="8" entrytime="00:05:10.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.48" />
                    <SPLIT distance="200" swimtime="00:02:31.88" />
                    <SPLIT distance="300" swimtime="00:03:50.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Braun Prado" birthdate="2008-04-07" gender="M" nation="BRA" license="307663" swrid="5484324" athleteid="2641" externalid="307663">
              <RESULTS>
                <RESULT eventid="1072" points="493" swimtime="00:02:21.62" resultid="2642" heatid="4277" lane="1" entrytime="00:02:19.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="537" swimtime="00:00:57.65" resultid="2643" heatid="4344" lane="3" entrytime="00:00:59.80" entrycourse="LCM" />
                <RESULT eventid="1236" points="454" swimtime="00:00:27.20" resultid="2644" heatid="4409" lane="6" />
                <RESULT eventid="1306" points="489" swimtime="00:00:29.88" resultid="2645" heatid="4476" lane="6" />
                <RESULT eventid="1374" points="517" swimtime="00:01:04.25" resultid="2646" heatid="4532" lane="6" entrytime="00:01:03.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nina" lastname="Rocha Ribeiro Da Silva" birthdate="2010-09-22" gender="F" nation="BRA" license="367216" swrid="5588884" athleteid="2916" externalid="367216">
              <RESULTS>
                <RESULT eventid="1080" points="401" swimtime="00:03:06.41" resultid="2917" heatid="4281" lane="6" entrytime="00:03:03.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="419" swimtime="00:01:09.05" resultid="2918" heatid="4326" lane="6" entrytime="00:01:09.78" entrycourse="LCM" />
                <RESULT eventid="1180" points="464" swimtime="00:00:37.64" resultid="2919" heatid="4358" lane="1" entrytime="00:00:41.02" entrycourse="LCM" />
                <RESULT eventid="1212" points="424" swimtime="00:01:25.33" resultid="2920" heatid="4383" lane="6" entrytime="00:01:23.50" entrycourse="LCM" />
                <RESULT eventid="1282" points="360" swimtime="00:02:38.57" resultid="2921" heatid="4454" lane="2" entrytime="00:02:32.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Novak Bredt" birthdate="2009-09-08" gender="F" nation="BRA" license="338909" swrid="5622297" athleteid="2531" externalid="338909">
              <RESULTS>
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="2532" heatid="4282" lane="1" entrytime="00:02:58.10" entrycourse="LCM" />
                <RESULT eventid="1180" status="DNS" swimtime="00:00:00.00" resultid="2533" heatid="4359" lane="1" entrytime="00:00:38.07" entrycourse="LCM" />
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="2534" heatid="4384" lane="7" entrytime="00:01:21.28" entrycourse="LCM" />
                <RESULT eventid="1266" status="DNS" swimtime="00:00:00.00" resultid="2535" heatid="4439" lane="1" entrytime="00:02:42.47" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Fontolan Gomes" birthdate="2010-07-02" gender="M" nation="BRA" license="356245" swrid="5588705" athleteid="2664" externalid="356245">
              <RESULTS>
                <RESULT eventid="1072" points="374" swimtime="00:02:35.27" resultid="2665" heatid="4275" lane="8" entrytime="00:02:36.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="354" swimtime="00:01:06.24" resultid="2666" heatid="4339" lane="3" entrytime="00:01:06.79" entrycourse="LCM" />
                <RESULT eventid="1290" points="366" swimtime="00:02:22.53" resultid="2667" heatid="4463" lane="7" entrytime="00:02:27.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="384" swimtime="00:05:02.63" resultid="2668" heatid="4513" lane="2" entrytime="00:05:17.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.42" />
                    <SPLIT distance="200" swimtime="00:02:29.60" />
                    <SPLIT distance="300" swimtime="00:03:47.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="351" swimtime="00:01:13.11" resultid="2669" heatid="4529" lane="5" entrytime="00:01:12.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Brandt De Macedo" birthdate="2010-01-13" gender="M" nation="BRA" license="338925" swrid="5588565" athleteid="2740" externalid="338925">
              <RESULTS>
                <RESULT eventid="1124" points="449" swimtime="00:09:50.38" resultid="2741" heatid="4313" lane="8" entrytime="00:09:34.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.61" />
                    <SPLIT distance="200" swimtime="00:02:17.52" />
                    <SPLIT distance="300" swimtime="00:03:31.44" />
                    <SPLIT distance="400" swimtime="00:04:46.20" />
                    <SPLIT distance="500" swimtime="00:06:01.99" />
                    <SPLIT distance="600" swimtime="00:07:18.56" />
                    <SPLIT distance="700" swimtime="00:08:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="455" swimtime="00:01:00.90" resultid="2742" heatid="4342" lane="4" entrytime="00:01:01.92" entrycourse="LCM" />
                <RESULT eventid="1258" points="457" swimtime="00:18:50.77" resultid="2743" heatid="4432" lane="3" entrytime="00:18:23.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.08" />
                    <SPLIT distance="200" swimtime="00:02:20.67" />
                    <SPLIT distance="300" swimtime="00:03:35.11" />
                    <SPLIT distance="400" swimtime="00:04:50.40" />
                    <SPLIT distance="500" swimtime="00:06:05.65" />
                    <SPLIT distance="600" swimtime="00:07:21.30" />
                    <SPLIT distance="700" swimtime="00:08:37.47" />
                    <SPLIT distance="800" swimtime="00:09:53.56" />
                    <SPLIT distance="900" swimtime="00:11:10.17" />
                    <SPLIT distance="1000" swimtime="00:12:26.56" />
                    <SPLIT distance="1100" swimtime="00:13:43.30" />
                    <SPLIT distance="1200" swimtime="00:15:00.35" />
                    <SPLIT distance="1300" swimtime="00:16:17.45" />
                    <SPLIT distance="1400" swimtime="00:17:34.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="455" swimtime="00:02:12.53" resultid="2744" heatid="4466" lane="7" entrytime="00:02:14.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="455" swimtime="00:04:45.97" resultid="2745" heatid="4515" lane="5" entrytime="00:04:40.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.24" />
                    <SPLIT distance="200" swimtime="00:02:19.75" />
                    <SPLIT distance="300" swimtime="00:03:33.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Braga Amatuzzi" birthdate="2006-01-18" gender="M" nation="BRA" license="296650" swrid="5465902" athleteid="2513" externalid="296650">
              <RESULTS>
                <RESULT eventid="1088" points="684" swimtime="00:02:22.37" resultid="2514" heatid="4289" lane="5" entrytime="00:02:16.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="638" swimtime="00:00:30.14" resultid="2515" heatid="4369" lane="2" entrytime="00:00:29.37" entrycourse="LCM" />
                <RESULT eventid="1220" points="605" swimtime="00:01:07.23" resultid="2516" heatid="4395" lane="3" entrytime="00:01:03.51" entrycourse="LCM" />
                <RESULT eventid="1290" points="664" swimtime="00:01:56.87" resultid="2517" heatid="4458" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Peret Saboia" birthdate="2009-11-25" gender="F" nation="BRA" license="342238" swrid="5600234" athleteid="2610" externalid="342238">
              <RESULTS>
                <RESULT eventid="1080" points="457" swimtime="00:02:58.57" resultid="2611" heatid="4281" lane="3" entrytime="00:03:03.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="473" swimtime="00:00:37.40" resultid="2612" heatid="4359" lane="7" entrytime="00:00:38.04" entrycourse="LCM" />
                <RESULT eventid="1212" points="476" swimtime="00:01:22.09" resultid="2613" heatid="4383" lane="4" entrytime="00:01:21.98" entrycourse="LCM" />
                <RESULT eventid="1266" points="415" swimtime="00:02:48.98" resultid="2614" heatid="4438" lane="4" entrytime="00:02:48.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo" lastname="De Lima Cavalcanti" birthdate="2009-12-17" gender="M" nation="BRA" license="380965" swrid="5634589" athleteid="2969" externalid="380965">
              <RESULTS>
                <RESULT eventid="1104" points="518" swimtime="00:00:27.72" resultid="2970" heatid="4301" lane="1" entrytime="00:00:30.28" entrycourse="LCM" />
                <RESULT eventid="1172" points="423" swimtime="00:02:26.98" resultid="2971" heatid="4353" lane="5" entrytime="00:02:25.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="504" swimtime="00:00:26.27" resultid="2972" heatid="4419" lane="1" entrytime="00:00:26.60" entrycourse="LCM" />
                <RESULT eventid="1342" points="491" swimtime="00:01:02.65" resultid="2973" heatid="4504" lane="3" entrytime="00:01:01.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carol" lastname="De Hertel" birthdate="2001-02-20" gender="F" nation="BRA" license="118424" athleteid="3002" externalid="118424">
              <RESULTS>
                <RESULT eventid="1116" status="DNS" swimtime="00:00:00.00" resultid="3003" heatid="4308" lane="3" entrytime="00:22:41.00" entrycourse="LCM" />
                <RESULT eventid="1250" points="618" swimtime="00:09:28.86" resultid="3004" heatid="4426" lane="1" entrytime="00:11:57.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.34" />
                    <SPLIT distance="200" swimtime="00:02:15.29" />
                    <SPLIT distance="300" swimtime="00:03:26.52" />
                    <SPLIT distance="400" swimtime="00:04:38.51" />
                    <SPLIT distance="500" swimtime="00:05:51.23" />
                    <SPLIT distance="600" swimtime="00:07:04.27" />
                    <SPLIT distance="700" swimtime="00:08:17.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="570" swimtime="00:04:43.74" resultid="3005" heatid="4506" lane="4" entrytime="00:05:46.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.59" />
                    <SPLIT distance="200" swimtime="00:02:17.62" />
                    <SPLIT distance="300" swimtime="00:03:30.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Valduga Artigas" birthdate="2009-06-01" gender="M" nation="BRA" license="339569" swrid="5600268" athleteid="2631" externalid="339569">
              <RESULTS>
                <RESULT eventid="1104" points="319" swimtime="00:00:32.57" resultid="2632" heatid="4298" lane="5" entrytime="00:00:36.27" entrycourse="LCM" />
                <RESULT eventid="1156" points="351" swimtime="00:01:06.37" resultid="2633" heatid="4340" lane="3" entrytime="00:01:05.80" entrycourse="LCM" />
                <RESULT eventid="1342" points="262" swimtime="00:01:17.25" resultid="2634" heatid="4501" lane="7" entrytime="00:01:15.33" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Felipe Paes Feres" birthdate="2008-07-28" gender="M" nation="BRA" license="307676" swrid="5600156" athleteid="2575" externalid="307676">
              <RESULTS>
                <RESULT eventid="1072" points="437" swimtime="00:02:27.45" resultid="2576" heatid="4276" lane="2" entrytime="00:02:28.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="477" swimtime="00:00:59.94" resultid="2577" heatid="4345" lane="3" entrytime="00:00:59.08" entrycourse="LCM" />
                <RESULT eventid="1236" points="460" swimtime="00:00:27.07" resultid="2578" heatid="4419" lane="7" entrytime="00:00:26.51" entrycourse="LCM" />
                <RESULT eventid="1306" points="406" swimtime="00:00:31.79" resultid="2579" heatid="4481" lane="1" entrytime="00:00:31.61" entrycourse="LCM" />
                <RESULT eventid="1374" points="428" swimtime="00:01:08.47" resultid="2580" heatid="4532" lane="1" entrytime="00:01:06.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Estevao" lastname="Valduga Artigas" birthdate="2009-06-01" gender="M" nation="BRA" license="339556" swrid="5600267" athleteid="2600" externalid="339556">
              <RESULTS>
                <RESULT eventid="1072" points="281" swimtime="00:02:50.77" resultid="2601" heatid="4273" lane="1" entrytime="00:03:25.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="340" swimtime="00:10:47.70" resultid="2602" heatid="4311" lane="7" entrytime="00:10:48.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.61" />
                    <SPLIT distance="200" swimtime="00:02:36.79" />
                    <SPLIT distance="300" swimtime="00:03:59.08" />
                    <SPLIT distance="400" swimtime="00:05:21.17" />
                    <SPLIT distance="500" swimtime="00:06:43.69" />
                    <SPLIT distance="600" swimtime="00:08:06.60" />
                    <SPLIT distance="700" swimtime="00:09:29.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="291" swimtime="00:00:31.53" resultid="2603" heatid="4412" lane="7" entrytime="00:00:32.50" entrycourse="LCM" />
                <RESULT eventid="1374" points="274" swimtime="00:01:19.41" resultid="2604" heatid="4528" lane="1" entrytime="00:01:19.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Vieira Motta" birthdate="2009-09-19" gender="M" nation="BRA" license="339064" swrid="5600271" athleteid="2635" externalid="339064">
              <RESULTS>
                <RESULT eventid="1072" points="454" swimtime="00:02:25.61" resultid="2636" heatid="4275" lane="2" entrytime="00:02:33.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="482" swimtime="00:09:36.45" resultid="2637" heatid="4312" lane="6" entrytime="00:09:53.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.44" />
                    <SPLIT distance="200" swimtime="00:02:18.59" />
                    <SPLIT distance="300" swimtime="00:03:30.31" />
                    <SPLIT distance="400" swimtime="00:04:43.43" />
                    <SPLIT distance="500" swimtime="00:05:57.14" />
                    <SPLIT distance="600" swimtime="00:07:11.17" />
                    <SPLIT distance="700" swimtime="00:08:25.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="437" swimtime="00:01:01.71" resultid="2638" heatid="4339" lane="7" entrytime="00:01:07.25" entrycourse="LCM" />
                <RESULT eventid="1258" points="461" swimtime="00:18:46.75" resultid="2639" heatid="4432" lane="9" entrytime="00:19:33.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.32" />
                    <SPLIT distance="200" swimtime="00:02:19.63" />
                    <SPLIT distance="300" swimtime="00:03:33.23" />
                    <SPLIT distance="400" swimtime="00:04:47.89" />
                    <SPLIT distance="500" swimtime="00:06:03.37" />
                    <SPLIT distance="600" swimtime="00:07:19.46" />
                    <SPLIT distance="700" swimtime="00:08:35.62" />
                    <SPLIT distance="800" swimtime="00:09:52.42" />
                    <SPLIT distance="900" swimtime="00:11:09.09" />
                    <SPLIT distance="1000" swimtime="00:12:25.89" />
                    <SPLIT distance="1100" swimtime="00:13:42.42" />
                    <SPLIT distance="1200" swimtime="00:14:59.92" />
                    <SPLIT distance="1300" swimtime="00:16:17.50" />
                    <SPLIT distance="1400" swimtime="00:17:33.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="457" swimtime="00:01:06.98" resultid="2640" heatid="4530" lane="4" entrytime="00:01:09.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariana" lastname="Stoberl" birthdate="2010-07-09" gender="F" nation="BRA" license="356250" swrid="5600265" athleteid="2676" externalid="356250">
              <RESULTS>
                <RESULT eventid="1148" points="510" swimtime="00:01:04.68" resultid="2677" heatid="4329" lane="5" entrytime="00:01:04.05" entrycourse="LCM" />
                <RESULT eventid="1228" points="534" swimtime="00:00:29.09" resultid="2678" heatid="4404" lane="3" entrytime="00:00:29.58" entrycourse="LCM" />
                <RESULT eventid="1282" points="509" swimtime="00:02:21.33" resultid="2679" heatid="4456" lane="6" entrytime="00:02:20.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="314" swimtime="00:01:21.55" resultid="2680" heatid="4494" lane="8" />
                <RESULT eventid="1350" points="465" swimtime="00:05:03.77" resultid="2681" heatid="4509" lane="6" entrytime="00:05:07.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.42" />
                    <SPLIT distance="200" swimtime="00:02:32.18" />
                    <SPLIT distance="300" swimtime="00:03:50.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Clara Fernandes Pereira" birthdate="2009-11-19" gender="F" nation="BRA" license="344340" swrid="5600137" athleteid="2449" externalid="344340">
              <RESULTS>
                <RESULT eventid="1132" points="460" swimtime="00:05:44.29" resultid="2450" heatid="4315" lane="5" entrytime="00:05:42.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.62" />
                    <SPLIT distance="200" swimtime="00:02:46.01" />
                    <SPLIT distance="300" swimtime="00:04:26.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="540" swimtime="00:09:55.28" resultid="2451" heatid="4428" lane="7" entrytime="00:10:05.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.20" />
                    <SPLIT distance="200" swimtime="00:02:26.26" />
                    <SPLIT distance="300" swimtime="00:03:41.22" />
                    <SPLIT distance="400" swimtime="00:04:56.42" />
                    <SPLIT distance="500" swimtime="00:06:11.42" />
                    <SPLIT distance="600" swimtime="00:07:26.64" />
                    <SPLIT distance="700" swimtime="00:08:41.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="551" swimtime="00:02:17.57" resultid="2452" heatid="4456" lane="4" entrytime="00:02:17.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="533" swimtime="00:04:50.27" resultid="2453" heatid="4510" lane="1" entrytime="00:04:49.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.46" />
                    <SPLIT distance="200" swimtime="00:02:21.66" />
                    <SPLIT distance="300" swimtime="00:03:36.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Emili Da Silva Gomes Xavier" birthdate="2010-09-08" gender="F" nation="BRA" license="372519" swrid="5717260" athleteid="2992" externalid="372519">
              <RESULTS>
                <RESULT eventid="1064" points="341" swimtime="00:02:56.11" resultid="2993" heatid="4269" lane="6" entrytime="00:02:57.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="417" swimtime="00:00:31.58" resultid="2994" heatid="4402" lane="7" entrytime="00:00:31.29" entrycourse="LCM" />
                <RESULT eventid="1212" points="402" swimtime="00:01:26.83" resultid="2995" heatid="4381" lane="5" entrytime="00:01:30.91" entrycourse="LCM" />
                <RESULT eventid="1282" points="417" swimtime="00:02:30.95" resultid="2996" heatid="4453" lane="7" entrytime="00:02:35.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="336" swimtime="00:01:22.44" resultid="2997" heatid="4521" lane="2" entrytime="00:01:22.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Ramos Marcon" birthdate="2008-01-12" gender="M" nation="BRA" license="372281" swrid="5600240" athleteid="2911" externalid="372281">
              <RESULTS>
                <RESULT eventid="1104" points="438" swimtime="00:00:29.32" resultid="2912" heatid="4301" lane="6" entrytime="00:00:29.86" entrycourse="LCM" />
                <RESULT eventid="1156" points="583" swimtime="00:00:56.08" resultid="2913" heatid="4346" lane="4" entrytime="00:00:56.51" entrycourse="LCM" />
                <RESULT eventid="1236" points="542" swimtime="00:00:25.64" resultid="2914" heatid="4420" lane="3" entrytime="00:00:25.53" entrycourse="LCM" />
                <RESULT eventid="1290" points="498" swimtime="00:02:08.62" resultid="2915" heatid="4467" lane="2" entrytime="00:02:09.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Saboia" birthdate="2009-01-25" gender="M" nation="BRA" license="342252" swrid="5600253" athleteid="2620" externalid="342252">
              <RESULTS>
                <RESULT eventid="1088" points="429" swimtime="00:02:46.30" resultid="2621" heatid="4287" lane="6" entrytime="00:02:47.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="456" swimtime="00:00:33.71" resultid="2622" heatid="4365" lane="5" entrytime="00:00:37.74" entrycourse="LCM" />
                <RESULT eventid="1220" points="420" swimtime="00:01:15.92" resultid="2623" heatid="4393" lane="8" entrytime="00:01:15.70" entrycourse="LCM" />
                <RESULT eventid="1274" points="401" swimtime="00:02:34.59" resultid="2624" heatid="4445" lane="4" entrytime="00:02:38.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Estela" lastname="Albuquerque" birthdate="2010-11-23" gender="F" nation="BRA" license="356344" swrid="5653285" athleteid="2688" externalid="356344">
              <RESULTS>
                <RESULT eventid="1064" points="363" swimtime="00:02:52.54" resultid="2689" heatid="4269" lane="5" entrytime="00:02:53.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="456" swimtime="00:01:07.16" resultid="2690" heatid="4326" lane="4" entrytime="00:01:09.04" entrycourse="LCM" />
                <RESULT eventid="1282" points="463" swimtime="00:02:25.79" resultid="2691" heatid="4455" lane="3" entrytime="00:02:27.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="366" swimtime="00:01:20.09" resultid="2692" heatid="4522" lane="3" entrytime="00:01:19.04" entrycourse="LCM" />
                <RESULT eventid="1350" points="428" swimtime="00:05:12.23" resultid="2693" heatid="4508" lane="5" entrytime="00:05:25.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.36" />
                    <SPLIT distance="200" swimtime="00:02:36.75" />
                    <SPLIT distance="300" swimtime="00:03:55.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Sachser Rocha" birthdate="2008-07-09" gender="M" nation="BRA" license="330072" swrid="5600254" athleteid="2581" externalid="330072">
              <RESULTS>
                <RESULT eventid="1104" points="567" swimtime="00:00:26.90" resultid="2582" heatid="4303" lane="7" entrytime="00:00:28.05" entrycourse="LCM" />
                <RESULT eventid="1156" points="542" swimtime="00:00:57.45" resultid="2583" heatid="4346" lane="6" entrytime="00:00:57.34" entrycourse="LCM" />
                <RESULT eventid="1236" points="553" swimtime="00:00:25.46" resultid="2584" heatid="4420" lane="6" entrytime="00:00:25.56" entrycourse="LCM" />
                <RESULT eventid="1342" points="530" swimtime="00:01:01.08" resultid="2585" heatid="4504" lane="1" entrytime="00:01:02.28" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Krupacz" birthdate="2008-04-18" gender="F" nation="BRA" license="329187" swrid="5634611" athleteid="2963" externalid="329187">
              <RESULTS>
                <RESULT eventid="1064" points="537" swimtime="00:02:31.44" resultid="2964" heatid="4271" lane="3" entrytime="00:02:32.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="488" swimtime="00:01:05.66" resultid="2965" heatid="4319" lane="4" />
                <RESULT eventid="1250" status="DNS" swimtime="00:00:00.00" resultid="2966" heatid="4428" lane="1" entrytime="00:10:10.08" entrycourse="LCM" />
                <RESULT eventid="1298" points="606" swimtime="00:00:31.74" resultid="2967" heatid="4470" lane="2" />
                <RESULT eventid="1366" points="564" swimtime="00:01:09.35" resultid="2968" heatid="4524" lane="6" entrytime="00:01:08.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fernandes" birthdate="2010-03-13" gender="M" nation="BRA" license="339266" swrid="5588695" athleteid="2928" externalid="339266">
              <RESULTS>
                <RESULT eventid="1072" points="429" swimtime="00:02:28.36" resultid="2929" heatid="4276" lane="8" entrytime="00:02:30.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="491" swimtime="00:00:59.38" resultid="2930" heatid="4345" lane="7" entrytime="00:00:59.39" entrycourse="LCM" />
                <RESULT eventid="1236" points="466" swimtime="00:00:26.96" resultid="2931" heatid="4418" lane="3" entrytime="00:00:26.94" entrycourse="LCM" />
                <RESULT eventid="1290" points="460" swimtime="00:02:12.08" resultid="2932" heatid="4466" lane="6" entrytime="00:02:14.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="425" swimtime="00:01:08.59" resultid="2933" heatid="4531" lane="8" entrytime="00:01:08.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raphael" lastname="Rached Windmuller" birthdate="2003-05-19" gender="M" nation="BRA" license="249770" swrid="5302329" athleteid="2559" externalid="249770">
              <RESULTS>
                <RESULT eventid="1088" points="804" swimtime="00:02:14.91" resultid="2560" heatid="4289" lane="4" entrytime="00:02:13.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="809" swimtime="00:00:27.84" resultid="2561" heatid="4369" lane="5" entrytime="00:00:27.96" entrycourse="LCM" />
                <RESULT eventid="1220" points="780" swimtime="00:01:01.79" resultid="2562" heatid="4395" lane="4" entrytime="00:01:01.22" entrycourse="LCM" />
                <RESULT eventid="1274" status="DNS" swimtime="00:00:00.00" resultid="2563" heatid="4441" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Pedro Pasqual" birthdate="2009-06-17" gender="M" nation="BRA" license="386136" swrid="5600232" athleteid="3006" externalid="386136">
              <RESULTS>
                <RESULT eventid="1072" points="517" swimtime="00:02:19.42" resultid="3007" heatid="4277" lane="7" entrytime="00:02:19.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="562" swimtime="00:00:56.78" resultid="3008" heatid="4346" lane="1" entrytime="00:00:58.18" entrycourse="LCM" />
                <RESULT eventid="1306" points="557" swimtime="00:00:28.62" resultid="3009" heatid="4481" lane="5" entrytime="00:00:30.25" entrycourse="LCM" />
                <RESULT eventid="1374" status="DSQ" swimtime="00:01:03.85" resultid="3010" heatid="4532" lane="3" entrytime="00:01:03.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Heloisa Souza" birthdate="2007-01-15" gender="F" nation="BRA" license="336615" swrid="5600184" athleteid="2542" externalid="336615">
              <RESULTS>
                <RESULT eventid="1148" points="646" swimtime="00:00:59.80" resultid="2543" heatid="4330" lane="5" entrytime="00:01:00.31" entrycourse="LCM" />
                <RESULT eventid="1250" points="579" swimtime="00:09:41.56" resultid="2544" heatid="4428" lane="3" entrytime="00:09:42.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.47" />
                    <SPLIT distance="200" swimtime="00:02:20.51" />
                    <SPLIT distance="300" swimtime="00:03:32.72" />
                    <SPLIT distance="400" swimtime="00:04:45.87" />
                    <SPLIT distance="500" swimtime="00:05:59.96" />
                    <SPLIT distance="600" swimtime="00:07:13.90" />
                    <SPLIT distance="700" swimtime="00:08:28.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="604" swimtime="00:02:13.50" resultid="2545" heatid="4457" lane="6" entrytime="00:02:11.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="581" swimtime="00:04:41.98" resultid="2546" heatid="4510" lane="7" entrytime="00:04:46.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.57" />
                    <SPLIT distance="200" swimtime="00:02:17.62" />
                    <SPLIT distance="300" swimtime="00:03:29.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Presiazniuk" birthdate="2010-10-14" gender="M" nation="BRA" license="356353" swrid="5600237" athleteid="2700" externalid="356353">
              <RESULTS>
                <RESULT eventid="1072" points="414" swimtime="00:02:30.10" resultid="2701" heatid="4275" lane="6" entrytime="00:02:33.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="469" swimtime="00:01:00.31" resultid="2702" heatid="4343" lane="3" entrytime="00:01:00.66" entrycourse="LCM" />
                <RESULT eventid="1236" points="422" swimtime="00:00:27.86" resultid="2703" heatid="4416" lane="3" entrytime="00:00:27.74" entrycourse="LCM" />
                <RESULT eventid="1290" points="462" swimtime="00:02:11.93" resultid="2704" heatid="4466" lane="2" entrytime="00:02:14.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="399" swimtime="00:01:10.08" resultid="2705" heatid="4530" lane="7" entrytime="00:01:11.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Mattioli" birthdate="2011-10-22" gender="F" nation="BRA" license="366896" swrid="5602559" athleteid="2775" externalid="366896">
              <RESULTS>
                <RESULT eventid="1080" points="378" swimtime="00:03:10.10" resultid="2776" heatid="4280" lane="1" entrytime="00:03:17.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="423" swimtime="00:01:08.88" resultid="2777" heatid="4326" lane="2" entrytime="00:01:09.84" entrycourse="LCM" />
                <RESULT eventid="1212" points="363" swimtime="00:01:29.85" resultid="2778" heatid="4381" lane="3" entrytime="00:01:32.25" entrycourse="LCM" />
                <RESULT eventid="1266" points="399" swimtime="00:02:51.27" resultid="2779" heatid="4437" lane="4" entrytime="00:02:59.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="427" swimtime="00:05:12.40" resultid="2780" heatid="4507" lane="7" entrytime="00:05:46.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.16" />
                    <SPLIT distance="200" swimtime="00:02:34.66" />
                    <SPLIT distance="300" swimtime="00:03:55.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Fontolan Gomes" birthdate="2008-05-01" gender="M" nation="BRA" license="307667" swrid="5600166" athleteid="2570" externalid="307667">
              <RESULTS>
                <RESULT eventid="1072" points="409" swimtime="00:02:30.77" resultid="2571" heatid="4275" lane="3" entrytime="00:02:32.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="422" swimtime="00:00:27.86" resultid="2572" heatid="4407" lane="6" />
                <RESULT eventid="1306" points="379" swimtime="00:00:32.53" resultid="2573" heatid="4480" lane="8" entrytime="00:00:33.52" entrycourse="LCM" />
                <RESULT eventid="1374" points="411" swimtime="00:01:09.36" resultid="2574" heatid="4530" lane="5" entrytime="00:01:09.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1204" points="486" swimtime="00:08:52.13" resultid="3030" heatid="4373" lane="2" entrytime="00:08:16.11">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.35" />
                    <SPLIT distance="200" swimtime="00:02:09.16" />
                    <SPLIT distance="300" swimtime="00:03:13.19" />
                    <SPLIT distance="400" swimtime="00:04:24.24" />
                    <SPLIT distance="500" swimtime="00:05:28.45" />
                    <SPLIT distance="600" swimtime="00:06:39.30" />
                    <SPLIT distance="700" swimtime="00:07:43.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2845" number="1" />
                    <RELAYPOSITION athleteid="2740" number="2" />
                    <RELAYPOSITION athleteid="2928" number="3" />
                    <RELAYPOSITION athleteid="2694" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="19" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1208" points="775" swimtime="00:07:35.59" resultid="3031" heatid="4375" lane="4" entrytime="00:07:43.98">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.33" />
                    <SPLIT distance="200" swimtime="00:01:51.59" />
                    <SPLIT distance="300" swimtime="00:02:46.26" />
                    <SPLIT distance="400" swimtime="00:03:44.44" />
                    <SPLIT distance="500" swimtime="00:04:40.77" />
                    <SPLIT distance="600" swimtime="00:05:40.49" />
                    <SPLIT distance="700" swimtime="00:06:36.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2503" number="1" />
                    <RELAYPOSITION athleteid="2982" number="2" />
                    <RELAYPOSITION athleteid="2513" number="3" />
                    <RELAYPOSITION athleteid="2547" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1206" points="576" swimtime="00:08:22.79" resultid="3032" heatid="4374" lane="7" entrytime="00:08:07.25">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.02" />
                    <SPLIT distance="200" swimtime="00:02:06.60" />
                    <SPLIT distance="300" swimtime="00:03:04.78" />
                    <SPLIT distance="400" swimtime="00:04:14.61" />
                    <SPLIT distance="500" swimtime="00:05:13.16" />
                    <SPLIT distance="600" swimtime="00:06:16.93" />
                    <SPLIT distance="700" swimtime="00:07:16.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2536" number="1" />
                    <RELAYPOSITION athleteid="2957" number="2" />
                    <RELAYPOSITION athleteid="2851" number="3" />
                    <RELAYPOSITION athleteid="2484" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1324" status="DSQ" swimtime="00:04:49.42" resultid="3033" heatid="4488" lane="4" entrytime="00:04:53.52">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.21" />
                    <SPLIT distance="200" swimtime="00:02:31.09" />
                    <SPLIT distance="300" swimtime="00:03:49.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2857" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2763" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="2793" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="2811" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1392" points="402" swimtime="00:04:14.90" resultid="3038" heatid="4539" lane="4" entrytime="00:04:04.42">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.42" />
                    <SPLIT distance="200" swimtime="00:02:04.63" />
                    <SPLIT distance="300" swimtime="00:03:09.31" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2811" number="1" />
                    <RELAYPOSITION athleteid="2857" number="2" />
                    <RELAYPOSITION athleteid="2751" number="3" />
                    <RELAYPOSITION athleteid="2763" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1326" points="410" swimtime="00:04:38.14" resultid="3034" heatid="4489" lane="4" entrytime="00:04:38.22">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.40" />
                    <SPLIT distance="200" swimtime="00:02:28.24" />
                    <SPLIT distance="300" swimtime="00:03:37.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2928" number="1" />
                    <RELAYPOSITION athleteid="2718" number="2" />
                    <RELAYPOSITION athleteid="2694" number="3" />
                    <RELAYPOSITION athleteid="2845" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1394" points="489" swimtime="00:03:58.89" resultid="3039" heatid="4540" lane="4" entrytime="00:03:57.05">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.88" />
                    <SPLIT distance="200" swimtime="00:02:00.21" />
                    <SPLIT distance="300" swimtime="00:03:00.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2658" number="1" />
                    <RELAYPOSITION athleteid="2845" number="2" />
                    <RELAYPOSITION athleteid="2928" number="3" />
                    <RELAYPOSITION athleteid="2694" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1330" points="587" swimtime="00:04:06.95" resultid="3035" heatid="4491" lane="4" entrytime="00:04:09.83">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.50" />
                    <SPLIT distance="200" swimtime="00:02:13.20" />
                    <SPLIT distance="300" swimtime="00:03:12.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2641" number="1" />
                    <RELAYPOSITION athleteid="2494" number="2" />
                    <RELAYPOSITION athleteid="2489" number="3" />
                    <RELAYPOSITION athleteid="2957" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1398" points="608" swimtime="00:03:42.13" resultid="3042" heatid="4542" lane="4" entrytime="00:03:46.37">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:54.55" />
                    <SPLIT distance="200" swimtime="00:01:50.55" />
                    <SPLIT distance="300" swimtime="00:02:45.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2957" number="1" />
                    <RELAYPOSITION athleteid="2851" number="2" />
                    <RELAYPOSITION athleteid="2489" number="3" />
                    <RELAYPOSITION athleteid="2911" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1328" points="519" swimtime="00:04:17.22" resultid="3036" heatid="4490" lane="4" entrytime="00:04:14.43">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.43" />
                    <SPLIT distance="200" swimtime="00:02:19.91" />
                    <SPLIT distance="300" swimtime="00:03:21.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3006" number="1" />
                    <RELAYPOSITION athleteid="2620" number="2" />
                    <RELAYPOSITION athleteid="2969" number="3" />
                    <RELAYPOSITION athleteid="2484" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1396" points="551" swimtime="00:03:49.60" resultid="3041" heatid="4541" lane="4" entrytime="00:03:49.59">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.60" />
                    <SPLIT distance="200" swimtime="00:01:53.40" />
                    <SPLIT distance="300" swimtime="00:02:52.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2484" number="1" />
                    <RELAYPOSITION athleteid="2536" number="2" />
                    <RELAYPOSITION athleteid="3006" number="3" />
                    <RELAYPOSITION athleteid="2969" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1332" points="711" swimtime="00:03:51.59" resultid="3037" heatid="4492" lane="4" entrytime="00:03:57.02">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:56.75" />
                    <SPLIT distance="200" swimtime="00:01:58.89" />
                    <SPLIT distance="300" swimtime="00:02:56.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2834" number="1" />
                    <RELAYPOSITION athleteid="2559" number="2" />
                    <RELAYPOSITION athleteid="2507" number="3" />
                    <RELAYPOSITION athleteid="2547" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1400" points="739" swimtime="00:03:28.16" resultid="3040" heatid="4543" lane="4" entrytime="00:03:39.00">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:50.93" />
                    <SPLIT distance="200" swimtime="00:01:42.51" />
                    <SPLIT distance="300" swimtime="00:02:35.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2547" number="1" />
                    <RELAYPOSITION athleteid="2982" number="2" />
                    <RELAYPOSITION athleteid="2513" number="3" />
                    <RELAYPOSITION athleteid="2503" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1324" points="307" swimtime="00:05:06.31" resultid="3052" heatid="4488" lane="5" entrytime="00:05:10.32">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.43" />
                    <SPLIT distance="200" swimtime="00:02:46.66" />
                    <SPLIT distance="300" swimtime="00:04:01.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2817" number="1" />
                    <RELAYPOSITION athleteid="2896" number="2" />
                    <RELAYPOSITION athleteid="2757" number="3" />
                    <RELAYPOSITION athleteid="2751" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1392" points="322" swimtime="00:04:34.42" resultid="3054" heatid="4539" lane="5" entrytime="00:04:17.28">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.14" />
                    <SPLIT distance="200" swimtime="00:02:15.12" />
                    <SPLIT distance="300" swimtime="00:03:25.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2757" number="1" />
                    <RELAYPOSITION athleteid="2793" number="2" />
                    <RELAYPOSITION athleteid="2817" number="3" />
                    <RELAYPOSITION athleteid="2769" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1326" points="369" swimtime="00:04:48.18" resultid="3053" heatid="4489" lane="6" entrytime="00:04:57.41">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.71" />
                    <SPLIT distance="200" swimtime="00:02:33.07" />
                    <SPLIT distance="300" swimtime="00:03:47.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2700" number="1" />
                    <RELAYPOSITION athleteid="2658" number="2" />
                    <RELAYPOSITION athleteid="2729" number="3" />
                    <RELAYPOSITION athleteid="2740" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1394" points="456" swimtime="00:04:04.56" resultid="3055" heatid="4540" lane="3" entrytime="00:04:26.97">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.68" />
                    <SPLIT distance="200" swimtime="00:02:00.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2718" number="1" />
                    <RELAYPOSITION athleteid="2700" number="2" />
                    <RELAYPOSITION athleteid="2740" number="3" />
                    <RELAYPOSITION athleteid="2706" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1196" points="508" swimtime="00:09:33.12" resultid="3017" heatid="4370" lane="2" entrytime="00:09:07.52">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.53" />
                    <SPLIT distance="200" swimtime="00:02:14.43" />
                    <SPLIT distance="300" swimtime="00:03:24.49" />
                    <SPLIT distance="400" swimtime="00:04:39.12" />
                    <SPLIT distance="500" swimtime="00:05:49.62" />
                    <SPLIT distance="600" swimtime="00:07:06.11" />
                    <SPLIT distance="700" swimtime="00:08:16.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2881" number="1" />
                    <RELAYPOSITION athleteid="2723" number="2" />
                    <RELAYPOSITION athleteid="2682" number="3" />
                    <RELAYPOSITION athleteid="2676" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="19" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1200" points="581" swimtime="00:09:08.09" resultid="3018" heatid="4372" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.14" />
                    <SPLIT distance="200" swimtime="00:02:11.62" />
                    <SPLIT distance="300" swimtime="00:03:19.39" />
                    <SPLIT distance="400" swimtime="00:04:34.19" />
                    <SPLIT distance="500" swimtime="00:05:40.77" />
                    <SPLIT distance="700" swimtime="00:07:58.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2542" number="1" />
                    <RELAYPOSITION athleteid="2978" number="2" />
                    <RELAYPOSITION athleteid="2498" number="3" />
                    <RELAYPOSITION athleteid="2887" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1198" points="556" swimtime="00:09:16.11" resultid="3019" heatid="4371" lane="6" entrytime="00:09:00.98">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.56" />
                    <SPLIT distance="200" swimtime="00:02:14.25" />
                    <SPLIT distance="300" swimtime="00:03:21.05" />
                    <SPLIT distance="400" swimtime="00:04:33.87" />
                    <SPLIT distance="500" swimtime="00:05:40.26" />
                    <SPLIT distance="600" swimtime="00:06:56.01" />
                    <SPLIT distance="700" swimtime="00:08:03.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2520" number="1" />
                    <RELAYPOSITION athleteid="2460" number="2" />
                    <RELAYPOSITION athleteid="2625" number="3" />
                    <RELAYPOSITION athleteid="2449" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1314" points="455" swimtime="00:04:59.39" resultid="3020" heatid="4483" lane="4" entrytime="00:05:09.57">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.85" />
                    <SPLIT distance="200" swimtime="00:02:45.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2823" number="1" />
                    <RELAYPOSITION athleteid="2775" number="2" />
                    <RELAYPOSITION athleteid="2881" number="3" />
                    <RELAYPOSITION athleteid="2805" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1382" points="458" swimtime="00:04:29.62" resultid="3029" heatid="4534" lane="4" entrytime="00:04:27.55">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:02:10.98" />
                    <SPLIT distance="300" swimtime="00:03:22.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2881" number="1" />
                    <RELAYPOSITION athleteid="2805" number="2" />
                    <RELAYPOSITION athleteid="2799" number="3" />
                    <RELAYPOSITION athleteid="2823" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1316" points="452" swimtime="00:05:00.15" resultid="3021" heatid="4484" lane="4" entrytime="00:04:57.86">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.58" />
                    <SPLIT distance="200" swimtime="00:02:39.09" />
                    <SPLIT distance="300" swimtime="00:03:53.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2682" number="1" />
                    <RELAYPOSITION athleteid="2526" number="2" />
                    <RELAYPOSITION athleteid="2723" number="3" />
                    <RELAYPOSITION athleteid="2676" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1384" points="466" swimtime="00:04:28.10" resultid="3027" heatid="4535" lane="4" entrytime="00:04:15.69">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.01" />
                    <SPLIT distance="200" swimtime="00:02:13.94" />
                    <SPLIT distance="300" swimtime="00:03:20.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2676" number="1" />
                    <RELAYPOSITION athleteid="2682" number="2" />
                    <RELAYPOSITION athleteid="2723" number="3" />
                    <RELAYPOSITION athleteid="2526" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1320" points="541" swimtime="00:04:42.72" resultid="3022" heatid="4486" lane="4" entrytime="00:04:45.68">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.31" />
                    <SPLIT distance="200" swimtime="00:02:30.15" />
                    <SPLIT distance="300" swimtime="00:03:38.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2963" number="1" />
                    <RELAYPOSITION athleteid="2445" number="2" />
                    <RELAYPOSITION athleteid="2454" number="3" />
                    <RELAYPOSITION athleteid="2875" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1388" points="536" swimtime="00:04:15.88" resultid="3025" heatid="4537" lane="4" entrytime="00:04:07.97">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.36" />
                    <SPLIT distance="200" swimtime="00:02:09.09" />
                    <SPLIT distance="300" swimtime="00:03:11.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2445" number="1" />
                    <RELAYPOSITION athleteid="2963" number="2" />
                    <RELAYPOSITION athleteid="2454" number="3" />
                    <RELAYPOSITION athleteid="2875" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1318" points="488" swimtime="00:04:52.51" resultid="3023" heatid="4485" lane="1">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:02:39.68" />
                    <SPLIT distance="300" swimtime="00:03:49.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2625" number="1" />
                    <RELAYPOSITION athleteid="2610" number="2" />
                    <RELAYPOSITION athleteid="2520" number="3" />
                    <RELAYPOSITION athleteid="2460" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1386" points="559" swimtime="00:04:12.44" resultid="3028" heatid="4536" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.47" />
                    <SPLIT distance="200" swimtime="00:02:07.24" />
                    <SPLIT distance="300" swimtime="00:03:11.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2460" number="1" />
                    <RELAYPOSITION athleteid="2625" number="2" />
                    <RELAYPOSITION athleteid="2449" number="3" />
                    <RELAYPOSITION athleteid="2520" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1322" points="544" swimtime="00:04:42.19" resultid="3024" heatid="4487" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.88" />
                    <SPLIT distance="200" swimtime="00:02:31.73" />
                    <SPLIT distance="300" swimtime="00:03:40.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2887" number="1" />
                    <RELAYPOSITION athleteid="2978" number="2" />
                    <RELAYPOSITION athleteid="2934" number="3" />
                    <RELAYPOSITION athleteid="2542" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1390" status="WDR" swimtime="00:00:00.00" resultid="3026" heatid="4538" lane="6" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1314" status="DSQ" swimtime="00:05:33.97" resultid="3048" heatid="4483" lane="5" entrytime="00:05:19.58">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:02:56.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2945" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2799" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="2951" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="2869" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1382" points="373" swimtime="00:04:48.87" resultid="3051" heatid="4534" lane="5" entrytime="00:04:37.58">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:02:20.87" />
                    <SPLIT distance="300" swimtime="00:03:34.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2869" number="1" />
                    <RELAYPOSITION athleteid="2775" number="2" />
                    <RELAYPOSITION athleteid="2945" number="3" />
                    <RELAYPOSITION athleteid="2787" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1316" points="387" swimtime="00:05:16.01" resultid="3049" heatid="4484" lane="5" entrytime="00:05:08.42">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:02:43.45" />
                    <SPLIT distance="300" swimtime="00:04:08.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2670" number="1" />
                    <RELAYPOSITION athleteid="2916" number="2" />
                    <RELAYPOSITION athleteid="2735" number="3" />
                    <RELAYPOSITION athleteid="2688" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1384" points="433" swimtime="00:04:34.77" resultid="3050" heatid="4535" lane="5" entrytime="00:04:31.87">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.98" />
                    <SPLIT distance="200" swimtime="00:02:17.53" />
                    <SPLIT distance="300" swimtime="00:03:26.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2688" number="1" />
                    <RELAYPOSITION athleteid="2916" number="2" />
                    <RELAYPOSITION athleteid="2712" number="3" />
                    <RELAYPOSITION athleteid="2992" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1112" points="406" swimtime="00:04:53.76" resultid="3043" heatid="4306" lane="4" entrytime="00:04:55.49">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:02:39.29" />
                    <SPLIT distance="300" swimtime="00:03:52.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2857" number="1" />
                    <RELAYPOSITION athleteid="2775" number="2" />
                    <RELAYPOSITION athleteid="2793" number="3" />
                    <RELAYPOSITION athleteid="2881" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1114" points="454" swimtime="00:04:42.95" resultid="3044" heatid="4307" lane="4" entrytime="00:04:45.86">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.67" />
                    <SPLIT distance="300" swimtime="00:03:44.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2928" number="1" />
                    <RELAYPOSITION athleteid="2916" number="2" />
                    <RELAYPOSITION athleteid="2723" number="3" />
                    <RELAYPOSITION athleteid="2845" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1248" points="571" swimtime="00:04:22.15" resultid="3045" heatid="4425" lane="4" entrytime="00:04:22.85">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.95" />
                    <SPLIT distance="200" swimtime="00:02:19.27" />
                    <SPLIT distance="300" swimtime="00:03:20.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2987" number="1" />
                    <RELAYPOSITION athleteid="2498" number="2" />
                    <RELAYPOSITION athleteid="2553" number="3" />
                    <RELAYPOSITION athleteid="2542" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1246" points="568" swimtime="00:04:22.58" resultid="3046" heatid="4424" lane="4" entrytime="00:04:25.85">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.02" />
                    <SPLIT distance="200" swimtime="00:02:19.48" />
                    <SPLIT distance="300" swimtime="00:03:19.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2963" number="1" />
                    <RELAYPOSITION athleteid="2494" number="2" />
                    <RELAYPOSITION athleteid="2489" number="3" />
                    <RELAYPOSITION athleteid="2445" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1244" points="527" swimtime="00:04:29.28" resultid="3047" heatid="4423" lane="4" entrytime="00:04:31.55">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.58" />
                    <SPLIT distance="200" swimtime="00:02:25.50" />
                    <SPLIT distance="300" swimtime="00:03:26.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3006" number="1" />
                    <RELAYPOSITION athleteid="2610" number="2" />
                    <RELAYPOSITION athleteid="2969" number="3" />
                    <RELAYPOSITION athleteid="2460" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1112" points="354" swimtime="00:05:07.33" resultid="3056" heatid="4306" lane="3" entrytime="00:05:02.39">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.60" />
                    <SPLIT distance="200" swimtime="00:02:43.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2805" number="1" />
                    <RELAYPOSITION athleteid="2811" number="2" />
                    <RELAYPOSITION athleteid="2751" number="3" />
                    <RELAYPOSITION athleteid="2823" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1114" points="407" swimtime="00:04:53.37" resultid="3057" heatid="4307" lane="3" entrytime="00:04:55.20">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.50" />
                    <SPLIT distance="200" swimtime="00:02:32.69" />
                    <SPLIT distance="300" swimtime="00:03:50.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2700" number="1" />
                    <RELAYPOSITION athleteid="2526" number="2" />
                    <RELAYPOSITION athleteid="2718" number="3" />
                    <RELAYPOSITION athleteid="2676" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="16131" nation="BRA" region="PR" clubid="3081" swrid="93766" name="Associação Nadar Colombo" shortname="Equipe Nadar">
          <ATHLETES>
            <ATHLETE firstname="Vitor" lastname="Rafael D Agostin Batistao" birthdate="2008-05-13" gender="M" nation="BRA" license="384738" swrid="5622300" athleteid="3082" externalid="384738">
              <RESULTS>
                <RESULT eventid="1188" points="371" swimtime="00:00:36.11" resultid="3083" heatid="4366" lane="5" entrytime="00:00:36.16" entrycourse="LCM" />
                <RESULT eventid="1220" points="310" swimtime="00:01:24.02" resultid="3084" heatid="4391" lane="1" entrytime="00:01:22.87" entrycourse="LCM" />
                <RESULT eventid="1236" points="315" swimtime="00:00:30.70" resultid="3085" heatid="4414" lane="6" entrytime="00:00:30.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Rosa De Souza" birthdate="2009-01-01" gender="F" nation="BRA" license="399926" swrid="5653301" athleteid="3099" externalid="399926">
              <RESULTS>
                <RESULT eventid="1080" points="191" swimtime="00:03:58.71" resultid="3100" heatid="4278" lane="3" entrytime="00:04:07.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="304" swimtime="00:01:16.90" resultid="3101" heatid="4321" lane="7" entrytime="00:01:25.31" entrycourse="LCM" />
                <RESULT eventid="1212" points="222" swimtime="00:01:45.89" resultid="3102" heatid="4380" lane="8" entrytime="00:01:46.07" entrycourse="LCM" />
                <RESULT eventid="1266" points="219" swimtime="00:03:29.17" resultid="3103" heatid="4435" lane="5" entrytime="00:03:31.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="164" swimtime="00:01:41.17" resultid="3104" heatid="4494" lane="6" entrytime="00:01:57.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Carvalho Ezaki" birthdate="2011-10-20" gender="F" nation="BRA" license="399927" swrid="5652882" athleteid="3105" externalid="399927">
              <RESULTS>
                <RESULT eventid="1180" points="244" swimtime="00:00:46.62" resultid="3106" heatid="4355" lane="6" />
                <RESULT eventid="1212" points="244" swimtime="00:01:42.53" resultid="3107" heatid="4380" lane="2" entrytime="00:01:43.02" entrycourse="LCM" />
                <RESULT eventid="1266" points="235" swimtime="00:03:24.24" resultid="3108" heatid="4435" lane="2" entrytime="00:03:43.63" entrycourse="LCM" />
                <RESULT eventid="1334" points="107" swimtime="00:01:56.67" resultid="3109" heatid="4494" lane="3" entrytime="00:01:45.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Felipe Glir" birthdate="2006-10-11" gender="M" nation="BRA" license="384741" swrid="5622280" athleteid="3090" externalid="384741">
              <RESULTS>
                <RESULT eventid="1104" points="349" swimtime="00:00:31.62" resultid="3091" heatid="4301" lane="7" entrytime="00:00:30.25" entrycourse="LCM" />
                <RESULT eventid="1236" points="404" swimtime="00:00:28.28" resultid="3092" heatid="4418" lane="6" entrytime="00:00:26.96" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Luiz Sartori" birthdate="2008-04-07" gender="M" nation="BRA" license="384742" swrid="5622287" athleteid="3093" externalid="384742">
              <RESULTS>
                <RESULT eventid="1104" points="400" swimtime="00:00:30.20" resultid="3094" heatid="4299" lane="5" entrytime="00:00:33.15" entrycourse="LCM" />
                <RESULT eventid="1156" points="473" swimtime="00:01:00.13" resultid="3095" heatid="4342" lane="6" entrytime="00:01:02.27" entrycourse="LCM" />
                <RESULT eventid="1188" points="212" swimtime="00:00:43.50" resultid="3096" heatid="4362" lane="1" />
                <RESULT eventid="1236" points="442" swimtime="00:00:27.43" resultid="3097" heatid="4416" lane="1" entrytime="00:00:28.45" entrycourse="LCM" />
                <RESULT eventid="1274" points="312" swimtime="00:02:48.02" resultid="3098" heatid="4444" lane="1" entrytime="00:02:57.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Krik" birthdate="2010-11-24" gender="F" nation="BRA" license="406702" swrid="5717277" athleteid="3114" externalid="406702">
              <RESULTS>
                <RESULT eventid="1148" points="174" swimtime="00:01:32.53" resultid="3115" heatid="4320" lane="6" entrytime="00:01:38.60" entrycourse="LCM" />
                <RESULT eventid="1212" points="125" swimtime="00:02:08.02" resultid="3116" heatid="4379" lane="8" entrytime="00:02:05.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaylaine" lastname="Sofia Vargas Bueno" birthdate="2006-11-28" gender="F" nation="BRA" license="384739" swrid="5622307" athleteid="3086" externalid="384739">
              <RESULTS>
                <RESULT eventid="1080" points="239" swimtime="00:03:41.55" resultid="3087" heatid="4278" lane="4" entrytime="00:03:45.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="231" swimtime="00:00:43.76" resultid="3088" heatid="4470" lane="6" />
                <RESULT eventid="1266" points="232" swimtime="00:03:25.07" resultid="3089" heatid="4435" lane="3" entrytime="00:03:33.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Guarise" birthdate="2008-11-28" gender="M" nation="BRA" license="408881" athleteid="3119" externalid="408881">
              <RESULTS>
                <RESULT eventid="1188" points="268" swimtime="00:00:40.23" resultid="3120" heatid="4361" lane="3" />
                <RESULT eventid="1236" points="339" swimtime="00:00:29.97" resultid="3121" heatid="4408" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Pavin" birthdate="2008-07-17" gender="F" nation="BRA" license="406703" swrid="5717287" athleteid="3117" externalid="406703">
              <RESULTS>
                <RESULT eventid="1228" points="269" swimtime="00:00:36.55" resultid="3118" heatid="4397" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Glir" birthdate="2010-07-01" gender="M" nation="BRA" license="406701" swrid="5717266" athleteid="3110" externalid="406701">
              <RESULTS>
                <RESULT eventid="1156" points="250" swimtime="00:01:14.37" resultid="3111" heatid="4333" lane="5" />
                <RESULT eventid="1188" points="173" swimtime="00:00:46.51" resultid="3112" heatid="4363" lane="2" />
                <RESULT eventid="1236" points="241" swimtime="00:00:33.57" resultid="3113" heatid="4410" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="36" nation="BRA" region="PR" clubid="2228" swrid="93753" name="Associação Atlética Comercial" shortname="Comercial Cascavel">
          <ATHLETES>
            <ATHLETE firstname="Flavia" lastname="De Metz" birthdate="2011-01-07" gender="F" nation="BRA" license="390846" swrid="5596887" athleteid="2397" externalid="390846">
              <RESULTS>
                <RESULT eventid="1064" status="DSQ" swimtime="00:02:56.97" resultid="2398" heatid="4268" lane="2" entrytime="00:03:07.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="349" swimtime="00:11:27.99" resultid="2399" heatid="4426" lane="0" entrytime="00:11:57.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.69" />
                    <SPLIT distance="200" swimtime="00:02:40.76" />
                    <SPLIT distance="300" swimtime="00:04:08.57" />
                    <SPLIT distance="400" swimtime="00:05:36.99" />
                    <SPLIT distance="500" swimtime="00:07:05.48" />
                    <SPLIT distance="600" swimtime="00:08:34.30" />
                    <SPLIT distance="700" swimtime="00:10:03.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="399" swimtime="00:02:33.22" resultid="2400" heatid="4453" lane="8" entrytime="00:02:39.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="319" swimtime="00:01:23.83" resultid="2401" heatid="4520" lane="6" entrytime="00:01:25.61" entrycourse="LCM" />
                <RESULT eventid="1350" points="360" swimtime="00:05:30.59" resultid="2402" heatid="4508" lane="6" entrytime="00:05:31.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.09" />
                    <SPLIT distance="200" swimtime="00:02:38.10" />
                    <SPLIT distance="300" swimtime="00:04:05.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Do Prado Martins" birthdate="2008-10-17" gender="F" nation="BRA" license="369419" swrid="5596893" athleteid="2313" externalid="369419">
              <RESULTS>
                <RESULT eventid="1080" points="416" swimtime="00:03:04.20" resultid="2314" heatid="4281" lane="8" entrytime="00:03:04.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="310" swimtime="00:02:59.83" resultid="2315" heatid="4350" lane="3" entrytime="00:02:45.29" entrycourse="LCM" />
                <RESULT eventid="1132" points="417" swimtime="00:05:55.86" resultid="2316" heatid="4315" lane="3" entrytime="00:05:44.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.89" />
                    <SPLIT distance="200" swimtime="00:02:53.11" />
                    <SPLIT distance="300" swimtime="00:04:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" status="DSQ" swimtime="00:02:41.33" resultid="2317" heatid="4439" lane="6" entrytime="00:02:37.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="452" swimtime="00:01:12.29" resultid="2318" heatid="4497" lane="2" entrytime="00:01:10.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Bertelli Weirich" birthdate="2011-03-18" gender="F" nation="BRA" license="369534" swrid="5588552" athleteid="2325" externalid="369534">
              <RESULTS>
                <RESULT eventid="1064" points="333" swimtime="00:02:57.65" resultid="2326" heatid="4267" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="388" swimtime="00:21:00.96" resultid="2327" heatid="4308" lane="5" entrytime="00:22:41.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.30" />
                    <SPLIT distance="200" swimtime="00:02:36.73" />
                    <SPLIT distance="300" swimtime="00:03:59.39" />
                    <SPLIT distance="400" swimtime="00:05:22.72" />
                    <SPLIT distance="500" swimtime="00:06:47.21" />
                    <SPLIT distance="600" swimtime="00:08:12.14" />
                    <SPLIT distance="700" swimtime="00:09:37.78" />
                    <SPLIT distance="800" swimtime="00:11:03.03" />
                    <SPLIT distance="900" swimtime="00:12:28.36" />
                    <SPLIT distance="1000" swimtime="00:13:54.28" />
                    <SPLIT distance="1100" swimtime="00:15:20.03" />
                    <SPLIT distance="1200" swimtime="00:16:47.24" />
                    <SPLIT distance="1300" swimtime="00:18:14.03" />
                    <SPLIT distance="1400" swimtime="00:19:39.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="385" swimtime="00:06:05.23" resultid="2328" heatid="4314" lane="4" entrytime="00:06:42.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.97" />
                    <SPLIT distance="200" swimtime="00:03:05.01" />
                    <SPLIT distance="300" swimtime="00:04:46.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" points="429" swimtime="00:02:47.11" resultid="2329" heatid="4438" lane="2" entrytime="00:02:52.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="329" swimtime="00:01:20.32" resultid="2330" heatid="4495" lane="4" entrytime="00:01:22.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Luisa Lottermann" birthdate="2011-08-26" gender="F" nation="BRA" license="382238" swrid="5596909" athleteid="2367" externalid="382238">
              <RESULTS>
                <RESULT eventid="1080" points="367" swimtime="00:03:11.97" resultid="2368" heatid="4279" lane="2" entrytime="00:03:23.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="307" swimtime="00:06:33.88" resultid="2369" heatid="4314" lane="3" entrytime="00:06:42.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.05" />
                    <SPLIT distance="200" swimtime="00:03:27.69" />
                    <SPLIT distance="300" swimtime="00:05:08.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="331" swimtime="00:01:32.62" resultid="2370" heatid="4380" lane="4" entrytime="00:01:35.40" entrycourse="LCM" />
                <RESULT eventid="1266" points="277" swimtime="00:03:13.31" resultid="2371" heatid="4435" lane="4" entrytime="00:03:23.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="181" swimtime="00:01:38.02" resultid="2372" heatid="4495" lane="1" entrytime="00:01:40.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luann" lastname="Miguel Mazur" birthdate="2007-01-10" gender="M" nation="BRA" license="365682" swrid="5596915" athleteid="2295" externalid="365682">
              <RESULTS>
                <RESULT eventid="1088" points="482" swimtime="00:02:39.97" resultid="2296" heatid="4288" lane="7" entrytime="00:02:43.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="436" swimtime="00:00:34.21" resultid="2297" heatid="4367" lane="7" entrytime="00:00:35.23" entrycourse="LCM" />
                <RESULT eventid="1140" points="488" swimtime="00:05:07.83" resultid="2298" heatid="4318" lane="7" entrytime="00:05:08.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.66" />
                    <SPLIT distance="200" swimtime="00:02:31.11" />
                    <SPLIT distance="300" swimtime="00:03:56.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="435" swimtime="00:01:15.06" resultid="2299" heatid="4393" lane="7" entrytime="00:01:15.41" entrycourse="LCM" />
                <RESULT eventid="1274" points="476" swimtime="00:02:25.97" resultid="2300" heatid="4447" lane="6" entrytime="00:02:25.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Tolentino Smarczewski" birthdate="2008-09-01" gender="M" nation="BRA" license="378818" swrid="5596941" athleteid="2355" externalid="378818">
              <RESULTS>
                <RESULT eventid="1088" points="426" swimtime="00:02:46.76" resultid="2356" heatid="4283" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="451" swimtime="00:09:49.47" resultid="2357" heatid="4312" lane="3" entrytime="00:09:48.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.35" />
                    <SPLIT distance="200" swimtime="00:02:22.39" />
                    <SPLIT distance="300" swimtime="00:03:38.25" />
                    <SPLIT distance="400" swimtime="00:04:54.87" />
                    <SPLIT distance="500" swimtime="00:06:10.05" />
                    <SPLIT distance="600" swimtime="00:07:25.00" />
                    <SPLIT distance="700" swimtime="00:08:38.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="458" swimtime="00:18:49.92" resultid="2358" heatid="4432" lane="7" entrytime="00:19:05.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.32" />
                    <SPLIT distance="200" swimtime="00:02:23.65" />
                    <SPLIT distance="300" swimtime="00:03:39.17" />
                    <SPLIT distance="400" swimtime="00:04:55.31" />
                    <SPLIT distance="500" swimtime="00:06:12.03" />
                    <SPLIT distance="600" swimtime="00:07:28.60" />
                    <SPLIT distance="700" swimtime="00:08:45.41" />
                    <SPLIT distance="800" swimtime="00:10:01.71" />
                    <SPLIT distance="900" swimtime="00:11:18.02" />
                    <SPLIT distance="1000" swimtime="00:12:34.69" />
                    <SPLIT distance="1100" swimtime="00:13:50.54" />
                    <SPLIT distance="1200" swimtime="00:15:07.42" />
                    <SPLIT distance="1300" swimtime="00:16:23.58" />
                    <SPLIT distance="1400" swimtime="00:17:37.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="468" swimtime="00:02:11.36" resultid="2359" heatid="4467" lane="1" entrytime="00:02:11.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="450" swimtime="00:04:47.12" resultid="2360" heatid="4515" lane="6" entrytime="00:04:41.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.57" />
                    <SPLIT distance="200" swimtime="00:02:18.35" />
                    <SPLIT distance="300" swimtime="00:03:33.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Kupicki" birthdate="2004-03-02" gender="F" nation="BRA" license="311897" swrid="5624094" athleteid="2235" externalid="311897">
              <RESULTS>
                <RESULT eventid="1096" points="386" swimtime="00:00:33.53" resultid="2236" heatid="4293" lane="4" entrytime="00:00:33.74" entrycourse="LCM" />
                <RESULT eventid="1148" points="383" swimtime="00:01:11.20" resultid="2237" heatid="4327" lane="1" entrytime="00:01:08.18" entrycourse="LCM" />
                <RESULT eventid="1180" points="345" swimtime="00:00:41.55" resultid="2238" heatid="4358" lane="2" entrytime="00:00:40.28" entrycourse="LCM" />
                <RESULT eventid="1228" points="374" swimtime="00:00:32.75" resultid="2239" heatid="4396" lane="4" />
                <RESULT eventid="1282" points="345" swimtime="00:02:40.88" resultid="2240" heatid="4450" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Danilo" lastname="Rodrigues" birthdate="2011-05-23" gender="M" nation="BRA" license="370763" swrid="5596934" athleteid="2337" externalid="370763">
              <RESULTS>
                <RESULT eventid="1088" points="317" swimtime="00:03:03.86" resultid="2338" heatid="4284" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="334" swimtime="00:10:51.28" resultid="2339" heatid="4310" lane="8" entrytime="00:11:24.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.50" />
                    <SPLIT distance="200" swimtime="00:02:37.85" />
                    <SPLIT distance="300" swimtime="00:04:01.08" />
                    <SPLIT distance="400" swimtime="00:05:24.92" />
                    <SPLIT distance="500" swimtime="00:06:49.26" />
                    <SPLIT distance="600" swimtime="00:08:11.56" />
                    <SPLIT distance="700" swimtime="00:09:34.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="298" swimtime="00:02:45.10" resultid="2340" heatid="4352" lane="5" entrytime="00:02:53.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="326" swimtime="00:02:28.13" resultid="2341" heatid="4458" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="294" swimtime="00:01:14.30" resultid="2342" heatid="4501" lane="2" entrytime="00:01:14.59" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Luiza Bezerra Sedlacek" birthdate="2008-04-18" gender="F" nation="BRA" license="344607" swrid="4496478" athleteid="2265" externalid="344607">
              <RESULTS>
                <RESULT eventid="1064" points="409" swimtime="00:02:45.86" resultid="2266" heatid="4270" lane="4" entrytime="00:02:44.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="524" swimtime="00:01:04.11" resultid="2267" heatid="4330" lane="1" entrytime="00:01:03.25" entrycourse="LCM" />
                <RESULT eventid="1228" points="507" swimtime="00:00:29.59" resultid="2268" heatid="4404" lane="5" entrytime="00:00:29.53" entrycourse="LCM" />
                <RESULT eventid="1282" points="459" swimtime="00:02:26.23" resultid="2269" heatid="4456" lane="3" entrytime="00:02:18.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" points="471" swimtime="00:02:42.07" resultid="2270" heatid="4439" lane="3" entrytime="00:02:36.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Pedro Signor" birthdate="2005-12-20" gender="M" nation="BRA" license="375814" swrid="5596925" athleteid="2349" externalid="375814">
              <RESULTS>
                <RESULT eventid="1104" points="522" swimtime="00:00:27.65" resultid="2350" heatid="4302" lane="3" entrytime="00:00:28.54" entrycourse="LCM" />
                <RESULT eventid="1140" status="DSQ" swimtime="00:05:51.13" resultid="2351" heatid="4317" lane="2" entrytime="00:05:34.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.97" />
                    <SPLIT distance="200" swimtime="00:02:50.54" />
                    <SPLIT distance="300" swimtime="00:04:36.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="419" swimtime="00:00:27.93" resultid="2352" heatid="4406" lane="7" />
                <RESULT eventid="1306" points="400" swimtime="00:00:31.95" resultid="2353" heatid="4481" lane="4" entrytime="00:00:30.21" entrycourse="LCM" />
                <RESULT eventid="1374" points="345" swimtime="00:01:13.54" resultid="2354" heatid="4531" lane="7" entrytime="00:01:08.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Breno" lastname="Zanella Janke" birthdate="2011-04-26" gender="M" nation="BRA" license="365697" swrid="5588970" athleteid="2319" externalid="365697">
              <RESULTS>
                <RESULT eventid="1088" points="353" swimtime="00:02:57.49" resultid="2320" heatid="4286" lane="8" entrytime="00:03:02.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="378" swimtime="00:05:35.23" resultid="2321" heatid="4316" lane="4" entrytime="00:06:23.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.23" />
                    <SPLIT distance="200" swimtime="00:02:42.41" />
                    <SPLIT distance="300" swimtime="00:04:19.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="336" swimtime="00:01:21.81" resultid="2322" heatid="4390" lane="5" entrytime="00:01:23.39" entrycourse="LCM" />
                <RESULT eventid="1274" points="390" swimtime="00:02:35.91" resultid="2323" heatid="4445" lane="3" entrytime="00:02:39.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="421" swimtime="00:04:53.51" resultid="2324" heatid="4514" lane="5" entrytime="00:04:56.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.64" />
                    <SPLIT distance="200" swimtime="00:02:26.01" />
                    <SPLIT distance="300" swimtime="00:03:42.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raul" lastname="Bonamigo" birthdate="2010-12-01" gender="M" nation="BRA" license="344397" swrid="5588559" athleteid="2379" externalid="344397">
              <RESULTS>
                <RESULT eventid="1072" points="355" swimtime="00:02:37.98" resultid="2380" heatid="4275" lane="7" entrytime="00:02:33.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="2381" heatid="4311" lane="4" entrytime="00:10:16.40" entrycourse="LCM" />
                <RESULT eventid="1258" status="WDR" swimtime="00:00:00.00" resultid="2382" heatid="4432" lane="2" entrytime="00:19:01.75" entrycourse="LCM" />
                <RESULT eventid="1274" status="DNS" swimtime="00:00:00.00" resultid="2383" heatid="4446" lane="7" entrytime="00:02:36.21" entrycourse="LCM" />
                <RESULT eventid="1374" points="334" swimtime="00:01:14.30" resultid="2384" heatid="4529" lane="4" entrytime="00:01:12.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Sehn Uren" birthdate="2009-10-15" gender="F" nation="BRA" license="357159" swrid="5596937" athleteid="2277" externalid="357159">
              <RESULTS>
                <RESULT eventid="1064" points="361" swimtime="00:02:52.93" resultid="2278" heatid="4269" lane="8" entrytime="00:03:01.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="363" swimtime="00:06:12.60" resultid="2279" heatid="4315" lane="1" entrytime="00:06:42.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.76" />
                    <SPLIT distance="200" swimtime="00:03:07.85" />
                    <SPLIT distance="300" swimtime="00:04:48.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="374" swimtime="00:01:28.98" resultid="2280" heatid="4377" lane="3" />
                <RESULT eventid="1266" points="408" swimtime="00:02:49.99" resultid="2281" heatid="4437" lane="6" entrytime="00:03:00.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="352" swimtime="00:01:21.19" resultid="2282" heatid="4520" lane="3" entrytime="00:01:25.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Mariotti De Castro" birthdate="2008-06-27" gender="M" nation="BRA" license="329200" swrid="5596912" athleteid="2247" externalid="329200">
              <RESULTS>
                <RESULT eventid="1124" points="627" swimtime="00:08:48.11" resultid="2248" heatid="4313" lane="4" entrytime="00:08:50.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.41" />
                    <SPLIT distance="200" swimtime="00:02:08.89" />
                    <SPLIT distance="300" swimtime="00:03:14.51" />
                    <SPLIT distance="400" swimtime="00:04:21.84" />
                    <SPLIT distance="500" swimtime="00:05:26.82" />
                    <SPLIT distance="600" swimtime="00:06:35.24" />
                    <SPLIT distance="700" swimtime="00:07:41.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="588" swimtime="00:02:11.67" resultid="2249" heatid="4354" lane="3" entrytime="00:02:12.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="600" swimtime="00:04:47.42" resultid="2250" heatid="4318" lane="4" entrytime="00:04:42.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.09" />
                    <SPLIT distance="200" swimtime="00:02:18.77" />
                    <SPLIT distance="300" swimtime="00:03:44.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1274" points="600" swimtime="00:02:15.14" resultid="2251" heatid="4448" lane="7" entrytime="00:02:17.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="646" swimtime="00:04:14.57" resultid="2252" heatid="4516" lane="6" entrytime="00:04:14.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.53" />
                    <SPLIT distance="200" swimtime="00:02:05.91" />
                    <SPLIT distance="300" swimtime="00:03:09.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Dillenburg Benetti" birthdate="2011-03-10" gender="M" nation="BRA" license="368119" swrid="5588656" athleteid="2307" externalid="368119">
              <RESULTS>
                <RESULT eventid="1072" points="349" swimtime="00:02:38.86" resultid="2308" heatid="4274" lane="7" entrytime="00:02:45.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="325" swimtime="00:05:52.58" resultid="2309" heatid="4316" lane="3" entrytime="00:06:23.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.86" />
                    <SPLIT distance="200" swimtime="00:02:51.71" />
                    <SPLIT distance="300" swimtime="00:04:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="270" swimtime="00:01:27.96" resultid="2310" heatid="4386" lane="6" />
                <RESULT eventid="1274" points="336" swimtime="00:02:43.88" resultid="2311" heatid="4444" lane="4" entrytime="00:02:49.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="335" swimtime="00:01:14.28" resultid="2312" heatid="4528" lane="6" entrytime="00:01:17.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Vitoria Gugel" birthdate="2011-12-08" gender="F" nation="BRA" license="365490" swrid="5588960" athleteid="2409" externalid="365490">
              <RESULTS>
                <RESULT eventid="1096" points="283" swimtime="00:00:37.21" resultid="2410" heatid="4292" lane="6" entrytime="00:00:37.98" entrycourse="LCM" />
                <RESULT eventid="1164" points="241" swimtime="00:03:15.56" resultid="2411" heatid="4349" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="334" swimtime="00:06:22.86" resultid="2412" heatid="4315" lane="8" entrytime="00:06:42.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.09" />
                    <SPLIT distance="200" swimtime="00:03:12.00" />
                    <SPLIT distance="300" swimtime="00:04:56.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" points="347" swimtime="00:02:59.39" resultid="2413" heatid="4437" lane="3" entrytime="00:03:00.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="256" swimtime="00:01:27.31" resultid="2414" heatid="4495" lane="3" entrytime="00:01:29.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Claudio" lastname="Rohnelt" birthdate="2010-03-08" gender="M" nation="BRA" license="357954" swrid="5596935" athleteid="2289" externalid="357954">
              <RESULTS>
                <RESULT eventid="1124" points="325" swimtime="00:10:57.07" resultid="2290" heatid="4310" lane="5" entrytime="00:11:08.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.41" />
                    <SPLIT distance="200" swimtime="00:02:34.32" />
                    <SPLIT distance="300" swimtime="00:03:57.59" />
                    <SPLIT distance="400" swimtime="00:05:21.72" />
                    <SPLIT distance="500" swimtime="00:06:45.61" />
                    <SPLIT distance="600" swimtime="00:08:10.03" />
                    <SPLIT distance="700" swimtime="00:09:33.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="268" swimtime="00:02:51.14" resultid="2291" heatid="4352" lane="2" entrytime="00:02:58.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="341" swimtime="00:20:46.26" resultid="2292" heatid="4431" lane="2" entrytime="00:21:09.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.08" />
                    <SPLIT distance="200" swimtime="00:02:38.81" />
                    <SPLIT distance="300" swimtime="00:04:02.29" />
                    <SPLIT distance="400" swimtime="00:05:26.25" />
                    <SPLIT distance="500" swimtime="00:06:50.35" />
                    <SPLIT distance="600" swimtime="00:08:14.70" />
                    <SPLIT distance="700" swimtime="00:09:38.80" />
                    <SPLIT distance="800" swimtime="00:11:03.03" />
                    <SPLIT distance="900" swimtime="00:12:27.47" />
                    <SPLIT distance="1000" swimtime="00:13:51.87" />
                    <SPLIT distance="1100" swimtime="00:15:16.24" />
                    <SPLIT distance="1200" swimtime="00:16:39.70" />
                    <SPLIT distance="1300" swimtime="00:18:03.31" />
                    <SPLIT distance="1400" swimtime="00:19:25.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="336" swimtime="00:02:26.67" resultid="2293" heatid="4458" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="216" swimtime="00:01:22.41" resultid="2294" heatid="4500" lane="7" entrytime="00:01:18.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Zital" birthdate="1991-05-03" gender="M" nation="BRA" license="093924" athleteid="2421" externalid="093924">
              <RESULTS>
                <RESULT eventid="1072" points="452" swimtime="00:02:25.79" resultid="2422" heatid="4272" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1306" points="500" swimtime="00:00:29.66" resultid="2423" heatid="4477" lane="2" />
                <RESULT eventid="1374" points="453" swimtime="00:01:07.16" resultid="2424" heatid="4525" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emanuel" lastname="Ranieri" birthdate="2011-01-24" gender="M" nation="BRA" license="390838" swrid="5596930" athleteid="2391" externalid="390838">
              <RESULTS>
                <RESULT eventid="1072" points="295" swimtime="00:02:48.02" resultid="2392" heatid="4273" lane="3" entrytime="00:03:00.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="306" swimtime="00:05:59.65" resultid="2393" heatid="4316" lane="2" entrytime="00:06:23.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.85" />
                    <SPLIT distance="200" swimtime="00:02:58.10" />
                    <SPLIT distance="300" swimtime="00:04:41.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="312" swimtime="00:00:30.80" resultid="2394" heatid="4412" lane="5" entrytime="00:00:31.46" entrycourse="LCM" />
                <RESULT eventid="1274" points="323" swimtime="00:02:46.14" resultid="2395" heatid="4441" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1374" points="267" swimtime="00:01:20.04" resultid="2396" heatid="4527" lane="3" entrytime="00:01:22.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hendrik" lastname="Alteiro Groenwold" birthdate="2011-03-23" gender="M" nation="BRA" license="365756" swrid="5588520" athleteid="2301" externalid="365756">
              <RESULTS>
                <RESULT eventid="1072" points="373" swimtime="00:02:35.38" resultid="2302" heatid="4272" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="391" swimtime="00:00:30.44" resultid="2303" heatid="4300" lane="2" entrytime="00:00:31.52" entrycourse="LCM" />
                <RESULT eventid="1172" points="369" swimtime="00:02:33.78" resultid="2304" heatid="4353" lane="8" entrytime="00:02:42.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="396" swimtime="00:02:18.86" resultid="2305" heatid="4464" lane="3" entrytime="00:02:21.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="383" swimtime="00:01:08.04" resultid="2306" heatid="4502" lane="8" entrytime="00:01:11.33" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Stein Duarte" birthdate="2010-10-03" gender="F" nation="BRA" license="351635" swrid="5588923" athleteid="2271" externalid="351635">
              <RESULTS>
                <RESULT eventid="1064" points="459" swimtime="00:02:39.62" resultid="2272" heatid="4271" lane="8" entrytime="00:02:43.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="449" swimtime="00:05:47.17" resultid="2273" heatid="4315" lane="2" entrytime="00:05:51.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.68" />
                    <SPLIT distance="200" swimtime="00:02:48.02" />
                    <SPLIT distance="300" swimtime="00:04:28.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" points="443" swimtime="00:02:45.43" resultid="2274" heatid="4439" lane="8" entrytime="00:02:47.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="319" swimtime="00:01:21.14" resultid="2275" heatid="4493" lane="4" />
                <RESULT eventid="1366" points="473" swimtime="00:01:13.58" resultid="2276" heatid="4523" lane="4" entrytime="00:01:15.53" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Colaco Da Conceicao" birthdate="2011-05-25" gender="F" nation="BRA" license="369535" swrid="5588601" athleteid="2331" externalid="369535">
              <RESULTS>
                <RESULT eventid="1116" points="358" swimtime="00:21:36.30" resultid="2332" heatid="4308" lane="4" entrytime="00:22:41.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.57" />
                    <SPLIT distance="200" swimtime="00:02:37.46" />
                    <SPLIT distance="300" swimtime="00:04:01.26" />
                    <SPLIT distance="400" swimtime="00:05:29.08" />
                    <SPLIT distance="500" swimtime="00:06:59.17" />
                    <SPLIT distance="600" swimtime="00:08:26.42" />
                    <SPLIT distance="700" swimtime="00:09:55.52" />
                    <SPLIT distance="800" swimtime="00:11:23.98" />
                    <SPLIT distance="900" swimtime="00:12:52.19" />
                    <SPLIT distance="1000" swimtime="00:14:21.73" />
                    <SPLIT distance="1100" swimtime="00:15:50.61" />
                    <SPLIT distance="1200" swimtime="00:17:19.45" />
                    <SPLIT distance="1300" swimtime="00:18:45.82" />
                    <SPLIT distance="1400" swimtime="00:20:12.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="278" swimtime="00:03:06.44" resultid="2333" heatid="4350" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:21.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="381" swimtime="00:11:08.61" resultid="2334" heatid="4426" lane="8" entrytime="00:11:57.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.56" />
                    <SPLIT distance="200" swimtime="00:02:38.36" />
                    <SPLIT distance="300" swimtime="00:04:03.23" />
                    <SPLIT distance="400" swimtime="00:05:29.45" />
                    <SPLIT distance="500" swimtime="00:06:55.94" />
                    <SPLIT distance="600" swimtime="00:08:20.62" />
                    <SPLIT distance="700" swimtime="00:09:46.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="416" swimtime="00:02:31.13" resultid="2335" heatid="4450" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="423" swimtime="00:05:13.56" resultid="2336" heatid="4507" lane="5" entrytime="00:05:45.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.06" />
                    <SPLIT distance="200" swimtime="00:02:35.08" />
                    <SPLIT distance="300" swimtime="00:03:56.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Paiz Ribeiro" birthdate="2006-02-17" gender="M" nation="BRA" license="297583" swrid="5596921" athleteid="2229" externalid="297583">
              <RESULTS>
                <RESULT eventid="1088" points="440" swimtime="00:02:44.90" resultid="2230" heatid="4287" lane="4" entrytime="00:02:45.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="494" swimtime="00:02:19.52" resultid="2231" heatid="4354" lane="1" entrytime="00:02:18.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="364" swimtime="00:01:19.65" resultid="2232" heatid="4386" lane="3" />
                <RESULT eventid="1274" points="478" swimtime="00:02:25.79" resultid="2233" heatid="4442" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="498" swimtime="00:01:02.38" resultid="2234" heatid="4504" lane="7" entrytime="00:01:02.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Rinaldini" birthdate="2009-04-09" gender="M" nation="BRA" license="348289" swrid="5596932" athleteid="2259" externalid="348289">
              <RESULTS>
                <RESULT eventid="1124" points="554" swimtime="00:09:10.47" resultid="2260" heatid="4313" lane="1" entrytime="00:09:27.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.62" />
                    <SPLIT distance="200" swimtime="00:02:12.46" />
                    <SPLIT distance="300" swimtime="00:03:22.06" />
                    <SPLIT distance="400" swimtime="00:04:31.71" />
                    <SPLIT distance="500" swimtime="00:05:42.07" />
                    <SPLIT distance="600" swimtime="00:06:52.46" />
                    <SPLIT distance="700" swimtime="00:08:02.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="522" swimtime="00:02:16.98" resultid="2261" heatid="4354" lane="7" entrytime="00:02:18.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="549" swimtime="00:17:43.11" resultid="2262" heatid="4432" lane="8" entrytime="00:19:12.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.36" />
                    <SPLIT distance="200" swimtime="00:02:18.32" />
                    <SPLIT distance="300" swimtime="00:03:30.81" />
                    <SPLIT distance="400" swimtime="00:04:42.72" />
                    <SPLIT distance="500" swimtime="00:05:54.47" />
                    <SPLIT distance="600" swimtime="00:07:05.96" />
                    <SPLIT distance="700" swimtime="00:08:16.95" />
                    <SPLIT distance="800" swimtime="00:09:27.80" />
                    <SPLIT distance="900" swimtime="00:10:38.18" />
                    <SPLIT distance="1000" swimtime="00:11:48.43" />
                    <SPLIT distance="1100" swimtime="00:12:59.70" />
                    <SPLIT distance="1200" swimtime="00:14:11.41" />
                    <SPLIT distance="1300" swimtime="00:15:23.19" />
                    <SPLIT distance="1400" swimtime="00:16:34.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1274" status="DSQ" swimtime="00:02:27.68" resultid="2263" heatid="4447" lane="1" entrytime="00:02:28.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="543" swimtime="00:04:29.61" resultid="2264" heatid="4516" lane="1" entrytime="00:04:31.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.41" />
                    <SPLIT distance="200" swimtime="00:02:11.62" />
                    <SPLIT distance="300" swimtime="00:03:21.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Gamero Prado" birthdate="2007-05-16" gender="F" nation="BRA" license="305973" swrid="5596903" athleteid="2241" externalid="305973">
              <RESULTS>
                <RESULT eventid="1116" points="392" swimtime="00:20:56.94" resultid="2242" heatid="4309" lane="2" entrytime="00:20:42.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.79" />
                    <SPLIT distance="200" swimtime="00:02:38.33" />
                    <SPLIT distance="300" swimtime="00:04:02.76" />
                    <SPLIT distance="400" swimtime="00:05:27.41" />
                    <SPLIT distance="500" swimtime="00:06:51.53" />
                    <SPLIT distance="600" swimtime="00:08:16.22" />
                    <SPLIT distance="700" swimtime="00:09:41.21" />
                    <SPLIT distance="800" swimtime="00:11:05.62" />
                    <SPLIT distance="900" swimtime="00:12:29.35" />
                    <SPLIT distance="1000" swimtime="00:13:54.45" />
                    <SPLIT distance="1100" swimtime="00:15:19.08" />
                    <SPLIT distance="1200" swimtime="00:16:43.47" />
                    <SPLIT distance="1300" swimtime="00:18:09.23" />
                    <SPLIT distance="1400" swimtime="00:19:33.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="351" swimtime="00:02:52.56" resultid="2243" heatid="4350" lane="2" entrytime="00:02:49.53" entrycourse="LCM" />
                <RESULT eventid="1132" points="387" swimtime="00:06:04.77" resultid="2244" heatid="4314" lane="5" entrytime="00:06:42.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.84" />
                    <SPLIT distance="200" swimtime="00:02:53.95" />
                    <SPLIT distance="300" swimtime="00:04:46.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="465" swimtime="00:10:25.38" resultid="2245" heatid="4427" lane="6" entrytime="00:10:41.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.02" />
                    <SPLIT distance="200" swimtime="00:02:31.94" />
                    <SPLIT distance="300" swimtime="00:03:51.62" />
                    <SPLIT distance="400" swimtime="00:05:11.71" />
                    <SPLIT distance="500" swimtime="00:06:30.15" />
                    <SPLIT distance="600" swimtime="00:07:49.34" />
                    <SPLIT distance="700" swimtime="00:09:08.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="393" swimtime="00:01:15.68" resultid="2246" heatid="4496" lane="2" entrytime="00:01:18.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Assakura" birthdate="2010-06-29" gender="F" nation="BRA" license="376473" swrid="5596868" athleteid="2373" externalid="376473">
              <RESULTS>
                <RESULT eventid="1080" points="456" swimtime="00:02:58.64" resultid="2374" heatid="4281" lane="1" entrytime="00:03:04.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="377" swimtime="00:00:40.34" resultid="2375" heatid="4357" lane="4" entrytime="00:00:41.78" entrycourse="LCM" />
                <RESULT eventid="1212" points="399" swimtime="00:01:27.08" resultid="2376" heatid="4382" lane="8" entrytime="00:01:29.72" entrycourse="LCM" />
                <RESULT eventid="1282" points="433" swimtime="00:02:29.15" resultid="2377" heatid="4454" lane="8" entrytime="00:02:34.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="400" swimtime="00:05:19.33" resultid="2378" heatid="4507" lane="6" entrytime="00:05:46.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.63" />
                    <SPLIT distance="200" swimtime="00:02:35.60" />
                    <SPLIT distance="300" swimtime="00:03:57.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jordana" lastname="Rinaldini" birthdate="2004-09-13" gender="F" nation="BRA" license="342426" swrid="5596933" athleteid="2253" externalid="342426">
              <RESULTS>
                <RESULT eventid="1080" points="349" swimtime="00:03:15.35" resultid="2254" heatid="4281" lane="7" entrytime="00:03:04.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="418" swimtime="00:00:38.99" resultid="2255" heatid="4358" lane="6" entrytime="00:00:39.55" entrycourse="LCM" />
                <RESULT eventid="1212" points="406" swimtime="00:01:26.59" resultid="2256" heatid="4382" lane="4" entrytime="00:01:26.41" entrycourse="LCM" />
                <RESULT eventid="1298" points="400" swimtime="00:00:36.43" resultid="2257" heatid="4473" lane="3" entrytime="00:00:37.94" entrycourse="LCM" />
                <RESULT eventid="1366" points="357" swimtime="00:01:20.74" resultid="2258" heatid="4521" lane="3" entrytime="00:01:22.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Borille Busetti" birthdate="2010-02-17" gender="F" nation="BRA" license="392830" swrid="5622263" athleteid="2415" externalid="392830">
              <RESULTS>
                <RESULT eventid="1064" points="244" swimtime="00:03:16.99" resultid="2416" heatid="4268" lane="8" entrytime="00:03:20.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="380" swimtime="00:01:11.38" resultid="2417" heatid="4324" lane="1" entrytime="00:01:13.20" entrycourse="LCM" />
                <RESULT eventid="1212" points="223" swimtime="00:01:45.75" resultid="2418" heatid="4378" lane="4" />
                <RESULT eventid="1282" points="350" swimtime="00:02:39.99" resultid="2419" heatid="4452" lane="5" entrytime="00:02:42.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="264" swimtime="00:01:29.26" resultid="2420" heatid="4519" lane="8" entrytime="00:01:34.13" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Cordeiro Silva" birthdate="2011-09-04" gender="M" nation="BRA" license="380664" swrid="5596877" athleteid="2361" externalid="380664">
              <RESULTS>
                <RESULT eventid="1088" points="251" swimtime="00:03:18.68" resultid="2362" heatid="4284" lane="4" entrytime="00:03:21.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="254" swimtime="00:00:40.96" resultid="2363" heatid="4365" lane="2" entrytime="00:00:40.75" entrycourse="LCM" />
                <RESULT eventid="1220" points="236" swimtime="00:01:32.04" resultid="2364" heatid="4389" lane="1" entrytime="00:01:32.44" entrycourse="LCM" />
                <RESULT eventid="1290" points="208" swimtime="00:02:51.96" resultid="2365" heatid="4459" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" status="DSQ" swimtime="00:01:29.91" resultid="2366" heatid="4499" lane="2" entrytime="00:01:31.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Balduíno" birthdate="2009-06-24" gender="M" nation="BRA" license="370764" swrid="5596870" athleteid="2343" externalid="370764">
              <RESULTS>
                <RESULT eventid="1088" points="321" swimtime="00:03:03.10" resultid="2344" heatid="4286" lane="7" entrytime="00:02:58.76" entrycourse="LCM" />
                <RESULT eventid="1140" points="392" swimtime="00:05:31.08" resultid="2345" heatid="4317" lane="5" entrytime="00:05:20.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.02" />
                    <SPLIT distance="200" swimtime="00:02:37.77" />
                    <SPLIT distance="300" swimtime="00:04:16.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="290" swimtime="00:01:25.93" resultid="2346" heatid="4386" lane="7" />
                <RESULT eventid="1274" points="405" swimtime="00:02:33.97" resultid="2347" heatid="4446" lane="6" entrytime="00:02:33.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="377" swimtime="00:01:08.42" resultid="2348" heatid="4502" lane="4" entrytime="00:01:05.33" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ramirez Vasconcelos" birthdate="2011-04-06" gender="M" nation="BRA" license="392013" swrid="4863662" athleteid="2403" externalid="392013">
              <RESULTS>
                <RESULT eventid="1088" points="249" swimtime="00:03:19.29" resultid="2404" heatid="4284" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="295" swimtime="00:11:18.86" resultid="2405" heatid="4310" lane="6" entrytime="00:11:24.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.14" />
                    <SPLIT distance="200" swimtime="00:02:42.66" />
                    <SPLIT distance="300" swimtime="00:04:10.74" />
                    <SPLIT distance="400" swimtime="00:05:38.65" />
                    <SPLIT distance="500" swimtime="00:07:06.96" />
                    <SPLIT distance="600" swimtime="00:08:32.46" />
                    <SPLIT distance="700" swimtime="00:09:59.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" status="DSQ" swimtime="00:00:39.19" resultid="2406" heatid="4360" lane="4" />
                <RESULT eventid="1220" points="252" swimtime="00:01:30.05" resultid="2407" heatid="4386" lane="1" />
                <RESULT eventid="1290" points="313" swimtime="00:02:30.11" resultid="2408" heatid="4460" lane="3" entrytime="00:02:45.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Zimmermann" birthdate="2010-01-19" gender="M" nation="BRA" license="357160" swrid="5588977" athleteid="2283" externalid="357160">
              <RESULTS>
                <RESULT eventid="1072" points="461" swimtime="00:02:24.86" resultid="2284" heatid="4276" lane="6" entrytime="00:02:27.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="483" swimtime="00:05:09.01" resultid="2285" heatid="4318" lane="1" entrytime="00:05:12.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.88" />
                    <SPLIT distance="200" swimtime="00:02:29.26" />
                    <SPLIT distance="300" swimtime="00:03:59.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="451" swimtime="00:02:12.96" resultid="2286" heatid="4459" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1274" points="466" swimtime="00:02:27.04" resultid="2287" heatid="4447" lane="8" entrytime="00:02:29.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="343" swimtime="00:01:10.58" resultid="2288" heatid="4498" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Alves Serafini" birthdate="2008-04-15" gender="M" nation="BRA" license="351644" swrid="5596867" athleteid="2385" externalid="351644">
              <RESULTS>
                <RESULT eventid="1104" points="489" swimtime="00:00:28.26" resultid="2386" heatid="4302" lane="6" entrytime="00:00:28.60" entrycourse="LCM" />
                <RESULT eventid="1172" points="516" swimtime="00:02:17.48" resultid="2387" heatid="4353" lane="4" entrytime="00:02:23.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="467" swimtime="00:00:26.95" resultid="2388" heatid="4418" lane="7" entrytime="00:00:27.04" entrycourse="LCM" />
                <RESULT eventid="1290" points="534" swimtime="00:02:05.68" resultid="2389" heatid="4467" lane="6" entrytime="00:02:09.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="512" swimtime="00:01:01.78" resultid="2390" heatid="4503" lane="5" entrytime="00:01:02.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1204" points="408" swimtime="00:09:23.96" resultid="2431" heatid="4373" lane="0">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.00" />
                    <SPLIT distance="200" swimtime="00:02:21.61" />
                    <SPLIT distance="300" swimtime="00:03:29.23" />
                    <SPLIT distance="400" swimtime="00:04:43.16" />
                    <SPLIT distance="500" swimtime="00:05:52.70" />
                    <SPLIT distance="600" swimtime="00:07:11.22" />
                    <SPLIT distance="700" swimtime="00:08:13.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2319" number="1" />
                    <RELAYPOSITION athleteid="2301" number="2" />
                    <RELAYPOSITION athleteid="2379" number="3" />
                    <RELAYPOSITION athleteid="2283" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1206" points="559" swimtime="00:08:28.02" resultid="2432" heatid="4374" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.65" />
                    <SPLIT distance="200" swimtime="00:02:02.39" />
                    <SPLIT distance="300" swimtime="00:03:02.86" />
                    <SPLIT distance="500" swimtime="00:05:10.31" />
                    <SPLIT distance="600" swimtime="00:06:17.51" />
                    <SPLIT distance="700" swimtime="00:07:19.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2247" number="1" />
                    <RELAYPOSITION athleteid="2385" number="2" />
                    <RELAYPOSITION athleteid="2259" number="3" />
                    <RELAYPOSITION athleteid="2355" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1324" points="369" swimtime="00:04:48.04" resultid="2433" heatid="4488" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.27" />
                    <SPLIT distance="200" swimtime="00:02:34.43" />
                    <SPLIT distance="300" swimtime="00:03:42.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2307" number="1" />
                    <RELAYPOSITION athleteid="2319" number="2" />
                    <RELAYPOSITION athleteid="2301" number="3" />
                    <RELAYPOSITION athleteid="2391" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1392" points="390" swimtime="00:04:17.63" resultid="2436" heatid="4539" lane="2">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:02:06.43" />
                    <SPLIT distance="300" swimtime="00:03:10.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2319" number="1" />
                    <RELAYPOSITION athleteid="2301" number="2" />
                    <RELAYPOSITION athleteid="2307" number="3" />
                    <RELAYPOSITION athleteid="2391" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1326" points="340" swimtime="00:04:56.12" resultid="2434" heatid="4489" lane="5" entrytime="00:04:39.35">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.06" />
                    <SPLIT distance="200" swimtime="00:02:33.69" />
                    <SPLIT distance="300" swimtime="00:03:49.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2283" number="1" />
                    <RELAYPOSITION athleteid="2337" number="2" />
                    <RELAYPOSITION athleteid="2289" number="3" />
                    <RELAYPOSITION athleteid="2379" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1394" points="360" swimtime="00:04:24.41" resultid="2437" heatid="4540" lane="1">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:02:08.62" />
                    <SPLIT distance="300" swimtime="00:03:18.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2283" number="1" />
                    <RELAYPOSITION athleteid="2337" number="2" />
                    <RELAYPOSITION athleteid="2289" number="3" />
                    <RELAYPOSITION athleteid="2379" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1330" points="481" swimtime="00:04:23.88" resultid="2435" heatid="4491" lane="5" entrytime="00:04:24.69">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.63" />
                    <SPLIT distance="200" swimtime="00:02:22.86" />
                    <SPLIT distance="300" swimtime="00:03:26.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2247" number="1" />
                    <RELAYPOSITION athleteid="2355" number="2" />
                    <RELAYPOSITION athleteid="2259" number="3" />
                    <RELAYPOSITION athleteid="2385" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1398" points="498" swimtime="00:03:57.40" resultid="2439" heatid="4542" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.73" />
                    <SPLIT distance="200" swimtime="00:01:56.54" />
                    <SPLIT distance="300" swimtime="00:02:56.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2247" number="1" />
                    <RELAYPOSITION athleteid="2385" number="2" />
                    <RELAYPOSITION athleteid="2259" number="3" />
                    <RELAYPOSITION athleteid="2355" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1400" points="447" swimtime="00:04:06.19" resultid="2438" heatid="4543" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.63" />
                    <SPLIT distance="200" swimtime="00:02:05.64" />
                    <SPLIT distance="300" swimtime="00:03:06.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2349" number="1" />
                    <RELAYPOSITION athleteid="2229" number="2" />
                    <RELAYPOSITION athleteid="2295" number="3" />
                    <RELAYPOSITION athleteid="2421" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1196" points="426" swimtime="00:10:07.55" resultid="2426" heatid="4370" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.64" />
                    <SPLIT distance="200" swimtime="00:02:31.55" />
                    <SPLIT distance="300" swimtime="00:03:45.98" />
                    <SPLIT distance="500" swimtime="00:06:19.87" />
                    <SPLIT distance="600" swimtime="00:07:37.88" />
                    <SPLIT distance="700" swimtime="00:08:49.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2397" number="1" />
                    <RELAYPOSITION athleteid="2271" number="2" />
                    <RELAYPOSITION athleteid="2325" number="3" />
                    <RELAYPOSITION athleteid="2373" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1316" points="379" swimtime="00:05:18.24" resultid="2428" heatid="4484" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.71" />
                    <SPLIT distance="200" swimtime="00:02:41.72" />
                    <SPLIT distance="300" swimtime="00:04:08.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2271" number="1" />
                    <RELAYPOSITION athleteid="2373" number="2" />
                    <RELAYPOSITION athleteid="2331" number="3" />
                    <RELAYPOSITION athleteid="2415" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1384" points="399" swimtime="00:04:42.25" resultid="2429" heatid="4535" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.72" />
                    <SPLIT distance="200" swimtime="00:02:22.73" />
                    <SPLIT distance="300" swimtime="00:03:33.43" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2271" number="1" />
                    <RELAYPOSITION athleteid="2373" number="2" />
                    <RELAYPOSITION athleteid="2415" number="3" />
                    <RELAYPOSITION athleteid="2397" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1382" points="348" swimtime="00:04:55.64" resultid="2430" heatid="4534" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.44" />
                    <SPLIT distance="200" swimtime="00:02:29.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2325" number="1" />
                    <RELAYPOSITION athleteid="2367" number="2" />
                    <RELAYPOSITION athleteid="2409" number="3" />
                    <RELAYPOSITION athleteid="2331" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="COMERCIAL CASCAVEL &quot;A&quot;" number="20">
              <RESULTS>
                <RESULT eventid="1314" points="343" swimtime="00:05:28.88" resultid="2427" heatid="4483" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2325" number="1" />
                    <RELAYPOSITION athleteid="2367" number="2" />
                    <RELAYPOSITION athleteid="2409" number="3" />
                    <RELAYPOSITION athleteid="2397" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1112" status="DSQ" swimtime="00:05:00.79" resultid="2440" heatid="4306" lane="6" entrytime="00:05:04.16">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:02:43.80" />
                    <SPLIT distance="300" swimtime="00:03:51.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2325" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2319" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="2301" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="2397" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1114" points="381" swimtime="00:04:59.95" resultid="2441" heatid="4307" lane="5" entrytime="00:04:53.53">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.80" />
                    <SPLIT distance="200" swimtime="00:02:44.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2271" number="1" />
                    <RELAYPOSITION athleteid="2373" number="2" />
                    <RELAYPOSITION athleteid="2283" number="3" />
                    <RELAYPOSITION athleteid="2379" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1248" points="440" swimtime="00:04:45.98" resultid="2442" heatid="4425" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.71" />
                    <SPLIT distance="200" swimtime="00:02:36.14" />
                    <SPLIT distance="300" swimtime="00:03:38.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2253" number="1" />
                    <RELAYPOSITION athleteid="2295" number="2" />
                    <RELAYPOSITION athleteid="2229" number="3" />
                    <RELAYPOSITION athleteid="2241" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1246" points="510" swimtime="00:04:32.26" resultid="2443" heatid="4424" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.29" />
                    <SPLIT distance="200" swimtime="00:02:26.62" />
                    <SPLIT distance="300" swimtime="00:03:28.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2247" number="1" />
                    <RELAYPOSITION athleteid="2313" number="2" />
                    <RELAYPOSITION athleteid="2385" number="3" />
                    <RELAYPOSITION athleteid="2265" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="COMERCIAL CASCAVEL &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1112" points="330" swimtime="00:05:14.58" resultid="2425" heatid="4305" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.42" />
                    <SPLIT distance="200" swimtime="00:02:47.15" />
                    <SPLIT distance="300" swimtime="00:04:00.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2307" number="1" />
                    <RELAYPOSITION athleteid="2367" number="2" />
                    <RELAYPOSITION athleteid="2337" number="3" />
                    <RELAYPOSITION athleteid="2409" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="2864" nation="BRA" region="PR" clubid="1452" swrid="93756" name="Associacao De Pais E Amigos Da Natacao De Ponta Gr" shortname="Apan Ponta Grossa">
          <ATHLETES>
            <ATHLETE firstname="Yoseph" lastname="Rigoni Moraes" birthdate="2006-04-17" gender="M" nation="BRA" license="295182" swrid="5622302" athleteid="1508" externalid="295182">
              <RESULTS>
                <RESULT eventid="1104" points="531" swimtime="00:00:27.50" resultid="1509" heatid="4303" lane="3" entrytime="00:00:27.65" entrycourse="LCM" />
                <RESULT eventid="1188" points="475" swimtime="00:00:33.25" resultid="1510" heatid="4368" lane="6" entrytime="00:00:32.60" entrycourse="LCM" />
                <RESULT eventid="1236" points="513" swimtime="00:00:26.11" resultid="1511" heatid="4420" lane="8" entrytime="00:00:25.97" entrycourse="LCM" />
                <RESULT eventid="1306" points="437" swimtime="00:00:31.03" resultid="1512" heatid="4482" lane="8" entrytime="00:00:30.19" entrycourse="LCM" />
                <RESULT eventid="1374" points="437" swimtime="00:01:07.99" resultid="1513" heatid="4531" lane="3" entrytime="00:01:07.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Dolinski Thomassewski" birthdate="2006-12-15" gender="M" nation="BRA" license="400409" swrid="5653289" athleteid="1543" externalid="400409">
              <RESULTS>
                <RESULT eventid="1156" points="291" swimtime="00:01:10.67" resultid="1544" heatid="4336" lane="3" entrytime="00:01:11.60" entrycourse="LCM" />
                <RESULT eventid="1188" points="274" swimtime="00:00:39.92" resultid="1545" heatid="4365" lane="1" entrytime="00:00:41.42" entrycourse="LCM" />
                <RESULT eventid="1220" points="238" swimtime="00:01:31.67" resultid="1546" heatid="4389" lane="4" entrytime="00:01:30.30" entrycourse="LCM" />
                <RESULT eventid="1236" status="DNS" swimtime="00:00:00.00" resultid="1547" heatid="4409" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Gueiber Montes" birthdate="2009-03-09" gender="M" nation="BRA" license="342154" swrid="5600179" athleteid="1453" externalid="342154">
              <RESULTS>
                <RESULT eventid="1156" points="625" swimtime="00:00:54.80" resultid="1454" heatid="4347" lane="8" entrytime="00:00:55.98" entrycourse="LCM" />
                <RESULT eventid="1236" points="573" swimtime="00:00:25.17" resultid="1455" heatid="4420" lane="1" entrytime="00:00:25.69" entrycourse="LCM" />
                <RESULT eventid="1290" points="556" swimtime="00:02:04.02" resultid="1456" heatid="4468" lane="2" entrytime="00:02:04.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1306" points="536" swimtime="00:00:28.99" resultid="1457" heatid="4482" lane="1" entrytime="00:00:28.83" entrycourse="LCM" />
                <RESULT eventid="1374" points="576" swimtime="00:01:02.00" resultid="1458" heatid="4533" lane="7" entrytime="00:01:01.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Augusto" lastname="Tramontin" birthdate="2011-11-29" gender="M" nation="BRA" license="399691" swrid="5652901" athleteid="1525" externalid="399691">
              <RESULTS>
                <RESULT eventid="1156" points="358" swimtime="00:01:05.94" resultid="1526" heatid="4337" lane="2" entrytime="00:01:10.07" entrycourse="LCM" />
                <RESULT eventid="1188" points="309" swimtime="00:00:38.38" resultid="1527" heatid="4364" lane="2" entrytime="00:00:44.78" entrycourse="LCM" />
                <RESULT eventid="1220" points="264" swimtime="00:01:28.65" resultid="1528" heatid="4389" lane="7" entrytime="00:01:31.92" entrycourse="LCM" />
                <RESULT eventid="1236" points="367" swimtime="00:00:29.18" resultid="1529" heatid="4412" lane="6" entrytime="00:00:31.95" entrycourse="LCM" />
                <RESULT eventid="1306" points="287" swimtime="00:00:35.69" resultid="1530" heatid="4479" lane="8" entrytime="00:00:38.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Brenda" lastname="Gabriele Carvalho" birthdate="2010-04-11" gender="F" nation="BRA" license="399557" swrid="5658060" athleteid="1514" externalid="399557">
              <RESULTS>
                <RESULT eventid="1180" points="219" swimtime="00:00:48.36" resultid="1515" heatid="4355" lane="5" />
                <RESULT eventid="1228" points="208" swimtime="00:00:39.83" resultid="1516" heatid="4398" lane="7" entrytime="00:00:38.78" entrycourse="LCM" />
                <RESULT eventid="1212" points="221" swimtime="00:01:46.06" resultid="1517" heatid="4379" lane="5" entrytime="00:01:49.61" entrycourse="LCM" />
                <RESULT eventid="1298" points="281" swimtime="00:00:40.96" resultid="1518" heatid="4472" lane="7" entrytime="00:00:44.53" entrycourse="LCM" />
                <RESULT eventid="1366" points="258" swimtime="00:01:30.02" resultid="1519" heatid="4518" lane="4" entrytime="00:01:35.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Delinski" birthdate="2009-11-28" gender="F" nation="BRA" license="385190" swrid="5600150" athleteid="1491" externalid="385190">
              <RESULTS>
                <RESULT eventid="1064" points="315" swimtime="00:03:00.95" resultid="1492" heatid="4267" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="314" swimtime="00:00:42.87" resultid="1493" heatid="4357" lane="6" entrytime="00:00:42.30" entrycourse="LCM" />
                <RESULT eventid="1212" points="319" swimtime="00:01:33.82" resultid="1494" heatid="4381" lane="7" entrytime="00:01:33.61" entrycourse="LCM" />
                <RESULT eventid="1298" points="365" swimtime="00:00:37.58" resultid="1495" heatid="4471" lane="7" />
                <RESULT eventid="1366" points="333" swimtime="00:01:22.68" resultid="1496" heatid="4521" lane="8" entrytime="00:01:23.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fegert" birthdate="2009-04-13" gender="M" nation="BRA" license="353813" swrid="5622279" athleteid="1497" externalid="353813">
              <RESULTS>
                <RESULT eventid="1104" points="431" swimtime="00:00:29.48" resultid="1498" heatid="4300" lane="7" entrytime="00:00:31.76" entrycourse="LCM" />
                <RESULT eventid="1156" points="467" swimtime="00:01:00.38" resultid="1499" heatid="4343" lane="7" entrytime="00:01:01.32" entrycourse="LCM" />
                <RESULT eventid="1236" points="445" swimtime="00:00:27.37" resultid="1500" heatid="4407" lane="1" />
                <RESULT eventid="1342" points="367" swimtime="00:01:09.02" resultid="1501" heatid="4502" lane="1" entrytime="00:01:10.21" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Allana" lastname="Lacerda" birthdate="2005-03-15" gender="F" nation="BRA" license="295186" swrid="5600197" athleteid="1469" externalid="295186">
              <RESULTS>
                <RESULT eventid="1080" status="DSQ" swimtime="00:03:03.36" resultid="1470" heatid="4282" lane="8" entrytime="00:02:58.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="422" swimtime="00:00:38.85" resultid="1471" heatid="4358" lane="4" entrytime="00:00:38.77" entrycourse="LCM" />
                <RESULT eventid="1212" points="425" swimtime="00:01:25.23" resultid="1472" heatid="4383" lane="5" entrytime="00:01:22.04" entrycourse="LCM" />
                <RESULT eventid="1266" points="422" swimtime="00:02:48.04" resultid="1473" heatid="4439" lane="7" entrytime="00:02:41.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="297" swimtime="00:01:23.08" resultid="1474" heatid="4496" lane="8" entrytime="00:01:20.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Carraro Borges" birthdate="2009-05-11" gender="M" nation="BRA" license="345590" swrid="5622267" athleteid="1502" externalid="345590">
              <RESULTS>
                <RESULT eventid="1124" points="381" swimtime="00:10:23.33" resultid="1503" heatid="4312" lane="1" entrytime="00:10:01.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.43" />
                    <SPLIT distance="200" swimtime="00:02:26.51" />
                    <SPLIT distance="300" swimtime="00:03:45.70" />
                    <SPLIT distance="400" swimtime="00:05:06.15" />
                    <SPLIT distance="500" swimtime="00:06:27.23" />
                    <SPLIT distance="600" swimtime="00:07:48.09" />
                    <SPLIT distance="700" swimtime="00:09:07.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="445" swimtime="00:01:01.34" resultid="1504" heatid="4342" lane="8" entrytime="00:01:03.46" entrycourse="LCM" />
                <RESULT eventid="1258" points="424" swimtime="00:19:19.25" resultid="1505" heatid="4431" lane="4" entrytime="00:20:07.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.43" />
                    <SPLIT distance="200" swimtime="00:02:26.13" />
                    <SPLIT distance="300" swimtime="00:03:44.69" />
                    <SPLIT distance="400" swimtime="00:05:03.15" />
                    <SPLIT distance="500" swimtime="00:06:21.06" />
                    <SPLIT distance="600" swimtime="00:07:40.74" />
                    <SPLIT distance="700" swimtime="00:08:59.08" />
                    <SPLIT distance="800" swimtime="00:10:17.03" />
                    <SPLIT distance="900" swimtime="00:11:35.46" />
                    <SPLIT distance="1000" swimtime="00:12:53.78" />
                    <SPLIT distance="1100" swimtime="00:14:11.60" />
                    <SPLIT distance="1200" swimtime="00:15:29.42" />
                    <SPLIT distance="1300" swimtime="00:16:47.76" />
                    <SPLIT distance="1400" swimtime="00:18:05.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="410" swimtime="00:00:28.14" resultid="1506" heatid="4415" lane="6" entrytime="00:00:29.31" entrycourse="LCM" />
                <RESULT eventid="1358" points="426" swimtime="00:04:52.44" resultid="1507" heatid="4514" lane="7" entrytime="00:05:02.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.30" />
                    <SPLIT distance="200" swimtime="00:02:21.34" />
                    <SPLIT distance="300" swimtime="00:03:37.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Carolina Babiuki" birthdate="2007-02-06" gender="F" nation="BRA" license="316227" swrid="5600131" athleteid="1485" externalid="316227">
              <RESULTS>
                <RESULT eventid="1064" points="432" swimtime="00:02:42.81" resultid="1486" heatid="4271" lane="7" entrytime="00:02:40.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="545" swimtime="00:01:03.28" resultid="1487" heatid="4329" lane="3" entrytime="00:01:04.18" entrycourse="LCM" />
                <RESULT eventid="1228" points="517" swimtime="00:00:29.41" resultid="1488" heatid="4405" lane="7" entrytime="00:00:29.00" entrycourse="LCM" />
                <RESULT eventid="1298" points="530" swimtime="00:00:33.17" resultid="1489" heatid="4475" lane="3" entrytime="00:00:32.70" entrycourse="LCM" />
                <RESULT eventid="1366" points="452" swimtime="00:01:14.68" resultid="1490" heatid="4524" lane="1" entrytime="00:01:12.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Viechineski Bernardes" birthdate="2011-02-26" gender="M" nation="BRA" license="390879" swrid="5602588" athleteid="1520" externalid="390879">
              <RESULTS>
                <RESULT eventid="1104" points="76" swimtime="00:00:52.43" resultid="1521" heatid="4295" lane="6" />
                <RESULT eventid="1156" points="229" swimtime="00:01:16.55" resultid="1522" heatid="4332" lane="2" />
                <RESULT eventid="1188" points="161" swimtime="00:00:47.69" resultid="1523" heatid="4362" lane="4" />
                <RESULT eventid="1236" points="233" swimtime="00:00:33.98" resultid="1524" heatid="4407" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Chi Kravchychyn" birthdate="2009-09-27" gender="M" nation="BRA" license="344268" swrid="5600134" athleteid="1459" externalid="344268">
              <RESULTS>
                <RESULT eventid="1088" points="520" swimtime="00:02:36.04" resultid="1460" heatid="4289" lane="1" entrytime="00:02:31.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="449" swimtime="00:02:24.07" resultid="1461" heatid="4354" lane="2" entrytime="00:02:16.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="508" swimtime="00:05:03.73" resultid="1462" heatid="4318" lane="3" entrytime="00:04:51.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.44" />
                    <SPLIT distance="200" swimtime="00:02:27.48" />
                    <SPLIT distance="300" swimtime="00:03:54.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1220" points="494" swimtime="00:01:11.92" resultid="1463" heatid="4394" lane="6" entrytime="00:01:09.95" entrycourse="LCM" />
                <RESULT eventid="1274" points="524" swimtime="00:02:21.35" resultid="1464" heatid="4448" lane="1" entrytime="00:02:17.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yohan" lastname="Rigoni Moraes" birthdate="2002-04-03" gender="M" nation="BRA" license="272187" swrid="5600245" athleteid="1465" externalid="272187">
              <RESULTS>
                <RESULT eventid="1088" points="553" swimtime="00:02:32.79" resultid="1466" heatid="4288" lane="5" entrytime="00:02:35.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="738" swimtime="00:00:28.71" resultid="1467" heatid="4369" lane="6" entrytime="00:00:29.15" entrycourse="LCM" />
                <RESULT eventid="1220" points="632" swimtime="00:01:06.25" resultid="1468" heatid="4395" lane="8" entrytime="00:01:07.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Sabedotti" birthdate="2011-04-20" gender="F" nation="BRA" license="390877" swrid="5602580" athleteid="1537" externalid="390877">
              <RESULTS>
                <RESULT eventid="1064" points="339" swimtime="00:02:56.53" resultid="1538" heatid="4269" lane="2" entrytime="00:02:57.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="428" swimtime="00:01:08.59" resultid="1539" heatid="4326" lane="5" entrytime="00:01:09.20" entrycourse="LCM" />
                <RESULT eventid="1228" points="440" swimtime="00:00:31.03" resultid="1540" heatid="4401" lane="8" entrytime="00:00:32.56" entrycourse="LCM" />
                <RESULT eventid="1298" points="455" swimtime="00:00:34.92" resultid="1541" heatid="4474" lane="5" entrytime="00:00:36.58" entrycourse="LCM" />
                <RESULT eventid="1366" status="DNS" swimtime="00:00:00.00" resultid="1542" heatid="4522" lane="1" entrytime="00:01:19.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Franca Berger" birthdate="2010-05-07" gender="F" nation="BRA" license="399692" swrid="5653290" athleteid="1531" externalid="399692">
              <RESULTS>
                <RESULT eventid="1080" points="218" swimtime="00:03:48.42" resultid="1532" heatid="4278" lane="5" entrytime="00:03:55.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="252" swimtime="00:01:21.86" resultid="1533" heatid="4322" lane="7" entrytime="00:01:21.34" entrycourse="LCM" />
                <RESULT eventid="1180" points="225" swimtime="00:00:47.88" resultid="1534" heatid="4356" lane="2" entrytime="00:00:52.07" entrycourse="LCM" />
                <RESULT eventid="1228" points="291" swimtime="00:00:35.62" resultid="1535" heatid="4398" lane="3" entrytime="00:00:37.82" entrycourse="LCM" />
                <RESULT eventid="1212" points="203" swimtime="00:01:49.08" resultid="1536" heatid="4380" lane="1" entrytime="00:01:44.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Campagnoli" birthdate="2009-04-13" gender="F" nation="BRA" license="366915" swrid="5600128" athleteid="1475" externalid="366915">
              <RESULTS>
                <RESULT eventid="1064" points="430" swimtime="00:02:43.14" resultid="1476" heatid="4271" lane="1" entrytime="00:02:42.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="514" swimtime="00:01:04.55" resultid="1477" heatid="4329" lane="7" entrytime="00:01:04.80" entrycourse="LCM" />
                <RESULT eventid="1228" points="478" swimtime="00:00:30.18" resultid="1478" heatid="4404" lane="8" entrytime="00:00:30.26" entrycourse="LCM" />
                <RESULT eventid="1298" points="517" swimtime="00:00:33.45" resultid="1479" heatid="4475" lane="2" entrytime="00:00:34.49" entrycourse="LCM" />
                <RESULT eventid="1366" points="458" swimtime="00:01:14.35" resultid="1480" heatid="4524" lane="8" entrytime="00:01:14.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Reda" birthdate="2007-05-21" gender="F" nation="BRA" license="316228" swrid="5600241" athleteid="1481" externalid="316228">
              <RESULTS>
                <RESULT eventid="1148" status="DSQ" swimtime="00:01:11.69" resultid="1482" heatid="4324" lane="5" entrytime="00:01:11.86" entrycourse="LCM" />
                <RESULT eventid="1228" points="398" swimtime="00:00:32.08" resultid="1483" heatid="4401" lane="6" entrytime="00:00:32.28" entrycourse="LCM" />
                <RESULT eventid="1298" points="362" swimtime="00:00:37.68" resultid="1484" heatid="4474" lane="2" entrytime="00:00:37.29" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/PONTA GROSSA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1328" points="482" swimtime="00:04:23.71" resultid="1548" heatid="4490" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.68" />
                    <SPLIT distance="200" swimtime="00:02:15.64" />
                    <SPLIT distance="300" swimtime="00:03:23.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1453" number="1" />
                    <RELAYPOSITION athleteid="1459" number="2" />
                    <RELAYPOSITION athleteid="1497" number="3" />
                    <RELAYPOSITION athleteid="1502" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1396" points="514" swimtime="00:03:54.97" resultid="1549" heatid="4541" lane="3">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:01:58.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1459" number="1" />
                    <RELAYPOSITION athleteid="1497" number="2" />
                    <RELAYPOSITION athleteid="1502" number="3" />
                    <RELAYPOSITION athleteid="1453" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/PONTA GROSSA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1248" points="470" swimtime="00:04:39.74" resultid="1550" heatid="4425" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.53" />
                    <SPLIT distance="200" swimtime="00:02:24.28" />
                    <SPLIT distance="300" swimtime="00:03:31.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1485" number="1" />
                    <RELAYPOSITION athleteid="1465" number="2" />
                    <RELAYPOSITION athleteid="1508" number="3" />
                    <RELAYPOSITION athleteid="1469" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/PONTA GROSSA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1244" points="421" swimtime="00:04:50.09" resultid="1551" heatid="4423" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.76" />
                    <SPLIT distance="200" swimtime="00:02:37.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1453" number="1" />
                    <RELAYPOSITION athleteid="1491" number="2" />
                    <RELAYPOSITION athleteid="1497" number="3" />
                    <RELAYPOSITION athleteid="1475" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="13068" nation="BRA" region="PR" clubid="3251" swrid="93787" name="Sociedade Morgenau" shortname="Morgenau">
          <ATHLETES>
            <ATHLETE firstname="Jhenyffer" lastname="Stefany Szaida" birthdate="2006-09-16" gender="F" nation="BRA" license="369326" swrid="5600264" athleteid="3312" externalid="369326">
              <RESULTS>
                <RESULT eventid="1096" points="298" swimtime="00:00:36.54" resultid="3313" heatid="4293" lane="8" entrytime="00:00:37.00" entrycourse="LCM" />
                <RESULT eventid="1298" points="298" swimtime="00:00:40.20" resultid="3314" heatid="4470" lane="3" />
                <RESULT eventid="1266" points="266" swimtime="00:03:15.96" resultid="3315" heatid="4436" lane="7" entrytime="00:03:12.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="200" swimtime="00:01:34.85" resultid="3316" heatid="4495" lane="2" entrytime="00:01:30.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Gabriel Sarmento Buski" birthdate="2010-04-05" gender="M" nation="BRA" license="399533" swrid="5717264" athleteid="3279" externalid="399533">
              <RESULTS>
                <RESULT eventid="1188" points="240" swimtime="00:00:41.70" resultid="3280" heatid="4362" lane="8" />
                <RESULT eventid="1220" points="210" swimtime="00:01:35.59" resultid="3281" heatid="4388" lane="5" entrytime="00:01:33.87" entrycourse="LCM" />
                <RESULT eventid="1258" points="309" swimtime="00:21:27.10" resultid="3282" heatid="4430" lane="6" entrytime="00:21:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.48" />
                    <SPLIT distance="200" swimtime="00:02:38.71" />
                    <SPLIT distance="300" swimtime="00:04:05.50" />
                    <SPLIT distance="400" swimtime="00:05:31.66" />
                    <SPLIT distance="500" swimtime="00:06:59.04" />
                    <SPLIT distance="600" swimtime="00:08:24.89" />
                    <SPLIT distance="700" swimtime="00:09:51.17" />
                    <SPLIT distance="800" swimtime="00:11:18.90" />
                    <SPLIT distance="900" swimtime="00:12:47.16" />
                    <SPLIT distance="1000" swimtime="00:14:15.01" />
                    <SPLIT distance="1100" swimtime="00:15:42.06" />
                    <SPLIT distance="1200" swimtime="00:17:09.86" />
                    <SPLIT distance="1300" swimtime="00:18:37.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="267" swimtime="00:02:38.27" resultid="3283" heatid="4461" lane="5" entrytime="00:02:36.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Fernanda Pinto" birthdate="2004-09-17" gender="F" nation="BRA" license="391144" swrid="5600157" athleteid="3378" externalid="391144">
              <RESULTS>
                <RESULT eventid="1096" points="242" swimtime="00:00:39.18" resultid="3379" heatid="4292" lane="2" entrytime="00:00:41.73" entrycourse="LCM" />
                <RESULT eventid="1148" points="377" swimtime="00:01:11.53" resultid="3380" heatid="4323" lane="6" entrytime="00:01:13.88" entrycourse="LCM" />
                <RESULT eventid="1298" points="286" swimtime="00:00:40.76" resultid="3381" heatid="4472" lane="8" entrytime="00:00:46.16" entrycourse="LCM" />
                <RESULT eventid="1334" points="199" swimtime="00:01:34.97" resultid="3382" heatid="4495" lane="7" entrytime="00:01:35.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stella" lastname="Magalhaes Birnbaum" birthdate="2009-05-14" gender="F" nation="BRA" license="399684" swrid="5653298" athleteid="3416" externalid="399684">
              <RESULTS>
                <RESULT eventid="1096" points="237" swimtime="00:00:39.45" resultid="3417" heatid="4291" lane="2" />
                <RESULT eventid="1148" points="381" swimtime="00:01:11.28" resultid="3418" heatid="4323" lane="7" entrytime="00:01:14.23" entrycourse="LCM" />
                <RESULT eventid="1228" points="367" swimtime="00:00:32.97" resultid="3419" heatid="4400" lane="6" entrytime="00:00:32.89" entrycourse="LCM" />
                <RESULT eventid="1298" points="329" swimtime="00:00:38.87" resultid="3420" heatid="4472" lane="3" entrytime="00:00:42.27" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monike" lastname="Lemos Carvalho" birthdate="2008-03-28" gender="F" nation="BRA" license="307796" swrid="5600199" athleteid="3352" externalid="307796">
              <RESULTS>
                <RESULT eventid="1148" points="479" swimtime="00:01:06.06" resultid="3353" heatid="4327" lane="2" entrytime="00:01:08.11" entrycourse="LCM" />
                <RESULT eventid="1250" points="384" swimtime="00:11:06.45" resultid="3354" heatid="4427" lane="8" entrytime="00:11:05.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.69" />
                    <SPLIT distance="200" swimtime="00:02:42.09" />
                    <SPLIT distance="300" swimtime="00:04:07.65" />
                    <SPLIT distance="400" swimtime="00:05:33.24" />
                    <SPLIT distance="500" swimtime="00:06:56.32" />
                    <SPLIT distance="600" swimtime="00:08:21.25" />
                    <SPLIT distance="700" swimtime="00:09:45.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="468" swimtime="00:02:25.33" resultid="3355" heatid="4456" lane="8" entrytime="00:02:25.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="356" swimtime="00:01:20.82" resultid="3356" heatid="4523" lane="2" entrytime="00:01:17.55" entrycourse="LCM" />
                <RESULT eventid="1350" points="401" swimtime="00:05:19.07" resultid="3357" heatid="4509" lane="8" entrytime="00:05:23.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.77" />
                    <SPLIT distance="200" swimtime="00:02:35.16" />
                    <SPLIT distance="300" swimtime="00:03:58.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Mingorance Martins" birthdate="2007-10-13" gender="M" nation="BRA" license="393920" swrid="5622295" athleteid="3404" externalid="393920">
              <RESULTS>
                <RESULT eventid="1072" points="347" swimtime="00:02:39.18" resultid="3405" heatid="4274" lane="2" entrytime="00:02:44.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="546" swimtime="00:00:57.30" resultid="3406" heatid="4346" lane="2" entrytime="00:00:57.58" entrycourse="LCM" />
                <RESULT eventid="1236" points="524" swimtime="00:00:25.92" resultid="3407" heatid="4419" lane="2" entrytime="00:00:26.50" entrycourse="LCM" />
                <RESULT eventid="1290" points="493" swimtime="00:02:09.07" resultid="3408" heatid="4466" lane="3" entrytime="00:02:13.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="418" swimtime="00:04:54.11" resultid="3409" heatid="4514" lane="1" entrytime="00:05:04.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.85" />
                    <SPLIT distance="200" swimtime="00:02:17.87" />
                    <SPLIT distance="300" swimtime="00:03:35.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Portella Da Silva" birthdate="2010-07-19" gender="M" nation="BRA" license="399534" swrid="5717288" athleteid="3284" externalid="399534">
              <RESULTS>
                <RESULT eventid="1188" points="217" swimtime="00:00:43.13" resultid="3285" heatid="4362" lane="7" />
                <RESULT eventid="1306" points="171" swimtime="00:00:42.39" resultid="3286" heatid="4477" lane="6" />
                <RESULT eventid="1274" points="152" swimtime="00:03:33.30" resultid="3287" heatid="4442" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Matos Oliveira" birthdate="2007-10-26" gender="M" nation="BRA" license="391136" swrid="5600215" athleteid="3358" externalid="391136">
              <RESULTS>
                <RESULT eventid="1124" points="328" swimtime="00:10:55.31" resultid="3359" heatid="4311" lane="8" entrytime="00:10:59.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.83" />
                    <SPLIT distance="200" swimtime="00:02:35.98" />
                    <SPLIT distance="300" swimtime="00:03:58.96" />
                    <SPLIT distance="500" swimtime="00:06:46.87" />
                    <SPLIT distance="600" swimtime="00:08:10.73" />
                    <SPLIT distance="700" swimtime="00:09:34.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="290" swimtime="00:00:33.63" resultid="3360" heatid="4298" lane="2" entrytime="00:00:38.92" entrycourse="LCM" />
                <RESULT eventid="1188" points="233" swimtime="00:00:42.15" resultid="3361" heatid="4364" lane="5" entrytime="00:00:42.71" entrycourse="LCM" />
                <RESULT eventid="1258" points="341" swimtime="00:20:45.87" resultid="3362" heatid="4431" lane="7" entrytime="00:21:37.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="200" swimtime="00:02:37.53" />
                    <SPLIT distance="300" swimtime="00:04:01.24" />
                    <SPLIT distance="400" swimtime="00:05:25.12" />
                    <SPLIT distance="500" swimtime="00:06:49.54" />
                    <SPLIT distance="600" swimtime="00:08:13.46" />
                    <SPLIT distance="700" swimtime="00:09:37.91" />
                    <SPLIT distance="800" swimtime="00:11:02.35" />
                    <SPLIT distance="900" swimtime="00:12:26.86" />
                    <SPLIT distance="1000" swimtime="00:13:50.35" />
                    <SPLIT distance="1100" swimtime="00:15:14.78" />
                    <SPLIT distance="1200" swimtime="00:16:39.23" />
                    <SPLIT distance="1300" swimtime="00:18:03.47" />
                    <SPLIT distance="1400" swimtime="00:19:26.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="351" swimtime="00:05:11.95" resultid="3363" heatid="4513" lane="7" entrytime="00:05:22.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.55" />
                    <SPLIT distance="200" swimtime="00:02:32.23" />
                    <SPLIT distance="300" swimtime="00:03:53.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauan" lastname="Araujo" birthdate="2009-12-17" gender="M" nation="BRA" license="385119" swrid="5653286" athleteid="3340" externalid="385119">
              <RESULTS>
                <RESULT eventid="1156" points="382" swimtime="00:01:04.56" resultid="3341" heatid="4341" lane="2" entrytime="00:01:04.73" entrycourse="LCM" />
                <RESULT eventid="1188" points="262" swimtime="00:00:40.53" resultid="3342" heatid="4364" lane="7" entrytime="00:00:45.93" entrycourse="LCM" />
                <RESULT eventid="1220" points="242" swimtime="00:01:31.17" resultid="3343" heatid="4389" lane="3" entrytime="00:01:30.76" entrycourse="LCM" />
                <RESULT eventid="1236" points="353" swimtime="00:00:29.56" resultid="3344" heatid="4413" lane="8" entrytime="00:00:31.41" entrycourse="LCM" />
                <RESULT eventid="1290" points="349" swimtime="00:02:24.87" resultid="3345" heatid="4463" lane="4" entrytime="00:02:25.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Luiz Fischer" birthdate="2009-06-07" gender="M" nation="BRA" license="400273" swrid="5653296" athleteid="3423" externalid="400273">
              <RESULTS>
                <RESULT eventid="1104" points="351" swimtime="00:00:31.55" resultid="3424" heatid="4299" lane="7" entrytime="00:00:34.58" entrycourse="LCM" />
                <RESULT eventid="1220" points="231" swimtime="00:01:32.69" resultid="3425" heatid="4387" lane="4" entrytime="00:01:39.46" entrycourse="LCM" />
                <RESULT eventid="1274" points="213" swimtime="00:03:10.78" resultid="3426" heatid="4442" lane="3" entrytime="00:03:18.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" points="234" swimtime="00:01:20.15" resultid="3427" heatid="4499" lane="3" entrytime="00:01:25.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Vitoria De Lima" birthdate="2011-06-10" gender="F" nation="BRA" license="400090" swrid="5652904" athleteid="3421" externalid="400090">
              <RESULTS>
                <RESULT eventid="1228" status="DSQ" swimtime="00:00:42.89" resultid="3422" heatid="4397" lane="4" entrytime="00:00:42.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thiago" lastname="Kozera Chiarato" birthdate="2008-01-22" gender="M" nation="BRA" license="406728" swrid="5717276" athleteid="3457" externalid="406728">
              <RESULTS>
                <RESULT eventid="1104" points="315" swimtime="00:00:32.70" resultid="3458" heatid="4296" lane="5" />
                <RESULT eventid="1172" points="222" swimtime="00:03:02.05" resultid="3459" heatid="4351" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="366" swimtime="00:00:29.23" resultid="3460" heatid="4407" lane="8" />
                <RESULT eventid="1290" points="319" swimtime="00:02:29.19" resultid="3461" heatid="4462" lane="6" entrytime="00:02:32.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" status="DSQ" swimtime="00:01:15.02" resultid="3462" heatid="4500" lane="8" entrytime="00:01:19.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Bora" birthdate="2005-01-06" gender="F" nation="BRA" license="358252" swrid="5600153" athleteid="3306" externalid="358252">
              <RESULTS>
                <RESULT eventid="1064" points="323" swimtime="00:02:59.29" resultid="3307" heatid="4269" lane="1" entrytime="00:02:59.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="215" swimtime="00:01:46.97" resultid="3308" heatid="4378" lane="7" />
                <RESULT eventid="1266" points="313" swimtime="00:03:05.68" resultid="3309" heatid="4437" lane="8" entrytime="00:03:01.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="298" swimtime="00:01:25.76" resultid="3310" heatid="4520" lane="4" entrytime="00:01:24.43" entrycourse="LCM" />
                <RESULT eventid="1350" points="339" swimtime="00:05:37.53" resultid="3311" heatid="4508" lane="8" entrytime="00:05:38.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.99" />
                    <SPLIT distance="200" swimtime="00:02:44.86" />
                    <SPLIT distance="300" swimtime="00:04:11.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Geovana" lastname="Dos Santos" birthdate="2011-01-20" gender="F" nation="BRA" license="367254" swrid="5602533" athleteid="3300" externalid="367254">
              <RESULTS>
                <RESULT eventid="1148" points="315" swimtime="00:01:15.96" resultid="3301" heatid="4322" lane="6" entrytime="00:01:18.67" entrycourse="LCM" />
                <RESULT eventid="1228" points="317" swimtime="00:00:34.62" resultid="3302" heatid="4399" lane="1" entrytime="00:00:35.62" entrycourse="LCM" />
                <RESULT eventid="1282" points="319" swimtime="00:02:45.06" resultid="3303" heatid="4452" lane="1" entrytime="00:02:49.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="287" swimtime="00:00:40.68" resultid="3304" heatid="4473" lane="7" entrytime="00:00:40.67" entrycourse="LCM" />
                <RESULT eventid="1366" points="267" swimtime="00:01:28.94" resultid="3305" heatid="4519" lane="5" entrytime="00:01:29.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Lima" birthdate="2006-12-03" gender="M" nation="BRA" license="366749" swrid="5600201" athleteid="3329" externalid="366749">
              <RESULTS>
                <RESULT eventid="1104" points="542" swimtime="00:00:27.31" resultid="3330" heatid="4303" lane="8" entrytime="00:00:28.12" entrycourse="LCM" />
                <RESULT eventid="1156" points="594" swimtime="00:00:55.72" resultid="3331" heatid="4347" lane="1" entrytime="00:00:55.97" entrycourse="LCM" />
                <RESULT eventid="1236" points="566" swimtime="00:00:25.27" resultid="3332" heatid="4420" lane="4" entrytime="00:00:25.44" entrycourse="LCM" />
                <RESULT eventid="1342" points="474" swimtime="00:01:03.42" resultid="3333" heatid="4503" lane="4" entrytime="00:01:02.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Luiza Rimbano De Jesus" birthdate="2008-09-02" gender="F" nation="BRA" license="366819" swrid="5653297" athleteid="3410" externalid="366819">
              <RESULTS>
                <RESULT eventid="1148" points="555" swimtime="00:01:02.89" resultid="3411" heatid="4328" lane="4" entrytime="00:01:05.51" entrycourse="LCM" />
                <RESULT eventid="1180" points="443" swimtime="00:00:38.24" resultid="3412" heatid="4358" lane="8" entrytime="00:00:41.52" entrycourse="LCM" />
                <RESULT eventid="1228" points="546" swimtime="00:00:28.87" resultid="3413" heatid="4404" lane="4" entrytime="00:00:29.40" entrycourse="LCM" />
                <RESULT eventid="1282" points="481" swimtime="00:02:24.01" resultid="3414" heatid="4455" lane="4" entrytime="00:02:25.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="341" swimtime="00:01:19.36" resultid="3415" heatid="4494" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauren" lastname="Dziura" birthdate="2010-01-11" gender="F" nation="BRA" license="369416" swrid="5588668" athleteid="3323" externalid="369416">
              <RESULTS>
                <RESULT eventid="1064" points="306" swimtime="00:03:02.56" resultid="3324" heatid="4268" lane="5" entrytime="00:03:03.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="331" swimtime="00:11:40.39" resultid="3325" heatid="4427" lane="0" entrytime="00:11:12.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.89" />
                    <SPLIT distance="200" swimtime="00:02:46.21" />
                    <SPLIT distance="300" swimtime="00:04:15.46" />
                    <SPLIT distance="400" swimtime="00:05:45.26" />
                    <SPLIT distance="500" swimtime="00:07:14.81" />
                    <SPLIT distance="600" swimtime="00:08:43.56" />
                    <SPLIT distance="700" swimtime="00:10:14.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="363" swimtime="00:02:38.18" resultid="3326" heatid="4453" lane="6" entrytime="00:02:34.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" points="344" swimtime="00:02:59.97" resultid="3327" heatid="4436" lane="2" entrytime="00:03:12.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="283" swimtime="00:01:27.25" resultid="3328" heatid="4520" lane="5" entrytime="00:01:24.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Kozera Chiarato" birthdate="2010-05-28" gender="M" nation="BRA" license="406722" swrid="5717275" athleteid="3439" externalid="406722">
              <RESULTS>
                <RESULT eventid="1104" points="257" swimtime="00:00:35.02" resultid="3440" heatid="4295" lane="4" />
                <RESULT eventid="1188" points="207" swimtime="00:00:43.85" resultid="3441" heatid="4363" lane="7" />
                <RESULT eventid="1220" points="191" swimtime="00:01:38.73" resultid="3442" heatid="4388" lane="8" entrytime="00:01:39.27" entrycourse="LCM" />
                <RESULT eventid="1236" points="251" swimtime="00:00:33.12" resultid="3443" heatid="4406" lane="2" />
                <RESULT eventid="1342" points="221" swimtime="00:01:21.70" resultid="3444" heatid="4499" lane="5" entrytime="00:01:25.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karine" lastname="Correa" birthdate="2002-08-01" gender="F" nation="BRA" license="385191" swrid="5600141" athleteid="3346" externalid="385191">
              <RESULTS>
                <RESULT eventid="1116" points="288" swimtime="00:23:12.84" resultid="3347" heatid="4308" lane="2" entrytime="00:22:41.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.52" />
                    <SPLIT distance="200" swimtime="00:02:50.73" />
                    <SPLIT distance="300" swimtime="00:04:23.43" />
                    <SPLIT distance="400" swimtime="00:05:57.18" />
                    <SPLIT distance="500" swimtime="00:07:31.37" />
                    <SPLIT distance="600" swimtime="00:09:05.72" />
                    <SPLIT distance="700" swimtime="00:10:40.14" />
                    <SPLIT distance="800" swimtime="00:12:14.67" />
                    <SPLIT distance="900" swimtime="00:13:51.33" />
                    <SPLIT distance="1000" swimtime="00:15:26.64" />
                    <SPLIT distance="1100" swimtime="00:17:01.50" />
                    <SPLIT distance="1200" swimtime="00:18:36.59" />
                    <SPLIT distance="1300" swimtime="00:20:11.44" />
                    <SPLIT distance="1400" swimtime="00:21:45.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="369" swimtime="00:01:12.05" resultid="3348" heatid="4324" lane="3" entrytime="00:01:12.16" entrycourse="LCM" />
                <RESULT eventid="1250" points="274" swimtime="00:12:25.87" resultid="3349" heatid="4426" lane="7" entrytime="00:11:50.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.41" />
                    <SPLIT distance="200" swimtime="00:03:04.79" />
                    <SPLIT distance="300" swimtime="00:04:43.01" />
                    <SPLIT distance="400" swimtime="00:06:21.33" />
                    <SPLIT distance="500" swimtime="00:07:59.86" />
                    <SPLIT distance="600" swimtime="00:09:37.95" />
                    <SPLIT distance="700" swimtime="00:11:14.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1266" points="272" swimtime="00:03:14.44" resultid="3350" heatid="4436" lane="1" entrytime="00:03:12.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1350" points="302" swimtime="00:05:50.46" resultid="3351" heatid="4508" lane="7" entrytime="00:05:36.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.41" />
                    <SPLIT distance="200" swimtime="00:02:47.80" />
                    <SPLIT distance="300" swimtime="00:04:20.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Madalena De Lima" birthdate="2006-05-04" gender="M" nation="BRA" license="307786" swrid="5600206" athleteid="3257" externalid="307786">
              <RESULTS>
                <RESULT eventid="1124" points="392" swimtime="00:10:17.74" resultid="3258" heatid="4312" lane="7" entrytime="00:09:57.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.23" />
                    <SPLIT distance="200" swimtime="00:02:20.79" />
                    <SPLIT distance="300" swimtime="00:03:36.47" />
                    <SPLIT distance="400" swimtime="00:04:53.39" />
                    <SPLIT distance="500" swimtime="00:06:12.35" />
                    <SPLIT distance="600" swimtime="00:07:34.42" />
                    <SPLIT distance="700" swimtime="00:08:57.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="468" swimtime="00:02:11.29" resultid="3259" heatid="4466" lane="4" entrytime="00:02:12.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="455" swimtime="00:04:45.98" resultid="3260" heatid="4515" lane="1" entrytime="00:04:45.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.72" />
                    <SPLIT distance="200" swimtime="00:02:17.11" />
                    <SPLIT distance="300" swimtime="00:03:31.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Herick" lastname="Dos Santos" birthdate="2009-06-11" gender="M" nation="BRA" license="406724" swrid="5717258" athleteid="3448" externalid="406724">
              <RESULTS>
                <RESULT eventid="1104" points="90" swimtime="00:00:49.52" resultid="3449" heatid="4297" lane="1" />
                <RESULT eventid="1156" points="182" swimtime="00:01:22.65" resultid="3450" heatid="4332" lane="4" />
                <RESULT eventid="1188" status="DSQ" swimtime="00:01:10.86" resultid="3451" heatid="4361" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kedny" lastname="Correa" birthdate="2004-11-05" gender="M" nation="BRA" license="383858" swrid="5600142" athleteid="3334" externalid="383858">
              <RESULTS>
                <RESULT eventid="1124" points="436" swimtime="00:09:55.97" resultid="3335" heatid="4312" lane="2" entrytime="00:09:54.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.18" />
                    <SPLIT distance="200" swimtime="00:02:18.21" />
                    <SPLIT distance="300" swimtime="00:03:32.12" />
                    <SPLIT distance="400" swimtime="00:04:48.02" />
                    <SPLIT distance="500" swimtime="00:06:04.96" />
                    <SPLIT distance="600" swimtime="00:07:21.77" />
                    <SPLIT distance="700" swimtime="00:08:39.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="290" swimtime="00:02:46.52" resultid="3336" heatid="4353" lane="1" entrytime="00:02:39.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="429" swimtime="00:19:14.79" resultid="3337" heatid="4432" lane="1" entrytime="00:19:10.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.60" />
                    <SPLIT distance="200" swimtime="00:02:17.78" />
                    <SPLIT distance="300" swimtime="00:03:33.34" />
                    <SPLIT distance="400" swimtime="00:04:50.42" />
                    <SPLIT distance="500" swimtime="00:06:08.50" />
                    <SPLIT distance="600" swimtime="00:07:26.92" />
                    <SPLIT distance="700" swimtime="00:08:44.74" />
                    <SPLIT distance="800" swimtime="00:10:03.43" />
                    <SPLIT distance="900" swimtime="00:11:21.68" />
                    <SPLIT distance="1000" swimtime="00:12:40.59" />
                    <SPLIT distance="1100" swimtime="00:13:59.19" />
                    <SPLIT distance="1200" swimtime="00:15:19.29" />
                    <SPLIT distance="1300" swimtime="00:16:38.82" />
                    <SPLIT distance="1400" swimtime="00:17:57.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1274" points="419" swimtime="00:02:32.26" resultid="3338" heatid="4441" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="421" swimtime="00:04:53.43" resultid="3339" heatid="4515" lane="2" entrytime="00:04:44.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.50" />
                    <SPLIT distance="200" swimtime="00:02:17.75" />
                    <SPLIT distance="300" swimtime="00:03:35.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Marcos Pinto" birthdate="2006-01-26" gender="M" nation="BRA" license="391143" swrid="5600209" athleteid="3373" externalid="391143">
              <RESULTS>
                <RESULT eventid="1156" points="317" swimtime="00:01:08.68" resultid="3374" heatid="4337" lane="6" entrytime="00:01:09.95" entrycourse="LCM" />
                <RESULT eventid="1188" points="248" swimtime="00:00:41.29" resultid="3375" heatid="4364" lane="3" entrytime="00:00:42.92" entrycourse="LCM" />
                <RESULT eventid="1290" points="273" swimtime="00:02:37.18" resultid="3376" heatid="4462" lane="8" entrytime="00:02:36.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1274" status="DSQ" swimtime="00:03:03.50" resultid="3377" heatid="4442" lane="2" entrytime="00:03:22.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mayara" lastname="Fieber" birthdate="2008-08-20" gender="F" nation="BRA" license="391147" swrid="5600161" athleteid="3395" externalid="391147">
              <RESULTS>
                <RESULT eventid="1064" points="278" swimtime="00:03:08.66" resultid="3396" heatid="4268" lane="6" entrytime="00:03:06.45" entrycourse="LCM" />
                <RESULT eventid="1228" points="374" swimtime="00:00:32.75" resultid="3397" heatid="4399" lane="6" entrytime="00:00:34.29" entrycourse="LCM" />
                <RESULT eventid="1298" points="316" swimtime="00:00:39.41" resultid="3398" heatid="4473" lane="8" entrytime="00:00:41.27" entrycourse="LCM" />
                <RESULT eventid="1266" points="307" swimtime="00:03:06.88" resultid="3399" heatid="4436" lane="8" entrytime="00:03:23.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1366" points="278" swimtime="00:01:27.81" resultid="3400" heatid="4520" lane="1" entrytime="00:01:28.13" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Capoia Soares" birthdate="2011-11-07" gender="M" nation="BRA" license="393257" swrid="5616440" athleteid="3401" externalid="393257">
              <RESULTS>
                <RESULT eventid="1104" points="64" swimtime="00:00:55.50" resultid="3402" heatid="4295" lane="1" />
                <RESULT eventid="1156" points="108" swimtime="00:01:38.27" resultid="3403" heatid="4334" lane="1" entrytime="00:01:38.47" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Henrique Opuchkevich" birthdate="2011-02-22" gender="M" nation="BRA" license="406720" swrid="5717273" athleteid="3434" externalid="406720">
              <RESULTS>
                <RESULT eventid="1156" points="230" swimtime="00:01:16.45" resultid="3435" heatid="4335" lane="3" entrytime="00:01:16.67" entrycourse="LCM" />
                <RESULT eventid="1188" points="206" swimtime="00:00:43.89" resultid="3436" heatid="4362" lane="5" />
                <RESULT eventid="1220" points="205" swimtime="00:01:36.33" resultid="3437" heatid="4388" lane="1" entrytime="00:01:38.52" entrycourse="LCM" />
                <RESULT eventid="1274" points="198" swimtime="00:03:15.34" resultid="3438" heatid="4441" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Rodrigues Galvao" birthdate="2007-04-19" gender="M" nation="BRA" license="376586" swrid="5600247" athleteid="3267" externalid="376586">
              <RESULTS>
                <RESULT eventid="1104" points="522" swimtime="00:00:27.65" resultid="3268" heatid="4302" lane="5" entrytime="00:00:28.31" entrycourse="LCM" />
                <RESULT eventid="1156" points="514" swimtime="00:00:58.47" resultid="3269" heatid="4346" lane="8" entrytime="00:00:58.39" entrycourse="LCM" />
                <RESULT eventid="1172" points="355" swimtime="00:02:35.79" resultid="3270" heatid="4353" lane="2" entrytime="00:02:36.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="510" swimtime="00:00:26.17" resultid="3271" heatid="4419" lane="5" entrytime="00:00:26.22" entrycourse="LCM" />
                <RESULT eventid="1342" points="430" swimtime="00:01:05.51" resultid="3272" heatid="4503" lane="3" entrytime="00:01:03.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Andreis Ramos" birthdate="2007-03-26" gender="M" nation="BRA" license="406719" swrid="5717243" athleteid="3428" externalid="406719">
              <RESULTS>
                <RESULT eventid="1104" points="321" swimtime="00:00:32.50" resultid="3429" heatid="4297" lane="7" />
                <RESULT eventid="1156" points="345" swimtime="00:01:06.75" resultid="3430" heatid="4340" lane="5" entrytime="00:01:05.69" entrycourse="LCM" />
                <RESULT eventid="1236" points="343" swimtime="00:00:29.87" resultid="3431" heatid="4409" lane="1" />
                <RESULT eventid="1306" points="262" swimtime="00:00:36.79" resultid="3432" heatid="4476" lane="4" />
                <RESULT eventid="1342" points="232" swimtime="00:01:20.38" resultid="3433" heatid="4499" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benito" lastname="Alves Sant&apos;Ana" birthdate="2009-06-01" gender="M" nation="BRA" license="376585" swrid="5351951" athleteid="3273" externalid="376585">
              <RESULTS>
                <RESULT eventid="1124" points="499" swimtime="00:09:29.92" resultid="3274" heatid="4313" lane="2" entrytime="00:09:22.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.76" />
                    <SPLIT distance="200" swimtime="00:02:13.56" />
                    <SPLIT distance="300" swimtime="00:03:24.77" />
                    <SPLIT distance="400" swimtime="00:04:35.46" />
                    <SPLIT distance="500" swimtime="00:05:49.87" />
                    <SPLIT distance="600" swimtime="00:07:04.58" />
                    <SPLIT distance="700" swimtime="00:08:19.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="451" swimtime="00:05:16.11" resultid="3275" heatid="4317" lane="4" entrytime="00:05:19.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.14" />
                    <SPLIT distance="200" swimtime="00:02:36.20" />
                    <SPLIT distance="300" swimtime="00:04:10.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1258" points="526" swimtime="00:17:58.38" resultid="3276" heatid="4430" lane="5" entrytime="00:21:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.71" />
                    <SPLIT distance="200" swimtime="00:02:16.76" />
                    <SPLIT distance="300" swimtime="00:03:29.45" />
                    <SPLIT distance="400" swimtime="00:04:41.65" />
                    <SPLIT distance="500" swimtime="00:05:54.41" />
                    <SPLIT distance="600" swimtime="00:07:07.15" />
                    <SPLIT distance="700" swimtime="00:08:19.68" />
                    <SPLIT distance="800" swimtime="00:09:30.45" />
                    <SPLIT distance="900" swimtime="00:10:42.97" />
                    <SPLIT distance="1000" swimtime="00:11:55.17" />
                    <SPLIT distance="1100" swimtime="00:13:08.52" />
                    <SPLIT distance="1200" swimtime="00:14:21.67" />
                    <SPLIT distance="1300" swimtime="00:15:35.24" />
                    <SPLIT distance="1400" swimtime="00:16:48.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1274" points="411" swimtime="00:02:33.26" resultid="3277" heatid="4446" lane="5" entrytime="00:02:31.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="491" swimtime="00:04:38.95" resultid="3278" heatid="4515" lane="7" entrytime="00:04:44.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.32" />
                    <SPLIT distance="200" swimtime="00:02:17.11" />
                    <SPLIT distance="300" swimtime="00:03:28.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Barros Zagonel" birthdate="2006-06-01" gender="M" nation="BRA" license="347856" swrid="5622261" athleteid="3252" externalid="347856">
              <RESULTS>
                <RESULT eventid="1088" points="264" swimtime="00:03:15.49" resultid="3253" heatid="4285" lane="8" entrytime="00:03:18.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="393" swimtime="00:00:35.42" resultid="3254" heatid="4367" lane="1" entrytime="00:00:35.44" entrycourse="LCM" />
                <RESULT eventid="1220" points="291" swimtime="00:01:25.76" resultid="3255" heatid="4390" lane="2" entrytime="00:01:26.03" entrycourse="LCM" />
                <RESULT eventid="1274" points="301" swimtime="00:02:50.05" resultid="3256" heatid="4444" lane="2" entrytime="00:02:53.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Isabel Santos" birthdate="2005-12-20" gender="F" nation="BRA" license="391141" swrid="5600191" athleteid="3370" externalid="391141">
              <RESULTS>
                <RESULT eventid="1282" points="296" swimtime="00:02:49.28" resultid="3371" heatid="4451" lane="2" entrytime="00:02:55.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="180" swimtime="00:01:38.18" resultid="3372" heatid="4495" lane="8" entrytime="00:01:40.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Yoshie Kimura" birthdate="2010-07-08" gender="F" nation="BRA" license="391142" swrid="5600277" athleteid="3288" externalid="391142">
              <RESULTS>
                <RESULT eventid="1080" points="424" swimtime="00:03:03.05" resultid="3289" heatid="4280" lane="4" entrytime="00:03:08.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="456" swimtime="00:00:37.87" resultid="3290" heatid="4358" lane="3" entrytime="00:00:39.48" entrycourse="LCM" />
                <RESULT eventid="1212" points="456" swimtime="00:01:23.30" resultid="3291" heatid="4383" lane="3" entrytime="00:01:23.31" entrycourse="LCM" />
                <RESULT eventid="1266" points="386" swimtime="00:02:53.13" resultid="3292" heatid="4437" lane="2" entrytime="00:03:00.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" status="DSQ" swimtime="00:01:29.56" resultid="3293" heatid="4494" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabryel" lastname="Denk" birthdate="2011-05-09" gender="M" nation="BRA" license="391138" swrid="5602531" athleteid="3364" externalid="391138">
              <RESULTS>
                <RESULT eventid="1156" points="297" swimtime="00:01:10.22" resultid="3365" heatid="4335" lane="6" entrytime="00:01:17.49" entrycourse="LCM" />
                <RESULT eventid="1188" points="206" swimtime="00:00:43.92" resultid="3366" heatid="4364" lane="1" entrytime="00:00:49.85" entrycourse="LCM" />
                <RESULT eventid="1258" points="333" swimtime="00:20:55.61" resultid="3367" heatid="4431" lane="1" entrytime="00:21:59.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.03" />
                    <SPLIT distance="200" swimtime="00:02:41.80" />
                    <SPLIT distance="300" swimtime="00:04:06.09" />
                    <SPLIT distance="400" swimtime="00:05:29.76" />
                    <SPLIT distance="500" swimtime="00:06:54.38" />
                    <SPLIT distance="600" swimtime="00:08:18.64" />
                    <SPLIT distance="700" swimtime="00:09:43.38" />
                    <SPLIT distance="800" swimtime="00:11:06.60" />
                    <SPLIT distance="900" swimtime="00:12:30.80" />
                    <SPLIT distance="1000" swimtime="00:13:55.93" />
                    <SPLIT distance="1100" swimtime="00:15:20.01" />
                    <SPLIT distance="1200" swimtime="00:16:45.45" />
                    <SPLIT distance="1300" swimtime="00:18:09.53" />
                    <SPLIT distance="1400" swimtime="00:19:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" status="DSQ" swimtime="00:00:32.85" resultid="3368" heatid="4410" lane="4" entrytime="00:00:36.19" entrycourse="LCM" />
                <RESULT eventid="1306" points="254" swimtime="00:00:37.15" resultid="3369" heatid="4478" lane="5" entrytime="00:00:42.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcus" lastname="Vinicius De Almeida" birthdate="2009-06-16" gender="M" nation="BRA" license="348099" swrid="5600272" athleteid="3294" externalid="348099">
              <RESULTS>
                <RESULT eventid="1088" points="458" swimtime="00:02:42.68" resultid="3295" heatid="4288" lane="8" entrytime="00:02:44.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="534" swimtime="00:00:31.97" resultid="3296" heatid="4367" lane="4" entrytime="00:00:33.88" entrycourse="LCM" />
                <RESULT eventid="1220" points="475" swimtime="00:01:12.85" resultid="3297" heatid="4393" lane="6" entrytime="00:01:14.27" entrycourse="LCM" />
                <RESULT eventid="1306" points="456" swimtime="00:00:30.59" resultid="3298" heatid="4481" lane="7" entrytime="00:00:31.55" entrycourse="LCM" />
                <RESULT eventid="1374" points="472" swimtime="00:01:06.23" resultid="3299" heatid="4531" lane="1" entrytime="00:01:08.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="De Mello Araujo" birthdate="2010-11-03" gender="F" nation="BRA" license="406723" swrid="5717254" athleteid="3445" externalid="406723">
              <RESULTS>
                <RESULT eventid="1228" points="231" swimtime="00:00:38.45" resultid="3446" heatid="4396" lane="5" />
                <RESULT eventid="1212" points="183" swimtime="00:01:52.95" resultid="3447" heatid="4379" lane="7" entrytime="00:01:52.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduarda" lastname="Azevedo Birsneek" birthdate="2010-03-31" gender="F" nation="BRA" license="391145" swrid="5389427" athleteid="3383" externalid="391145">
              <RESULTS>
                <RESULT eventid="1064" points="197" swimtime="00:03:31.28" resultid="3384" heatid="4267" lane="4" entrytime="00:03:33.25" entrycourse="LCM" />
                <RESULT eventid="1096" points="120" swimtime="00:00:49.44" resultid="3385" heatid="4291" lane="3" entrytime="00:00:57.13" entrycourse="LCM" />
                <RESULT eventid="1148" points="200" swimtime="00:01:28.42" resultid="3386" heatid="4320" lane="3" entrytime="00:01:37.90" entrycourse="LCM" />
                <RESULT eventid="1298" points="203" swimtime="00:00:45.68" resultid="3387" heatid="4472" lane="1" entrytime="00:00:45.60" entrycourse="LCM" />
                <RESULT eventid="1366" points="189" swimtime="00:01:39.85" resultid="3388" heatid="4518" lane="5" entrytime="00:01:36.29" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaylane" lastname="Marques Ferreira" birthdate="2010-03-06" gender="F" nation="BRA" license="391146" swrid="5600211" athleteid="3389" externalid="391146">
              <RESULTS>
                <RESULT eventid="1096" points="346" swimtime="00:00:34.77" resultid="3390" heatid="4292" lane="7" entrytime="00:00:41.84" entrycourse="LCM" />
                <RESULT eventid="1148" points="269" swimtime="00:01:20.10" resultid="3391" heatid="4322" lane="1" entrytime="00:01:22.04" entrycourse="LCM" />
                <RESULT eventid="1228" points="319" swimtime="00:00:34.55" resultid="3392" heatid="4398" lane="6" entrytime="00:00:37.88" entrycourse="LCM" />
                <RESULT eventid="1282" points="224" swimtime="00:03:05.60" resultid="3393" heatid="4451" lane="1" entrytime="00:03:16.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="250" swimtime="00:01:27.96" resultid="3394" heatid="4494" lane="4" entrytime="00:01:43.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Vitor Navarro Zanini" birthdate="2008-06-30" gender="M" nation="BRA" license="369415" swrid="5600273" athleteid="3317" externalid="369415">
              <RESULTS>
                <RESULT eventid="1088" status="DSQ" swimtime="00:02:58.80" resultid="3318" heatid="4285" lane="3" entrytime="00:03:08.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="361" swimtime="00:00:36.42" resultid="3319" heatid="4365" lane="3" entrytime="00:00:39.53" entrycourse="LCM" />
                <RESULT eventid="1220" points="354" swimtime="00:01:20.37" resultid="3320" heatid="4390" lane="4" entrytime="00:01:23.36" entrycourse="LCM" />
                <RESULT eventid="1274" status="DSQ" swimtime="00:02:43.84" resultid="3321" heatid="4444" lane="7" entrytime="00:02:56.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1358" points="376" swimtime="00:05:04.77" resultid="3322" heatid="4512" lane="3" entrytime="00:05:29.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.72" />
                    <SPLIT distance="200" swimtime="00:02:30.26" />
                    <SPLIT distance="300" swimtime="00:03:49.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Liz Skowronski" birthdate="2008-01-24" gender="F" nation="BRA" license="358245" swrid="5600202" athleteid="3261" externalid="358245">
              <RESULTS>
                <RESULT eventid="1064" points="375" swimtime="00:02:50.61" resultid="3262" heatid="4270" lane="1" entrytime="00:02:49.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="307" swimtime="00:06:33.87" resultid="3263" heatid="4315" lane="7" entrytime="00:06:33.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.99" />
                    <SPLIT distance="200" swimtime="00:03:08.98" />
                    <SPLIT distance="300" swimtime="00:05:03.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1250" points="364" swimtime="00:11:18.75" resultid="3264" heatid="4427" lane="9" entrytime="00:11:13.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.02" />
                    <SPLIT distance="200" swimtime="00:02:38.26" />
                    <SPLIT distance="300" swimtime="00:04:04.68" />
                    <SPLIT distance="400" swimtime="00:05:30.33" />
                    <SPLIT distance="500" swimtime="00:06:56.41" />
                    <SPLIT distance="600" swimtime="00:08:24.23" />
                    <SPLIT distance="700" swimtime="00:09:52.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1298" points="368" swimtime="00:00:37.45" resultid="3265" heatid="4474" lane="3" entrytime="00:00:36.71" entrycourse="LCM" />
                <RESULT eventid="1366" points="361" swimtime="00:01:20.46" resultid="3266" heatid="4522" lane="7" entrytime="00:01:19.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Bilecki" birthdate="2007-05-28" gender="M" nation="BRA" license="406726" swrid="5717247" athleteid="3452" externalid="406726">
              <RESULTS>
                <RESULT eventid="1104" points="309" swimtime="00:00:32.94" resultid="3453" heatid="4296" lane="4" />
                <RESULT eventid="1156" points="357" swimtime="00:01:06.02" resultid="3454" heatid="4332" lane="7" />
                <RESULT eventid="1290" points="278" swimtime="00:02:36.26" resultid="3455" heatid="4459" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1342" status="DSQ" swimtime="00:01:19.15" resultid="3456" heatid="4500" lane="2" entrytime="00:01:17.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1204" points="267" swimtime="00:10:49.84" resultid="3470" heatid="4373" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.95" />
                    <SPLIT distance="200" swimtime="00:02:33.02" />
                    <SPLIT distance="300" swimtime="00:03:49.01" />
                    <SPLIT distance="400" swimtime="00:05:12.34" />
                    <SPLIT distance="500" swimtime="00:06:30.79" />
                    <SPLIT distance="600" swimtime="00:07:58.08" />
                    <SPLIT distance="700" swimtime="00:09:20.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3364" number="1" />
                    <RELAYPOSITION athleteid="3279" number="2" />
                    <RELAYPOSITION athleteid="3439" number="3" />
                    <RELAYPOSITION athleteid="3434" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="19" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1208" points="499" swimtime="00:08:47.67" resultid="3471" heatid="4375" lane="3" entrytime="00:09:07.36">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.14" />
                    <SPLIT distance="200" swimtime="00:02:09.12" />
                    <SPLIT distance="300" swimtime="00:03:10.94" />
                    <SPLIT distance="400" swimtime="00:04:21.53" />
                    <SPLIT distance="500" swimtime="00:05:24.28" />
                    <SPLIT distance="600" swimtime="00:06:34.71" />
                    <SPLIT distance="700" swimtime="00:07:36.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3329" number="1" />
                    <RELAYPOSITION athleteid="3257" number="2" />
                    <RELAYPOSITION athleteid="3404" number="3" />
                    <RELAYPOSITION athleteid="3267" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1206" points="438" swimtime="00:09:11.00" resultid="3472" heatid="4374" lane="9">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.71" />
                    <SPLIT distance="200" swimtime="00:02:12.13" />
                    <SPLIT distance="300" swimtime="00:03:18.84" />
                    <SPLIT distance="400" swimtime="00:04:36.24" />
                    <SPLIT distance="500" swimtime="00:05:44.74" />
                    <SPLIT distance="600" swimtime="00:06:58.90" />
                    <SPLIT distance="700" swimtime="00:08:03.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3294" number="1" />
                    <RELAYPOSITION athleteid="3340" number="2" />
                    <RELAYPOSITION athleteid="3317" number="3" />
                    <RELAYPOSITION athleteid="3273" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1326" points="217" swimtime="00:05:43.84" resultid="3473" heatid="4489" lane="7" entrytime="00:05:28.10">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.33" />
                    <SPLIT distance="200" swimtime="00:02:57.68" />
                    <SPLIT distance="300" swimtime="00:04:23.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3364" number="1" />
                    <RELAYPOSITION athleteid="3279" number="2" />
                    <RELAYPOSITION athleteid="3439" number="3" />
                    <RELAYPOSITION athleteid="3284" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1328" points="355" swimtime="00:04:51.76" resultid="3474" heatid="4490" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                    <SPLIT distance="200" swimtime="00:02:28.14" />
                    <SPLIT distance="300" swimtime="00:03:46.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3273" number="1" />
                    <RELAYPOSITION athleteid="3294" number="2" />
                    <RELAYPOSITION athleteid="3423" number="3" />
                    <RELAYPOSITION athleteid="3340" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1396" points="363" swimtime="00:04:23.75" resultid="3477" heatid="4541" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.43" />
                    <SPLIT distance="200" swimtime="00:02:00.38" />
                    <SPLIT distance="300" swimtime="00:03:19.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3294" number="1" />
                    <RELAYPOSITION athleteid="3273" number="2" />
                    <RELAYPOSITION athleteid="3423" number="3" />
                    <RELAYPOSITION athleteid="3340" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1332" points="425" swimtime="00:04:34.86" resultid="3475" heatid="4492" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.39" />
                    <SPLIT distance="200" swimtime="00:02:33.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3404" number="1" />
                    <RELAYPOSITION athleteid="3257" number="2" />
                    <RELAYPOSITION athleteid="3267" number="3" />
                    <RELAYPOSITION athleteid="3329" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1400" points="539" swimtime="00:03:51.24" resultid="3476" heatid="4543" lane="6" entrytime="00:04:00.82">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.09" />
                    <SPLIT distance="200" swimtime="00:01:56.52" />
                    <SPLIT distance="300" swimtime="00:02:55.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3404" number="1" />
                    <RELAYPOSITION athleteid="3257" number="2" />
                    <RELAYPOSITION athleteid="3267" number="3" />
                    <RELAYPOSITION athleteid="3329" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1196" points="318" swimtime="00:11:09.67" resultid="3463" heatid="4370" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.15" />
                    <SPLIT distance="200" swimtime="00:02:38.83" />
                    <SPLIT distance="300" swimtime="00:04:05.47" />
                    <SPLIT distance="400" swimtime="00:05:43.53" />
                    <SPLIT distance="500" swimtime="00:06:55.85" />
                    <SPLIT distance="600" swimtime="00:08:20.38" />
                    <SPLIT distance="700" swimtime="00:09:39.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3288" number="1" />
                    <RELAYPOSITION athleteid="3389" number="2" />
                    <RELAYPOSITION athleteid="3323" number="3" />
                    <RELAYPOSITION athleteid="3300" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="F" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1198" points="420" swimtime="00:10:10.67" resultid="3464" heatid="4371" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.34" />
                    <SPLIT distance="200" swimtime="00:02:26.15" />
                    <SPLIT distance="300" swimtime="00:03:40.31" />
                    <SPLIT distance="500" swimtime="00:06:19.71" />
                    <SPLIT distance="600" swimtime="00:07:42.14" />
                    <SPLIT distance="700" swimtime="00:08:52.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3410" number="1" />
                    <RELAYPOSITION athleteid="3416" number="2" />
                    <RELAYPOSITION athleteid="3261" number="3" />
                    <RELAYPOSITION athleteid="3352" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1316" points="272" swimtime="00:05:55.27" resultid="3465" heatid="4484" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.69" />
                    <SPLIT distance="200" swimtime="00:02:52.27" />
                    <SPLIT distance="300" swimtime="00:04:20.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3323" number="1" />
                    <RELAYPOSITION athleteid="3288" number="2" />
                    <RELAYPOSITION athleteid="3389" number="3" />
                    <RELAYPOSITION athleteid="3383" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1384" points="286" swimtime="00:05:15.43" resultid="3469" heatid="4535" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.55" />
                    <SPLIT distance="200" swimtime="00:02:23.24" />
                    <SPLIT distance="300" swimtime="00:03:42.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3288" number="1" />
                    <RELAYPOSITION athleteid="3323" number="2" />
                    <RELAYPOSITION athleteid="3389" number="3" />
                    <RELAYPOSITION athleteid="3383" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1320" points="317" swimtime="00:05:37.58" resultid="3466" heatid="4486" lane="3">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:02:52.61" />
                    <SPLIT distance="300" swimtime="00:04:23.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3352" number="1" />
                    <RELAYPOSITION athleteid="3410" number="2" />
                    <RELAYPOSITION athleteid="3261" number="3" />
                    <RELAYPOSITION athleteid="3395" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1388" points="421" swimtime="00:04:37.31" resultid="3467" heatid="4537" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.54" />
                    <SPLIT distance="200" swimtime="00:02:16.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3410" number="1" />
                    <RELAYPOSITION athleteid="3261" number="2" />
                    <RELAYPOSITION athleteid="3395" number="3" />
                    <RELAYPOSITION athleteid="3352" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="F" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1390" points="355" swimtime="00:04:53.48" resultid="3468" heatid="4538" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3306" number="1" />
                    <RELAYPOSITION athleteid="3370" number="2" />
                    <RELAYPOSITION athleteid="3378" number="3" />
                    <RELAYPOSITION athleteid="3346" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1248" points="349" swimtime="00:05:09.03" resultid="3478" heatid="4425" lane="3" entrytime="00:05:01.80">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.53" />
                    <SPLIT distance="200" swimtime="00:02:51.04" />
                    <SPLIT distance="300" swimtime="00:03:56.51" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3306" number="1" />
                    <RELAYPOSITION athleteid="3252" number="2" />
                    <RELAYPOSITION athleteid="3329" number="3" />
                    <RELAYPOSITION athleteid="3346" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1246" points="369" swimtime="00:05:03.15" resultid="3479" heatid="4424" lane="6" entrytime="00:05:03.44">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3352" number="1" />
                    <RELAYPOSITION athleteid="3317" number="2" />
                    <RELAYPOSITION athleteid="3457" number="3" />
                    <RELAYPOSITION athleteid="3410" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="16816" nation="BRA" region="SC" clubid="3778" swrid="94375" name="Jurerê Sports Center" shortname="Swimfloripa - Jurerê">
          <ATHLETES>
            <ATHLETE firstname="José" lastname="Roberto Vaz Guimarães Neto" birthdate="1996-11-14" gender="M" nation="BRA" license="109462" swrid="5206816" athleteid="3779" externalid="109462">
              <RESULTS>
                <RESULT eventid="1104" points="736" status="EXH" swimtime="00:00:24.66" resultid="3780" heatid="4304" lane="4" entrytime="00:00:24.75" entrycourse="LCM" />
                <RESULT eventid="1236" points="689" status="EXH" swimtime="00:00:23.67" resultid="3781" heatid="4422" lane="5" entrytime="00:00:23.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3133" nation="BRA" region="PR" clubid="3782" swrid="93768" name="Associação Toledo Natação" shortname="Toledo Natação">
          <ATHLETES>
            <ATHLETE firstname="Gabriel" lastname="Marafon" birthdate="2006-06-17" gender="M" nation="BRA" license="380288" swrid="5622291" athleteid="3800" externalid="380288">
              <RESULTS>
                <RESULT eventid="1088" points="373" swimtime="00:02:54.25" resultid="3801" heatid="4287" lane="1" entrytime="00:02:52.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="490" swimtime="00:00:32.90" resultid="3802" heatid="4367" lane="5" entrytime="00:00:34.13" entrycourse="LCM" />
                <RESULT eventid="1220" points="379" swimtime="00:01:18.54" resultid="3803" heatid="4392" lane="4" entrytime="00:01:15.75" entrycourse="LCM" />
                <RESULT eventid="1236" points="425" swimtime="00:00:27.80" resultid="3804" heatid="4417" lane="6" entrytime="00:00:27.45" entrycourse="LCM" />
                <RESULT eventid="1290" points="362" swimtime="00:02:23.06" resultid="3805" heatid="4459" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrielly" lastname="Luiza Horn" birthdate="2004-04-03" gender="F" nation="BRA" license="315145" swrid="5622288" athleteid="3788" externalid="315145">
              <RESULTS>
                <RESULT eventid="1096" points="372" swimtime="00:00:33.94" resultid="3789" heatid="4293" lane="5" entrytime="00:00:34.81" entrycourse="LCM" />
                <RESULT eventid="1180" points="338" swimtime="00:00:41.85" resultid="3790" heatid="4357" lane="2" entrytime="00:00:43.56" entrycourse="LCM" />
                <RESULT eventid="1228" points="378" swimtime="00:00:32.64" resultid="3791" heatid="4402" lane="8" entrytime="00:00:31.74" entrycourse="LCM" />
                <RESULT eventid="1298" points="379" swimtime="00:00:37.08" resultid="3792" heatid="4473" lane="4" entrytime="00:00:37.68" entrycourse="LCM" />
                <RESULT eventid="1366" points="299" swimtime="00:01:25.66" resultid="3793" heatid="4517" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Marafon" birthdate="2011-03-23" gender="F" nation="BRA" license="380287" swrid="5652623" athleteid="3821" externalid="380287">
              <RESULTS>
                <RESULT eventid="1080" points="331" swimtime="00:03:18.75" resultid="3822" heatid="4278" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:52.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="423" swimtime="00:01:08.85" resultid="3823" heatid="4320" lane="7" />
                <RESULT eventid="1180" points="377" swimtime="00:00:40.33" resultid="3824" heatid="4356" lane="8" />
                <RESULT eventid="1228" points="410" swimtime="00:00:31.78" resultid="3825" heatid="4396" lane="6" />
                <RESULT eventid="1212" points="362" swimtime="00:01:29.95" resultid="3826" heatid="4377" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Welter Levandowski" birthdate="2011-05-06" gender="F" nation="BRA" license="380286" swrid="5652626" athleteid="3816" externalid="380286">
              <RESULTS>
                <RESULT eventid="1096" points="259" swimtime="00:00:38.31" resultid="3817" heatid="4291" lane="6" />
                <RESULT eventid="1164" points="206" swimtime="00:03:26.18" resultid="3818" heatid="4349" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="360" swimtime="00:02:38.63" resultid="3819" heatid="4449" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1334" points="238" swimtime="00:01:29.45" resultid="3820" heatid="4493" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Feder" birthdate="2008-11-13" gender="M" nation="BRA" license="347224" swrid="5622278" athleteid="3783" externalid="347224">
              <RESULTS>
                <RESULT eventid="1072" points="397" swimtime="00:02:32.21" resultid="3784" heatid="4275" lane="1" entrytime="00:02:35.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="495" swimtime="00:00:28.15" resultid="3785" heatid="4297" lane="3" />
                <RESULT eventid="1306" points="467" swimtime="00:00:30.34" resultid="3786" heatid="4481" lane="3" entrytime="00:00:30.96" entrycourse="LCM" />
                <RESULT eventid="1374" points="437" swimtime="00:01:07.96" resultid="3787" heatid="4531" lane="6" entrytime="00:01:08.11" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Torres Romancini" birthdate="2010-05-28" gender="F" nation="BRA" license="347218" swrid="5622309" athleteid="3806" externalid="347218">
              <RESULTS>
                <RESULT eventid="1064" points="388" swimtime="00:02:48.70" resultid="3807" heatid="4267" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="352" swimtime="00:00:34.57" resultid="3808" heatid="4293" lane="1" entrytime="00:00:36.81" entrycourse="LCM" />
                <RESULT eventid="1228" points="399" swimtime="00:00:32.07" resultid="3809" heatid="4399" lane="4" entrytime="00:00:33.62" entrycourse="LCM" />
                <RESULT eventid="1298" points="465" swimtime="00:00:34.67" resultid="3810" heatid="4474" lane="8" entrytime="00:00:37.52" entrycourse="LCM" />
                <RESULT eventid="1366" points="418" swimtime="00:01:16.66" resultid="3811" heatid="4521" lane="5" entrytime="00:01:21.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lavinia" lastname="Martins Paludo" birthdate="2010-09-30" gender="F" nation="BRA" license="347217" swrid="5652624" athleteid="3812" externalid="347217">
              <RESULTS>
                <RESULT eventid="1080" status="DSQ" swimtime="00:03:46.59" resultid="3813" heatid="4279" lane="8" entrytime="00:03:40.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="233" swimtime="00:00:47.35" resultid="3814" heatid="4357" lane="7" entrytime="00:00:45.47" entrycourse="LCM" />
                <RESULT eventid="1212" points="231" swimtime="00:01:44.43" resultid="3815" heatid="4380" lane="7" entrytime="00:01:43.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giullia" lastname="Lagni" birthdate="2006-11-22" gender="F" nation="BRA" license="337671" swrid="5622285" athleteid="3794" externalid="337671">
              <RESULTS>
                <RESULT eventid="1064" points="342" swimtime="00:02:56.02" resultid="3795" heatid="4267" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="368" swimtime="00:01:12.14" resultid="3796" heatid="4323" lane="1" entrytime="00:01:14.48" entrycourse="LCM" />
                <RESULT eventid="1228" points="369" swimtime="00:00:32.91" resultid="3797" heatid="4399" lane="5" entrytime="00:00:33.65" entrycourse="LCM" />
                <RESULT eventid="1298" points="383" swimtime="00:00:36.97" resultid="3798" heatid="4471" lane="8" />
                <RESULT eventid="1366" points="354" swimtime="00:01:21.00" resultid="3799" heatid="4517" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="ASSOCIAÇÃO TOLEDO NATAÇAO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1316" points="319" swimtime="00:05:37.18" resultid="3827" heatid="4484" lane="7">
                  <SPLITS>
                    <SPLIT distance="200" swimtime="00:02:43.76" />
                    <SPLIT distance="300" swimtime="00:04:16.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3806" number="1" />
                    <RELAYPOSITION athleteid="3821" number="2" />
                    <RELAYPOSITION athleteid="3816" number="3" />
                    <RELAYPOSITION athleteid="3812" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1384" points="352" swimtime="00:04:54.44" resultid="3828" heatid="4535" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.61" />
                    <SPLIT distance="200" swimtime="00:02:24.22" />
                    <SPLIT distance="300" swimtime="00:03:45.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3806" number="1" />
                    <RELAYPOSITION athleteid="3816" number="2" />
                    <RELAYPOSITION athleteid="3812" number="3" />
                    <RELAYPOSITION athleteid="3821" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
