<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.79125">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Maringá" name="Torneio Regional da 2ª Região (Pré-Mirim/Sênior)" course="SCM" deadline="2024-03-04" entrystartdate="2024-02-28" entrytype="INVITATION" hostclub="Universidade Estadual de Maringá" hostclub.url="http://www.uem.br/" number="38298" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/evento/natacao/38298" startmethod="2" timing="AUTOMATIC" masters="F" withdrawuntil="2024-03-06" state="PR" nation="BRA">
      <AGEDATE value="2024-03-09" type="YEAR" />
      <POOL name="Universidade Estadual de Maringá" lanemin="1" lanemax="6" />
      <FACILITY city="Maringá" name="Universidade Estadual de Maringá" nation="BRA" state="PR" street="M19" street2="Vila Esperança" zip="87020-900" />
      <POINTTABLE pointtableid="3016" name="FINA Point Scoring" version="2023" />
      <QUALIFY from="2023-03-09" until="2024-03-08" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99206-4448" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99206-4448" street="Avenida do Batel, 1230" street2="Batel" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-03-09" daytime="09:10" endtime="11:58" number="1" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1060" daytime="09:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1780" />
                    <RANKING order="2" place="2" resultid="1364" />
                    <RANKING order="3" place="3" resultid="1473" />
                    <RANKING order="4" place="4" resultid="1677" />
                    <RANKING order="5" place="5" resultid="1494" />
                    <RANKING order="6" place="6" resultid="1518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1735" />
                    <RANKING order="2" place="2" resultid="1751" />
                    <RANKING order="3" place="3" resultid="1490" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1871" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1872" daytime="09:14" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1063" daytime="09:20" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1064" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1835" />
                    <RANKING order="2" place="2" resultid="1502" />
                    <RANKING order="3" place="3" resultid="1577" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1506" />
                    <RANKING order="2" place="2" resultid="1498" />
                    <RANKING order="3" place="3" resultid="1776" />
                    <RANKING order="4" place="4" resultid="1510" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1873" daytime="09:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1874" daytime="09:24" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1066" daytime="09:28" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1067" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1368" />
                    <RANKING order="2" place="2" resultid="1469" />
                    <RANKING order="3" place="3" resultid="1555" />
                    <RANKING order="4" place="4" resultid="1965" />
                    <RANKING order="5" place="-1" resultid="1802" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1529" />
                    <RANKING order="2" place="2" resultid="1686" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1070" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1071" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1072" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1073" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1875" daytime="09:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1960" daytime="09:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1074" daytime="09:38" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1075" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1463" />
                    <RANKING order="2" place="2" resultid="1762" />
                    <RANKING order="3" place="3" resultid="1405" />
                    <RANKING order="4" place="4" resultid="1738" />
                    <RANKING order="5" place="-1" resultid="1787" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1076" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1387" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1077" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1745" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1438" />
                    <RANKING order="2" place="2" resultid="1699" />
                    <RANKING order="3" place="3" resultid="1400" />
                    <RANKING order="4" place="4" resultid="1559" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1080" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1081" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1681" />
                    <RANKING order="2" place="-1" resultid="1379" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1876" daytime="09:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1877" daytime="09:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1878" daytime="09:46" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1082" daytime="09:52" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1083" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1602" />
                    <RANKING order="2" place="2" resultid="1759" />
                    <RANKING order="3" place="3" resultid="1794" />
                    <RANKING order="4" place="4" resultid="1755" />
                    <RANKING order="5" place="5" resultid="1676" />
                    <RANKING order="6" place="-1" resultid="1823" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1705" />
                    <RANKING order="2" place="2" resultid="1514" />
                    <RANKING order="3" place="3" resultid="1552" />
                    <RANKING order="4" place="4" resultid="1486" />
                    <RANKING order="5" place="-1" resultid="1723" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1879" daytime="09:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1880" daytime="09:54" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1085" daytime="09:58" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1086" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1573" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1775" />
                    <RANKING order="2" place="2" resultid="1505" />
                    <RANKING order="3" place="3" resultid="1727" />
                    <RANKING order="4" place="4" resultid="1719" />
                    <RANKING order="5" place="5" resultid="1610" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1881" daytime="09:58" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1088" daytime="10:02" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1089" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1468" />
                    <RANKING order="2" place="2" resultid="1476" />
                    <RANKING order="3" place="3" resultid="1357" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1345" />
                    <RANKING order="2" place="2" resultid="1534" />
                    <RANKING order="3" place="3" resultid="1339" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1427" />
                    <RANKING order="2" place="2" resultid="1432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1092" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1327" />
                    <RANKING order="2" place="2" resultid="1447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1093" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1333" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1415" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1882" daytime="10:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1883" daytime="10:06" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1096" daytime="10:08" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1097" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1459" />
                    <RANKING order="2" place="2" resultid="1737" />
                    <RANKING order="3" place="3" resultid="1351" />
                    <RANKING order="4" place="4" resultid="1848" />
                    <RANKING order="5" place="5" resultid="1797" />
                    <RANKING order="6" place="-1" resultid="1786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1712" />
                    <RANKING order="2" place="-1" resultid="1584" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1744" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1392" />
                    <RANKING order="2" place="2" resultid="1558" />
                    <RANKING order="3" place="3" resultid="1698" />
                    <RANKING order="4" place="4" resultid="1692" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1321" />
                    <RANKING order="2" place="2" resultid="1659" />
                    <RANKING order="3" place="-1" resultid="1525" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1374" />
                    <RANKING order="2" place="2" resultid="1452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1884" daytime="10:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1885" daytime="10:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1886" daytime="10:14" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1104" daytime="10:16" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1105" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1754" />
                    <RANKING order="2" place="2" resultid="1822" />
                    <RANKING order="3" place="3" resultid="1472" />
                    <RANKING order="4" place="4" resultid="1675" />
                    <RANKING order="5" place="5" resultid="1493" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1722" />
                    <RANKING order="2" place="2" resultid="1489" />
                    <RANKING order="3" place="3" resultid="1839" />
                    <RANKING order="4" place="4" resultid="1513" />
                    <RANKING order="5" place="5" resultid="1869" />
                    <RANKING order="6" place="6" resultid="1551" />
                    <RANKING order="7" place="7" resultid="1815" />
                    <RANKING order="8" place="8" resultid="1540" />
                    <RANKING order="9" place="9" resultid="1485" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1887" daytime="10:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1888" daytime="10:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1889" daytime="10:22" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1107" daytime="10:24" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1108" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1501" />
                    <RANKING order="2" place="2" resultid="1576" />
                    <RANKING order="3" place="3" resultid="1581" />
                    <RANKING order="4" place="-1" resultid="1772" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1726" />
                    <RANKING order="2" place="2" resultid="1718" />
                    <RANKING order="3" place="3" resultid="1482" />
                    <RANKING order="4" place="4" resultid="1831" />
                    <RANKING order="5" place="5" resultid="1509" />
                    <RANKING order="6" place="6" resultid="1569" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1890" daytime="10:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1891" daytime="10:26" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1110" daytime="10:30" gender="F" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1111" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1112" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1685" />
                    <RANKING order="2" place="2" resultid="1528" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1114" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1115" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1117" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1892" daytime="10:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1118" daytime="10:48" gender="M" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1119" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1120" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1122" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1123" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1124" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1125" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1893" daytime="10:48" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1126" daytime="11:24" gender="F" number="13" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1127" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1758" />
                    <RANKING order="2" place="2" resultid="1779" />
                    <RANKING order="3" place="3" resultid="1601" />
                    <RANKING order="4" place="4" resultid="1517" />
                    <RANKING order="5" place="-1" resultid="1709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1734" />
                    <RANKING order="2" place="2" resultid="1838" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1894" daytime="11:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1895" daytime="11:26" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1129" daytime="11:30" gender="M" number="14" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1130" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1580" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="12" agemin="12" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1896" daytime="11:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1132" daytime="11:32" gender="F" number="15" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1133" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1367" />
                    <RANKING order="2" place="2" resultid="1554" />
                    <RANKING order="3" place="3" resultid="1475" />
                    <RANKING order="4" place="4" resultid="1356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1134" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1135" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1137" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1663" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1139" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1897" daytime="11:32" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1140" daytime="11:34" gender="M" number="16" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1141" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1671" />
                    <RANKING order="2" place="2" resultid="1854" />
                    <RANKING order="3" place="3" resultid="1796" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1143" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1144" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1437" />
                    <RANKING order="2" place="2" resultid="1391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1658" />
                    <RANKING order="2" place="-1" resultid="1524" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1147" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1411" />
                    <RANKING order="2" place="2" resultid="1680" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1898" daytime="11:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1899" daytime="11:38" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1148" daytime="11:40" gender="F" number="17" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1149" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1757" />
                    <RANKING order="2" place="2" resultid="1363" />
                    <RANKING order="3" place="3" resultid="1471" />
                    <RANKING order="4" place="4" resultid="1753" />
                    <RANKING order="5" place="4" resultid="1793" />
                    <RANKING order="6" place="6" resultid="1492" />
                    <RANKING order="7" place="-1" resultid="1708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1733" />
                    <RANKING order="2" place="2" resultid="1488" />
                    <RANKING order="3" place="3" resultid="1704" />
                    <RANKING order="4" place="4" resultid="1750" />
                    <RANKING order="5" place="5" resultid="1550" />
                    <RANKING order="6" place="6" resultid="1539" />
                    <RANKING order="7" place="-1" resultid="1814" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1900" daytime="11:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1901" daytime="11:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1902" daytime="11:46" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1151" daytime="11:50" gender="M" number="18" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1152" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1500" />
                    <RANKING order="2" place="2" resultid="1834" />
                    <RANKING order="3" place="3" resultid="1575" />
                    <RANKING order="4" place="4" resultid="1572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1504" />
                    <RANKING order="2" place="2" resultid="1497" />
                    <RANKING order="3" place="3" resultid="1481" />
                    <RANKING order="4" place="4" resultid="1774" />
                    <RANKING order="5" place="5" resultid="1568" />
                    <RANKING order="6" place="6" resultid="1609" />
                    <RANKING order="7" place="-1" resultid="1830" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1903" daytime="11:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1904" daytime="11:52" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1154" daytime="11:56" gender="F" number="19" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1155" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1467" />
                    <RANKING order="2" place="2" resultid="1801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1533" />
                    <RANKING order="2" place="2" resultid="1344" />
                    <RANKING order="3" place="3" resultid="1338" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1158" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1420" />
                    <RANKING order="2" place="2" resultid="1326" />
                    <RANKING order="3" place="3" resultid="1446" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1160" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1161" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1905" daytime="11:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1906" daytime="11:58" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1162" daytime="12:02" gender="M" number="20" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1163" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1458" />
                    <RANKING order="2" place="2" resultid="1761" />
                    <RANKING order="3" place="3" resultid="1670" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1164" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1165" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1382" />
                    <RANKING order="2" place="2" resultid="1442" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1424" />
                    <RANKING order="2" place="2" resultid="1451" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1907" daytime="12:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1908" daytime="12:04" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1170" daytime="12:08" gender="F" number="21" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1171" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1600" />
                    <RANKING order="2" place="2" resultid="1362" />
                    <RANKING order="3" place="3" resultid="1778" />
                    <RANKING order="4" place="4" resultid="1821" />
                    <RANKING order="5" place="5" resultid="1792" />
                    <RANKING order="6" place="6" resultid="1516" />
                    <RANKING order="7" place="-1" resultid="1707" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1721" />
                    <RANKING order="2" place="2" resultid="1512" />
                    <RANKING order="3" place="3" resultid="1703" />
                    <RANKING order="4" place="4" resultid="1837" />
                    <RANKING order="5" place="5" resultid="1868" />
                    <RANKING order="6" place="6" resultid="1749" />
                    <RANKING order="7" place="7" resultid="1538" />
                    <RANKING order="8" place="8" resultid="1484" />
                    <RANKING order="9" place="9" resultid="1813" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1909" daytime="12:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1910" daytime="12:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1911" daytime="12:10" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1173" daytime="12:12" gender="M" number="22" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1174" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1833" />
                    <RANKING order="2" place="2" resultid="1579" />
                    <RANKING order="3" place="3" resultid="1571" />
                    <RANKING order="4" place="4" resultid="1771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1496" />
                    <RANKING order="2" place="2" resultid="1725" />
                    <RANKING order="3" place="3" resultid="1480" />
                    <RANKING order="4" place="3" resultid="1717" />
                    <RANKING order="5" place="5" resultid="1508" />
                    <RANKING order="6" place="6" resultid="1829" />
                    <RANKING order="7" place="7" resultid="1567" />
                    <RANKING order="8" place="8" resultid="1608" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1912" daytime="12:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1913" daytime="12:14" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1176" daytime="12:18" gender="F" number="23" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1177" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1179" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1180" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1181" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1182" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1183" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1966" daytime="12:18" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1184" daytime="12:20" gender="M" number="24" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1185" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1462" />
                    <RANKING order="2" place="2" resultid="1404" />
                    <RANKING order="3" place="3" resultid="1350" />
                    <RANKING order="4" place="4" resultid="1669" />
                    <RANKING order="5" place="-1" resultid="1853" />
                    <RANKING order="6" place="-1" resultid="1847" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1711" />
                    <RANKING order="2" place="-1" resultid="1583" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1396" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1188" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1436" />
                    <RANKING order="2" place="2" resultid="1691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1189" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1190" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1191" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1378" />
                    <RANKING order="2" place="2" resultid="1679" />
                    <RANKING order="3" place="-1" resultid="1409" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1914" daytime="12:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1915" daytime="12:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1916" daytime="12:22" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-03-09" daytime="15:40" endtime="17:40" number="2" officialmeeting="15:00" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1192" daytime="15:40" gender="F" number="25" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1193" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1194" daytime="15:40" gender="M" number="26" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1195" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1858" />
                    <RANKING order="2" place="2" resultid="1643" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1917" daytime="15:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1196" daytime="15:42" gender="F" number="27" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1197" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1594" />
                    <RANKING order="2" place="2" resultid="1623" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1731" />
                    <RANKING order="2" place="2" resultid="1769" />
                    <RANKING order="3" place="3" resultid="1627" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1918" daytime="15:42" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1199" daytime="15:46" gender="M" number="28" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1200" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1784" />
                    <RANKING order="2" place="2" resultid="1638" />
                    <RANKING order="3" place="3" resultid="1565" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1201" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1544" />
                    <RANKING order="2" place="2" resultid="1827" />
                    <RANKING order="3" place="3" resultid="1656" />
                    <RANKING order="4" place="4" resultid="1617" />
                    <RANKING order="5" place="5" resultid="1845" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1919" daytime="15:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1920" daytime="15:48" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1202" daytime="15:52" gender="F" number="29" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1203" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1360" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1204" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1536" />
                    <RANKING order="2" place="2" resultid="1689" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1205" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1429" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1206" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1422" />
                    <RANKING order="2" place="2" resultid="1449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1336" />
                    <RANKING order="2" place="2" resultid="1667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1921" daytime="15:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1922" daytime="15:58" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1210" daytime="16:04" gender="M" number="30" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1211" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1741" />
                    <RANKING order="2" place="-1" resultid="1790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1212" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1389" />
                    <RANKING order="2" place="2" resultid="1715" />
                    <RANKING order="3" place="3" resultid="1456" />
                    <RANKING order="4" place="-1" resultid="1586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1213" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1384" />
                    <RANKING order="2" place="2" resultid="1747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1216" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1683" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1923" daytime="16:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1924" daytime="16:12" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1218" daytime="16:18" gender="F" number="31" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1219" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1220" daytime="16:18" gender="M" number="32" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1221" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1642" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1925" daytime="16:18" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1222" daytime="16:20" gender="F" number="33" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1223" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1593" />
                    <RANKING order="2" place="2" resultid="1622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1224" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1730" />
                    <RANKING order="2" place="2" resultid="1631" />
                    <RANKING order="3" place="3" resultid="1819" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1926" daytime="16:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1225" daytime="16:24" gender="M" number="34" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1226" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1606" />
                    <RANKING order="2" place="2" resultid="1564" />
                    <RANKING order="3" place="3" resultid="1598" />
                    <RANKING order="4" place="-1" resultid="1807" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1227" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1548" />
                    <RANKING order="2" place="2" resultid="1590" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1927" daytime="16:24" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1228" daytime="16:26" gender="F" number="35" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1229" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1974" />
                    <RANKING order="2" place="2" resultid="1805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1531" />
                    <RANKING order="2" place="2" resultid="1688" />
                    <RANKING order="3" place="3" resultid="1348" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1232" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1235" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1928" daytime="16:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1973" daytime="16:28" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1236" daytime="16:32" gender="M" number="36" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1237" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1465" />
                    <RANKING order="2" place="2" resultid="1407" />
                    <RANKING order="3" place="3" resultid="1765" />
                    <RANKING order="4" place="4" resultid="1354" />
                    <RANKING order="5" place="-1" resultid="1851" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1238" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1714" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1239" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1398" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1240" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1402" />
                    <RANKING order="2" place="2" resultid="1695" />
                    <RANKING order="3" place="3" resultid="1561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1241" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1243" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1380" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1929" daytime="16:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1930" daytime="16:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1244" daytime="16:38" gender="F" number="37" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1245" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1246" daytime="16:38" gender="M" number="38" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1247" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1641" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1931" daytime="16:38" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1248" daytime="16:56" gender="F" number="39" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1249" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1634" />
                    <RANKING order="2" place="2" resultid="1613" />
                    <RANKING order="3" place="-1" resultid="1811" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1250" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1626" />
                    <RANKING order="2" place="2" resultid="1768" />
                    <RANKING order="3" place="3" resultid="1522" />
                    <RANKING order="4" place="4" resultid="1620" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1932" daytime="16:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1933" daytime="16:58" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1251" daytime="17:02" gender="M" number="40" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1252" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1783" />
                    <RANKING order="2" place="2" resultid="1597" />
                    <RANKING order="3" place="3" resultid="1649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1253" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1543" />
                    <RANKING order="2" place="2" resultid="1646" />
                    <RANKING order="3" place="3" resultid="1652" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1934" daytime="17:02" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1254" daytime="17:04" gender="F" number="41" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1255" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1371" />
                    <RANKING order="2" place="2" resultid="1478" />
                    <RANKING order="3" place="3" resultid="1359" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1256" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1257" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1258" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1666" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1261" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1935" daytime="17:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1936" daytime="17:06" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1262" daytime="17:08" gender="M" number="42" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1263" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1764" />
                    <RANKING order="2" place="2" resultid="1673" />
                    <RANKING order="3" place="3" resultid="1353" />
                    <RANKING order="4" place="-1" resultid="1850" />
                    <RANKING order="5" place="-1" resultid="1799" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1265" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1444" />
                    <RANKING order="2" place="2" resultid="1397" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1700" />
                    <RANKING order="2" place="2" resultid="1694" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1267" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1268" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1375" />
                    <RANKING order="2" place="2" resultid="1425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1269" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1413" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1937" daytime="17:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1938" daytime="17:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1270" daytime="17:12" gender="F" number="43" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1271" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1862" />
                    <RANKING order="2" place="2" resultid="1860" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1939" daytime="17:12" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1272" daytime="17:14" gender="M" number="44" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1273" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1857" />
                    <RANKING order="2" place="2" resultid="1640" />
                    <RANKING order="3" place="3" resultid="1864" />
                    <RANKING order="4" place="4" resultid="1866" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1940" daytime="17:14" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1274" daytime="17:16" gender="F" number="45" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1275" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1592" />
                    <RANKING order="2" place="-1" resultid="1810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1729" />
                    <RANKING order="2" place="2" resultid="1630" />
                    <RANKING order="3" place="3" resultid="1521" />
                    <RANKING order="4" place="4" resultid="1818" />
                    <RANKING order="5" place="5" resultid="1842" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1941" daytime="17:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1942" daytime="17:18" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1277" daytime="17:20" gender="M" number="46" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1278" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1605" />
                    <RANKING order="2" place="2" resultid="1637" />
                    <RANKING order="3" place="3" resultid="1563" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1542" />
                    <RANKING order="2" place="2" resultid="1826" />
                    <RANKING order="3" place="3" resultid="1655" />
                    <RANKING order="4" place="4" resultid="1589" />
                    <RANKING order="5" place="5" resultid="1844" />
                    <RANKING order="6" place="6" resultid="1547" />
                    <RANKING order="7" place="7" resultid="1616" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1943" daytime="17:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1944" daytime="17:22" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1280" daytime="17:26" gender="F" number="47" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1281" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1370" />
                    <RANKING order="2" place="2" resultid="1804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1282" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1530" />
                    <RANKING order="2" place="2" resultid="1341" />
                    <RANKING order="3" place="3" resultid="1347" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1283" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1428" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1284" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1329" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1665" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1286" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1417" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1287" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1945" daytime="17:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1946" daytime="17:28" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1288" daytime="17:32" gender="M" number="48" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1289" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1460" />
                    <RANKING order="2" place="2" resultid="1740" />
                    <RANKING order="3" place="3" resultid="1672" />
                    <RANKING order="4" place="-1" resultid="1789" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1290" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1388" />
                    <RANKING order="2" place="2" resultid="1455" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1291" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1746" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1440" />
                    <RANKING order="2" place="2" resultid="1394" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1293" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1323" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1294" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1295" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1947" daytime="17:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1948" daytime="17:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1296" daytime="17:38" gender="F" number="49" order="26" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1297" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1633" />
                    <RANKING order="2" place="2" resultid="1612" />
                    <RANKING order="3" place="-1" resultid="1809" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1298" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1767" />
                    <RANKING order="2" place="2" resultid="1629" />
                    <RANKING order="3" place="3" resultid="1625" />
                    <RANKING order="4" place="4" resultid="1841" />
                    <RANKING order="5" place="5" resultid="1520" />
                    <RANKING order="6" place="6" resultid="1817" />
                    <RANKING order="7" place="7" resultid="1619" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1949" daytime="17:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1950" daytime="17:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1299" daytime="17:42" gender="M" number="50" order="27" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1300" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1782" />
                    <RANKING order="2" place="2" resultid="1596" />
                    <RANKING order="3" place="3" resultid="1604" />
                    <RANKING order="4" place="4" resultid="1636" />
                    <RANKING order="5" place="5" resultid="1648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1301" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1546" />
                    <RANKING order="2" place="2" resultid="1825" />
                    <RANKING order="3" place="3" resultid="1654" />
                    <RANKING order="4" place="4" resultid="1615" />
                    <RANKING order="5" place="5" resultid="1588" />
                    <RANKING order="6" place="6" resultid="1645" />
                    <RANKING order="7" place="7" resultid="1651" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1951" daytime="17:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1952" daytime="17:44" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1302" daytime="17:46" gender="F" number="51" order="28" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1303" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1369" />
                    <RANKING order="2" place="2" resultid="1556" />
                    <RANKING order="3" place="3" resultid="1477" />
                    <RANKING order="4" place="4" resultid="1970" />
                    <RANKING order="5" place="5" resultid="1803" />
                    <RANKING order="6" place="6" resultid="1358" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1304" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1346" />
                    <RANKING order="2" place="2" resultid="1340" />
                    <RANKING order="3" place="3" resultid="1535" />
                    <RANKING order="4" place="4" resultid="1687" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1305" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1306" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1328" />
                    <RANKING order="2" place="-1" resultid="1448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1307" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1334" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1308" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1416" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1309" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1953" daytime="17:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1954" daytime="17:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1955" daytime="17:50" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1310" daytime="17:52" gender="M" number="52" order="29" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1311" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1739" />
                    <RANKING order="2" place="2" resultid="1464" />
                    <RANKING order="3" place="3" resultid="1406" />
                    <RANKING order="4" place="4" resultid="1763" />
                    <RANKING order="5" place="5" resultid="1352" />
                    <RANKING order="6" place="6" resultid="1855" />
                    <RANKING order="7" place="7" resultid="1849" />
                    <RANKING order="8" place="-1" resultid="1788" />
                    <RANKING order="9" place="-1" resultid="1798" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1312" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1713" />
                    <RANKING order="2" place="-1" resultid="1585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1313" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1383" />
                    <RANKING order="2" place="2" resultid="1443" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1314" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1393" />
                    <RANKING order="2" place="2" resultid="1439" />
                    <RANKING order="3" place="3" resultid="1401" />
                    <RANKING order="4" place="4" resultid="1560" />
                    <RANKING order="5" place="5" resultid="1693" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1315" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1322" />
                    <RANKING order="2" place="2" resultid="1660" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1316" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1453" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1317" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1412" />
                    <RANKING order="2" place="2" resultid="1682" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1956" daytime="17:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1957" daytime="17:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1958" daytime="17:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="1959" daytime="17:58" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="2864" nation="BRA" region="PR" clubid="1365" swrid="93756" name="Associacao De Pais E Amigos Da Natacao De Ponta Gr" shortname="Apan Ponta Grossa">
          <ATHLETES>
            <ATHLETE firstname="Sofia" lastname="Pontes Mattioli" birthdate="2011-09-10" gender="F" nation="BRA" license="366914" swrid="5602572" athleteid="1366" externalid="366914">
              <RESULTS>
                <RESULT eventid="1132" points="294" swimtime="00:00:37.97" resultid="1367" heatid="1897" lane="2" entrytime="00:00:38.94" entrycourse="SCM" />
                <RESULT eventid="1066" points="290" swimtime="00:03:03.97" resultid="1368" heatid="1875" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:01:24.60" />
                    <SPLIT distance="150" swimtime="00:02:23.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="328" swimtime="00:00:33.22" resultid="1369" heatid="1954" lane="6" entrytime="00:00:34.75" entrycourse="SCM" />
                <RESULT eventid="1280" points="270" swimtime="00:01:24.89" resultid="1370" heatid="1945" lane="3" entrytime="00:01:25.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="241" swimtime="00:00:39.15" resultid="1371" heatid="1935" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2416" nation="BRA" region="PR" clubid="1372" swrid="93758" name="Apan/Maringá">
          <ATHLETES>
            <ATHLETE firstname="Sarah" lastname="Chaim" birthdate="2011-05-29" gender="F" nation="BRA" license="370662" swrid="5409721" athleteid="1474" externalid="370662">
              <RESULTS>
                <RESULT eventid="1132" points="179" swimtime="00:00:44.75" resultid="1475" heatid="1897" lane="1" entrytime="00:00:43.17" entrycourse="SCM" />
                <RESULT eventid="1088" points="245" swimtime="00:01:20.24" resultid="1476" heatid="1882" lane="1" entrytime="00:01:19.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="274" swimtime="00:00:35.27" resultid="1477" heatid="1954" lane="1" entrytime="00:00:34.71" entrycourse="SCM" />
                <RESULT eventid="1254" points="184" swimtime="00:00:42.81" resultid="1478" heatid="1936" lane="5" entrytime="00:00:45.09" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laion" lastname="Miguel Simoes" birthdate="2016-04-02" gender="M" nation="BRA" license="407179" athleteid="1639" externalid="407179">
              <RESULTS>
                <RESULT eventid="1272" points="33" swimtime="00:00:28.13" resultid="1640" heatid="1940" lane="3" />
                <RESULT eventid="1246" points="27" swimtime="00:00:37.92" resultid="1641" heatid="1931" lane="3" />
                <RESULT eventid="1220" points="29" swimtime="00:00:33.37" resultid="1642" heatid="1925" lane="3" />
                <RESULT eventid="1194" points="19" swimtime="00:00:36.50" resultid="1643" heatid="1917" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Bessa" birthdate="2003-06-19" gender="M" nation="BRA" license="317841" swrid="5312237" athleteid="1377" externalid="317841">
              <RESULTS>
                <RESULT eventid="1184" points="588" swimtime="00:00:29.77" resultid="1378" heatid="1916" lane="3" entrytime="00:00:29.02" entrycourse="SCM" />
                <RESULT eventid="1074" status="DSQ" swimtime="00:02:24.50" resultid="1379" heatid="1876" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                    <SPLIT distance="150" swimtime="00:01:45.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="624" swimtime="00:01:04.67" resultid="1380" heatid="1930" lane="3" entrytime="00:01:03.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Marques" birthdate="2015-10-15" gender="F" nation="BRA" license="399738" swrid="5651346" athleteid="1611" externalid="399738">
              <RESULTS>
                <RESULT eventid="1296" points="21" swimtime="00:01:22.02" resultid="1612" heatid="1949" lane="3" />
                <RESULT eventid="1248" points="38" swimtime="00:01:15.08" resultid="1613" heatid="1932" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Pacheco" birthdate="2006-12-20" gender="M" nation="BRA" license="336850" swrid="5603854" athleteid="1423" externalid="336850">
              <RESULTS>
                <RESULT eventid="1162" points="446" swimtime="00:01:02.53" resultid="1424" heatid="1908" lane="2" entrytime="00:01:02.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1262" points="438" swimtime="00:00:28.63" resultid="1425" heatid="1937" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Vitoria Moreira Ferreira" birthdate="2012-08-04" gender="F" nation="BRA" license="392098" swrid="5603928" athleteid="1549" externalid="392098">
              <RESULTS>
                <RESULT eventid="1148" points="144" swimtime="00:01:47.70" resultid="1550" heatid="1900" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="125" swimtime="00:00:50.38" resultid="1551" heatid="1887" lane="4" />
                <RESULT eventid="1082" points="131" swimtime="00:02:02.48" resultid="1552" heatid="1880" lane="5" entrytime="00:02:11.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Peroni Passafaro" birthdate="2013-09-17" gender="F" nation="BRA" license="370659" swrid="5603893" athleteid="1470" externalid="370659">
              <RESULTS>
                <RESULT eventid="1148" points="163" swimtime="00:01:43.33" resultid="1471" heatid="1902" lane="6" entrytime="00:01:51.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="174" swimtime="00:00:45.15" resultid="1472" heatid="1889" lane="1" entrytime="00:00:45.82" entrycourse="SCM" />
                <RESULT eventid="1060" points="203" swimtime="00:03:07.52" resultid="1473" heatid="1872" lane="6" entrytime="00:03:31.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                    <SPLIT distance="100" swimtime="00:01:31.66" />
                    <SPLIT distance="150" swimtime="00:02:20.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Hugo Santos" birthdate="2007-03-26" gender="M" nation="BRA" license="384355" swrid="5603855" athleteid="1523" externalid="384355">
              <RESULTS>
                <RESULT eventid="1140" status="DNS" swimtime="00:00:00.00" resultid="1524" heatid="1899" lane="6" entrytime="00:00:38.94" entrycourse="SCM" />
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="1525" heatid="1885" lane="5" entrytime="00:01:08.85" entrycourse="SCM" />
                <RESULT eventid="1210" status="DNS" swimtime="00:00:00.00" resultid="1526" heatid="1923" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Garcia Cavalcante" birthdate="2011-11-21" gender="M" nation="BRA" license="378200" swrid="5603840" athleteid="1403" externalid="378200">
              <RESULTS>
                <RESULT eventid="1184" points="222" swimtime="00:00:41.15" resultid="1404" heatid="1915" lane="3" entrytime="00:00:42.20" entrycourse="SCM" />
                <RESULT eventid="1074" points="221" swimtime="00:03:01.19" resultid="1405" heatid="1877" lane="5" entrytime="00:03:09.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.05" />
                    <SPLIT distance="100" swimtime="00:01:30.82" />
                    <SPLIT distance="150" swimtime="00:02:21.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="234" swimtime="00:00:32.70" resultid="1406" heatid="1957" lane="4" entrytime="00:00:33.60" entrycourse="SCM" />
                <RESULT eventid="1236" points="222" swimtime="00:01:31.29" resultid="1407" heatid="1929" lane="2" entrytime="00:01:35.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Casavechia Carraro" birthdate="2009-07-28" gender="M" nation="BRA" license="368150" swrid="5384752" athleteid="1381" externalid="368150">
              <RESULTS>
                <RESULT eventid="1162" points="491" swimtime="00:01:00.55" resultid="1382" heatid="1908" lane="4" entrytime="00:01:00.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="503" swimtime="00:00:25.34" resultid="1383" heatid="1959" lane="4" entrytime="00:00:24.99" entrycourse="SCM" />
                <RESULT eventid="1210" points="514" swimtime="00:04:24.87" resultid="1384" heatid="1924" lane="4" entrytime="00:04:29.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                    <SPLIT distance="100" swimtime="00:01:03.25" />
                    <SPLIT distance="150" swimtime="00:01:36.90" />
                    <SPLIT distance="200" swimtime="00:02:09.97" />
                    <SPLIT distance="250" swimtime="00:02:43.39" />
                    <SPLIT distance="300" swimtime="00:03:17.07" />
                    <SPLIT distance="350" swimtime="00:03:50.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Altoé" birthdate="2003-01-29" gender="M" nation="BRA" license="251546" swrid="5616194" athleteid="1408" externalid="251546">
              <RESULTS>
                <RESULT eventid="1184" status="DSQ" swimtime="00:00:24.11" resultid="1409" heatid="1915" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Coleto Arcanjo" birthdate="2015-08-17" gender="F" nation="BRA" license="407176" athleteid="1632" externalid="407176">
              <RESULTS>
                <RESULT eventid="1296" points="38" swimtime="00:01:07.66" resultid="1633" heatid="1950" lane="6" />
                <RESULT eventid="1248" points="40" swimtime="00:01:13.77" resultid="1634" heatid="1932" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Forti Francisco" birthdate="2015-07-08" gender="M" nation="BRA" license="392104" swrid="5534395" athleteid="1562" externalid="392104">
              <RESULTS>
                <RESULT eventid="1277" points="70" swimtime="00:01:00.48" resultid="1563" heatid="1944" lane="1" />
                <RESULT eventid="1225" points="54" swimtime="00:00:57.51" resultid="1564" heatid="1927" lane="1" />
                <RESULT eventid="1199" points="66" swimtime="00:01:50.67" resultid="1565" heatid="1920" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wellington" lastname="De Lima" birthdate="2008-03-01" gender="M" nation="BRA" license="370024" swrid="5470912" athleteid="1390" externalid="370024">
              <RESULTS>
                <RESULT eventid="1140" points="388" swimtime="00:00:30.29" resultid="1391" heatid="1898" lane="4" />
                <RESULT eventid="1096" points="495" swimtime="00:00:56.67" resultid="1392" heatid="1886" lane="2" entrytime="00:00:56.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="434" swimtime="00:00:26.62" resultid="1393" heatid="1959" lane="2" entrytime="00:00:26.36" entrycourse="SCM" />
                <RESULT eventid="1288" points="325" swimtime="00:01:10.23" resultid="1394" heatid="1948" lane="2" entrytime="00:01:07.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Antônio Boeing" birthdate="2004-06-04" gender="M" nation="BRA" license="317474" swrid="5184340" athleteid="1410" externalid="317474">
              <RESULTS>
                <RESULT eventid="1140" points="574" swimtime="00:00:26.59" resultid="1411" heatid="1899" lane="3" entrytime="00:00:25.65" entrycourse="SCM" />
                <RESULT eventid="1310" points="629" swimtime="00:00:23.52" resultid="1412" heatid="1959" lane="3" entrytime="00:00:24.15" entrycourse="SCM" />
                <RESULT eventid="1262" points="627" swimtime="00:00:25.41" resultid="1413" heatid="1938" lane="3" entrytime="00:00:24.01" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Pacheco" birthdate="2012-10-03" gender="M" nation="BRA" license="370663" swrid="5603883" athleteid="1479" externalid="370663">
              <RESULTS>
                <RESULT eventid="1173" points="225" swimtime="00:00:33.12" resultid="1480" heatid="1913" lane="2" entrytime="00:00:33.58" entrycourse="SCM" />
                <RESULT eventid="1151" points="174" swimtime="00:01:28.19" resultid="1481" heatid="1903" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="154" swimtime="00:00:41.22" resultid="1482" heatid="1890" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Furuchi Martins" birthdate="2011-10-05" gender="F" nation="BRA" license="367001" swrid="5602616" athleteid="1964" externalid="367001">
              <RESULTS>
                <RESULT eventid="1066" points="216" swimtime="00:03:23.01" resultid="1965" heatid="1875" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.13" />
                    <SPLIT distance="100" swimtime="00:01:41.68" />
                    <SPLIT distance="150" swimtime="00:02:38.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="273" swimtime="00:00:43.69" resultid="1967" heatid="1966" lane="3" late="yes" />
                <RESULT eventid="1302" points="238" swimtime="00:00:36.99" resultid="1970" heatid="1953" lane="2" late="yes" />
                <RESULT eventid="1228" points="270" swimtime="00:01:36.47" resultid="1974" heatid="1928" lane="2" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Otavio Luz" birthdate="2013-07-27" gender="M" nation="BRA" license="392111" swrid="5603882" athleteid="1578" externalid="392111">
              <RESULTS>
                <RESULT eventid="1173" points="160" swimtime="00:00:37.09" resultid="1579" heatid="1913" lane="6" entrytime="00:00:36.95" entrycourse="SCM" />
                <RESULT eventid="1129" status="DSQ" swimtime="00:01:42.43" resultid="1580" heatid="1896" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="118" swimtime="00:00:45.05" resultid="1581" heatid="1890" lane="3" entrytime="00:00:51.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Muniz" birthdate="2012-09-03" gender="M" nation="BRA" license="392106" swrid="5603877" athleteid="1566" externalid="392106">
              <RESULTS>
                <RESULT eventid="1173" points="118" swimtime="00:00:41.10" resultid="1567" heatid="1912" lane="5" entrytime="00:00:40.27" entrycourse="SCM" />
                <RESULT eventid="1151" points="86" swimtime="00:01:51.34" resultid="1568" heatid="1903" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="73" swimtime="00:00:52.84" resultid="1569" heatid="1890" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Donato De Morais" birthdate="2009-03-28" gender="F" nation="BRA" license="345588" swrid="5485198" athleteid="1426" externalid="345588">
              <RESULTS>
                <RESULT eventid="1088" points="343" swimtime="00:01:11.77" resultid="1427" heatid="1883" lane="6" entrytime="00:01:10.41" entrycourse="SCM" />
                <RESULT eventid="1280" points="337" swimtime="00:01:18.80" resultid="1428" heatid="1946" lane="2" entrytime="00:01:16.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="347" swimtime="00:05:28.96" resultid="1429" heatid="1922" lane="2" entrytime="00:05:22.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                    <SPLIT distance="100" swimtime="00:01:18.06" />
                    <SPLIT distance="150" swimtime="00:02:00.30" />
                    <SPLIT distance="200" swimtime="00:02:42.09" />
                    <SPLIT distance="250" swimtime="00:03:24.81" />
                    <SPLIT distance="300" swimtime="00:04:06.78" />
                    <SPLIT distance="350" swimtime="00:04:49.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raphael" lastname="Piai Pellegrini" birthdate="2012-03-24" gender="M" nation="BRA" license="377261" swrid="5603894" athleteid="1495" externalid="377261">
              <RESULTS>
                <RESULT eventid="1173" points="275" swimtime="00:00:31.00" resultid="1496" heatid="1913" lane="3" entrytime="00:00:32.16" entrycourse="SCM" />
                <RESULT eventid="1151" points="190" swimtime="00:01:25.60" resultid="1497" heatid="1903" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="263" swimtime="00:02:35.01" resultid="1498" heatid="1874" lane="4" entrytime="00:02:38.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                    <SPLIT distance="100" swimtime="00:01:13.13" />
                    <SPLIT distance="150" swimtime="00:01:54.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Fernandes Rivadavia" birthdate="2015-11-15" gender="F" nation="BRA" license="393774" swrid="5651342" athleteid="1591" externalid="393774">
              <RESULTS>
                <RESULT eventid="1274" points="122" swimtime="00:00:57.20" resultid="1592" heatid="1942" lane="5" />
                <RESULT eventid="1222" points="95" swimtime="00:00:53.26" resultid="1593" heatid="1926" lane="1" />
                <RESULT eventid="1196" points="152" swimtime="00:01:34.01" resultid="1594" heatid="1918" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Martins Pedro" birthdate="2015-01-19" gender="F" nation="BRA" license="403390" swrid="5676290" athleteid="1621" externalid="403390">
              <RESULTS>
                <RESULT eventid="1222" points="37" swimtime="00:01:12.55" resultid="1622" heatid="1926" lane="4" />
                <RESULT eventid="1196" points="71" swimtime="00:02:01.07" resultid="1623" heatid="1918" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Camila Cuenca" birthdate="2005-10-06" gender="F" nation="BRA" license="308081" swrid="5357445" athleteid="1414" externalid="308081">
              <RESULTS>
                <RESULT eventid="1088" points="426" swimtime="00:01:06.78" resultid="1415" heatid="1883" lane="4" entrytime="00:01:03.20" entrycourse="SCM" />
                <RESULT eventid="1302" points="429" swimtime="00:00:30.38" resultid="1416" heatid="1955" lane="3" entrytime="00:00:28.93" entrycourse="SCM" />
                <RESULT eventid="1280" points="374" swimtime="00:01:16.14" resultid="1417" heatid="1945" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="438" swimtime="00:05:04.53" resultid="1418" heatid="1921" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                    <SPLIT distance="100" swimtime="00:01:13.56" />
                    <SPLIT distance="150" swimtime="00:01:52.17" />
                    <SPLIT distance="200" swimtime="00:02:31.36" />
                    <SPLIT distance="250" swimtime="00:03:10.06" />
                    <SPLIT distance="300" swimtime="00:03:49.03" />
                    <SPLIT distance="350" swimtime="00:04:27.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Marques Picolo Vinha" birthdate="2010-07-01" gender="M" nation="BRA" license="366990" swrid="5603869" athleteid="1582" externalid="366990">
              <RESULTS>
                <RESULT eventid="1184" status="DNS" swimtime="00:00:00.00" resultid="1583" heatid="1915" lane="4" />
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="1584" heatid="1885" lane="4" entrytime="00:01:05.40" entrycourse="SCM" />
                <RESULT eventid="1310" status="DNS" swimtime="00:00:00.00" resultid="1585" heatid="1958" lane="3" entrytime="00:00:29.57" entrycourse="SCM" />
                <RESULT eventid="1210" status="DNS" swimtime="00:00:00.00" resultid="1586" heatid="1923" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Constantino" birthdate="2012-06-02" gender="F" nation="BRA" license="382208" swrid="5420069" athleteid="1511" externalid="382208">
              <RESULTS>
                <RESULT eventid="1170" points="257" swimtime="00:00:36.06" resultid="1512" heatid="1911" lane="2" entrytime="00:00:35.62" entrycourse="SCM" />
                <RESULT eventid="1104" points="172" swimtime="00:00:45.37" resultid="1513" heatid="1889" lane="5" entrytime="00:00:45.63" entrycourse="SCM" />
                <RESULT eventid="1082" points="237" swimtime="00:01:40.72" resultid="1514" heatid="1880" lane="2" entrytime="00:01:46.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Passafaro" birthdate="2009-02-01" gender="F" nation="BRA" license="370673" swrid="5603885" athleteid="1430" externalid="370673">
              <RESULTS>
                <RESULT eventid="1132" points="251" swimtime="00:00:40.02" resultid="1431" heatid="1897" lane="5" entrytime="00:00:40.89" entrycourse="SCM" />
                <RESULT eventid="1088" points="310" swimtime="00:01:14.19" resultid="1432" heatid="1883" lane="1" entrytime="00:01:09.23" entrycourse="SCM" />
                <RESULT eventid="1302" points="344" swimtime="00:00:32.72" resultid="1433" heatid="1955" lane="1" entrytime="00:00:30.79" entrycourse="SCM" />
                <RESULT eventid="1254" points="346" swimtime="00:00:34.72" resultid="1434" heatid="1936" lane="4" entrytime="00:00:34.84" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicole" lastname="De Meira" birthdate="2012-01-21" gender="F" nation="BRA" license="377257" swrid="5615583" athleteid="1483" externalid="377257">
              <RESULTS>
                <RESULT eventid="1170" points="117" swimtime="00:00:46.75" resultid="1484" heatid="1909" lane="2" entrytime="00:00:47.89" entrycourse="SCM" />
                <RESULT eventid="1104" points="83" swimtime="00:00:57.72" resultid="1485" heatid="1887" lane="3" />
                <RESULT eventid="1082" points="108" swimtime="00:02:10.94" resultid="1486" heatid="1880" lane="1" entrytime="00:02:22.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Beatriz Meira" birthdate="2012-04-11" gender="F" nation="BRA" license="392094" swrid="5305414" athleteid="1537" externalid="392094">
              <RESULTS>
                <RESULT eventid="1170" points="160" swimtime="00:00:42.21" resultid="1538" heatid="1909" lane="4" entrytime="00:00:45.90" entrycourse="SCM" />
                <RESULT eventid="1148" points="102" swimtime="00:02:00.90" resultid="1539" heatid="1900" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="116" swimtime="00:00:51.68" resultid="1540" heatid="1888" lane="1" entrytime="00:01:10.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Corsine Ferreira" birthdate="2010-03-10" gender="F" nation="BRA" license="353591" swrid="5588608" athleteid="1527" externalid="353591">
              <RESULTS>
                <RESULT eventid="1110" points="294" swimtime="00:22:45.06" resultid="1528" heatid="1892" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="360" swimtime="00:02:51.26" resultid="1529" heatid="1960" lane="4" entrytime="00:02:53.30" entrycourse="SCM" />
                <RESULT eventid="1280" points="374" swimtime="00:01:16.12" resultid="1530" heatid="1946" lane="3" entrytime="00:01:13.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="301" swimtime="00:01:33.00" resultid="1531" heatid="1928" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Allyce" lastname="Rodrigues Tavares" birthdate="2014-10-13" gender="F" nation="BRA" license="403389" swrid="5676291" athleteid="1618" externalid="403389">
              <RESULTS>
                <RESULT eventid="1296" points="17" swimtime="00:01:27.50" resultid="1619" heatid="1949" lane="5" />
                <RESULT eventid="1248" points="34" swimtime="00:01:17.76" resultid="1620" heatid="1932" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Yukio Tacaiama" birthdate="2014-06-29" gender="M" nation="BRA" license="407184" athleteid="1653" externalid="407184">
              <RESULTS>
                <RESULT eventid="1299" points="97" swimtime="00:00:43.78" resultid="1654" heatid="1951" lane="3" />
                <RESULT eventid="1277" points="78" swimtime="00:00:58.37" resultid="1655" heatid="1944" lane="5" />
                <RESULT eventid="1199" points="99" swimtime="00:01:36.82" resultid="1656" heatid="1919" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heitor" lastname="Bello Paula" birthdate="2015-06-14" gender="M" nation="BRA" license="393776" swrid="5507529" athleteid="1595" externalid="393776">
              <RESULTS>
                <RESULT eventid="1299" points="89" swimtime="00:00:45.12" resultid="1596" heatid="1952" lane="6" entrytime="00:00:58.94" entrycourse="SCM" />
                <RESULT eventid="1251" points="61" swimtime="00:00:56.00" resultid="1597" heatid="1934" lane="6" />
                <RESULT eventid="1225" points="41" swimtime="00:01:02.80" resultid="1598" heatid="1927" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Campos" birthdate="2013-02-17" gender="M" nation="BRA" license="377262" swrid="5641756" athleteid="1499" externalid="377262">
              <RESULTS>
                <RESULT eventid="1151" points="146" swimtime="00:01:33.51" resultid="1500" heatid="1904" lane="3" entrytime="00:01:39.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="146" swimtime="00:00:41.97" resultid="1501" heatid="1891" lane="4" entrytime="00:00:38.73" entrycourse="SCM" />
                <RESULT eventid="1063" points="171" swimtime="00:02:59.02" resultid="1502" heatid="1874" lane="5" entrytime="00:02:56.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:01:26.29" />
                    <SPLIT distance="150" swimtime="00:02:13.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Arthur Da Silva Ortiz" birthdate="2015-04-20" gender="M" nation="BRA" license="399733" swrid="5676285" athleteid="1603" externalid="399733">
              <RESULTS>
                <RESULT eventid="1299" points="79" swimtime="00:00:46.87" resultid="1604" heatid="1951" lane="1" />
                <RESULT eventid="1277" points="86" swimtime="00:00:56.36" resultid="1605" heatid="1943" lane="4" />
                <RESULT eventid="1225" points="57" swimtime="00:00:56.35" resultid="1606" heatid="1927" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Sol Reolon Gomes" birthdate="2011-02-28" gender="F" nation="BRA" license="392100" swrid="5603914" athleteid="1553" externalid="392100">
              <RESULTS>
                <RESULT eventid="1132" points="267" swimtime="00:00:39.18" resultid="1554" heatid="1897" lane="4" entrytime="00:00:38.80" entrycourse="SCM" />
                <RESULT eventid="1066" points="247" swimtime="00:03:14.08" resultid="1555" heatid="1960" lane="5" entrytime="00:03:22.24" entrycourse="SCM" />
                <RESULT eventid="1302" points="324" swimtime="00:00:33.36" resultid="1556" heatid="1954" lane="2" entrytime="00:00:33.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Dos Reis Monteiro" birthdate="2014-08-05" gender="M" nation="BRA" license="392095" swrid="5697226" athleteid="1541" externalid="392095">
              <RESULTS>
                <RESULT eventid="1277" points="167" swimtime="00:00:45.28" resultid="1542" heatid="1944" lane="3" entrytime="00:00:43.78" entrycourse="SCM" />
                <RESULT eventid="1251" points="111" swimtime="00:00:45.97" resultid="1543" heatid="1934" lane="2" />
                <RESULT eventid="1199" points="205" swimtime="00:01:15.98" resultid="1544" heatid="1920" lane="3" entrytime="00:01:18.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Rampasi" birthdate="2013-10-16" gender="F" nation="BRA" license="382209" swrid="5603866" athleteid="1515" externalid="382209">
              <RESULTS>
                <RESULT eventid="1170" points="160" swimtime="00:00:42.16" resultid="1516" heatid="1910" lane="5" entrytime="00:00:43.13" entrycourse="SCM" />
                <RESULT eventid="1126" points="92" swimtime="00:01:59.47" resultid="1517" heatid="1894" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="158" swimtime="00:03:23.64" resultid="1518" heatid="1871" lane="3" entrytime="00:03:36.58" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Izzo Breschiliare" birthdate="2015-09-23" gender="M" nation="BRA" license="407182" athleteid="1647" externalid="407182">
              <RESULTS>
                <RESULT eventid="1299" points="37" swimtime="00:01:00.12" resultid="1648" heatid="1951" lane="4" />
                <RESULT eventid="1251" points="39" swimtime="00:01:04.74" resultid="1649" heatid="1934" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Ficher Delmont Pais" birthdate="2010-07-15" gender="M" nation="BRA" license="338533" swrid="5588701" athleteid="1385" externalid="338533">
              <RESULTS>
                <RESULT eventid="1118" points="346" swimtime="00:20:05.61" resultid="1386" heatid="1893" lane="3" />
                <RESULT eventid="1074" points="426" swimtime="00:02:25.66" resultid="1387" heatid="1878" lane="3" entrytime="00:02:23.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                    <SPLIT distance="100" swimtime="00:01:07.08" />
                    <SPLIT distance="150" swimtime="00:01:51.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="366" swimtime="00:01:07.53" resultid="1388" heatid="1948" lane="4" entrytime="00:01:04.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1210" points="408" swimtime="00:04:45.98" resultid="1389" heatid="1924" lane="2" entrytime="00:04:51.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                    <SPLIT distance="100" swimtime="00:01:06.29" />
                    <SPLIT distance="150" swimtime="00:01:42.21" />
                    <SPLIT distance="200" swimtime="00:02:18.92" />
                    <SPLIT distance="250" swimtime="00:02:56.65" />
                    <SPLIT distance="300" swimtime="00:03:33.60" />
                    <SPLIT distance="350" swimtime="00:04:09.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Batista Sanchez" birthdate="2009-05-22" gender="M" nation="BRA" license="370668" swrid="5255779" athleteid="1395" externalid="370668">
              <RESULTS>
                <RESULT eventid="1184" points="332" swimtime="00:00:36.01" resultid="1396" heatid="1916" lane="2" entrytime="00:00:36.89" entrycourse="SCM" />
                <RESULT eventid="1262" points="245" swimtime="00:00:34.73" resultid="1397" heatid="1938" lane="1" entrytime="00:00:33.23" entrycourse="SCM" />
                <RESULT eventid="1236" points="381" swimtime="00:01:16.25" resultid="1398" heatid="1930" lane="6" entrytime="00:01:18.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Sossai Altoe" birthdate="2006-09-04" gender="M" nation="BRA" license="296488" swrid="5603915" athleteid="1373" externalid="296488">
              <RESULTS>
                <RESULT eventid="1096" points="564" swimtime="00:00:54.25" resultid="1374" heatid="1886" lane="3" entrytime="00:00:52.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1262" points="485" swimtime="00:00:27.68" resultid="1375" heatid="1938" lane="4" entrytime="00:00:26.82" entrycourse="SCM" />
                <RESULT eventid="1210" points="544" swimtime="00:04:19.95" resultid="1376" heatid="1924" lane="3" entrytime="00:04:18.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                    <SPLIT distance="100" swimtime="00:01:01.31" />
                    <SPLIT distance="150" swimtime="00:01:35.12" />
                    <SPLIT distance="200" swimtime="00:02:09.40" />
                    <SPLIT distance="250" swimtime="00:02:41.59" />
                    <SPLIT distance="300" swimtime="00:03:14.20" />
                    <SPLIT distance="350" swimtime="00:03:47.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Reolon Gomes" birthdate="2014-06-21" gender="M" nation="BRA" license="407183" athleteid="1650" externalid="407183">
              <RESULTS>
                <RESULT eventid="1299" points="45" swimtime="00:00:56.36" resultid="1651" heatid="1951" lane="5" />
                <RESULT eventid="1251" points="37" swimtime="00:01:05.85" resultid="1652" heatid="1934" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Quental De Meireles" birthdate="2008-11-20" gender="M" nation="BRA" license="392103" swrid="5603898" athleteid="1557" externalid="392103">
              <RESULTS>
                <RESULT eventid="1096" points="339" swimtime="00:01:04.27" resultid="1558" heatid="1885" lane="6" entrytime="00:01:10.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="318" swimtime="00:02:40.58" resultid="1559" heatid="1876" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:16.82" />
                    <SPLIT distance="150" swimtime="00:02:03.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="324" swimtime="00:00:29.34" resultid="1560" heatid="1958" lane="5" entrytime="00:00:30.35" entrycourse="SCM" />
                <RESULT eventid="1236" points="319" swimtime="00:01:20.84" resultid="1561" heatid="1929" lane="4" entrytime="00:01:26.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Bassil" birthdate="2015-07-02" gender="M" nation="BRA" license="407178" athleteid="1635" externalid="407178">
              <RESULTS>
                <RESULT eventid="1299" points="69" swimtime="00:00:49.14" resultid="1636" heatid="1951" lane="6" />
                <RESULT eventid="1277" points="74" swimtime="00:00:59.32" resultid="1637" heatid="1943" lane="3" />
                <RESULT eventid="1199" points="72" swimtime="00:01:47.33" resultid="1638" heatid="1919" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Paiva Boeing" birthdate="2008-01-22" gender="F" nation="BRA" license="318185" swrid="5603884" athleteid="1419" externalid="318185">
              <RESULTS>
                <RESULT eventid="1154" points="332" swimtime="00:01:17.98" resultid="1420" heatid="1905" lane="3" />
                <RESULT eventid="1254" points="377" swimtime="00:00:33.73" resultid="1421" heatid="1936" lane="3" entrytime="00:00:33.46" entrycourse="SCM" />
                <RESULT eventid="1202" points="370" swimtime="00:05:21.99" resultid="1422" heatid="1921" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                    <SPLIT distance="100" swimtime="00:01:16.23" />
                    <SPLIT distance="150" swimtime="00:01:58.17" />
                    <SPLIT distance="200" swimtime="00:02:40.18" />
                    <SPLIT distance="250" swimtime="00:03:20.97" />
                    <SPLIT distance="300" swimtime="00:04:02.87" />
                    <SPLIT distance="350" swimtime="00:04:43.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mochiutti Carneiro" birthdate="2010-04-22" gender="F" nation="BRA" license="370670" swrid="5588817" athleteid="1532" externalid="370670">
              <RESULTS>
                <RESULT eventid="1154" points="341" swimtime="00:01:17.34" resultid="1533" heatid="1906" lane="3" entrytime="00:01:16.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="451" swimtime="00:01:05.48" resultid="1534" heatid="1883" lane="2" entrytime="00:01:06.28" entrycourse="SCM" />
                <RESULT eventid="1302" points="427" swimtime="00:00:30.44" resultid="1535" heatid="1955" lane="2" entrytime="00:00:30.51" entrycourse="SCM" />
                <RESULT eventid="1202" points="408" swimtime="00:05:11.84" resultid="1536" heatid="1922" lane="5" entrytime="00:05:23.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.36" />
                    <SPLIT distance="100" swimtime="00:01:15.05" />
                    <SPLIT distance="150" swimtime="00:01:55.42" />
                    <SPLIT distance="200" swimtime="00:02:35.04" />
                    <SPLIT distance="250" swimtime="00:03:14.58" />
                    <SPLIT distance="300" swimtime="00:03:54.48" />
                    <SPLIT distance="350" swimtime="00:04:33.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Pastre" birthdate="2014-03-10" gender="F" nation="BRA" license="403760" swrid="5684593" athleteid="1624" externalid="403760">
              <RESULTS>
                <RESULT eventid="1296" points="117" swimtime="00:00:46.81" resultid="1625" heatid="1950" lane="5" entrytime="00:00:49.24" entrycourse="SCM" />
                <RESULT eventid="1248" points="144" swimtime="00:00:48.08" resultid="1626" heatid="1933" lane="3" entrytime="00:00:53.06" entrycourse="SCM" />
                <RESULT eventid="1196" points="104" swimtime="00:01:46.80" resultid="1627" heatid="1918" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Antonio Mendes" birthdate="2008-12-04" gender="M" nation="BRA" license="366962" swrid="5196287" athleteid="1435" externalid="366962">
              <RESULTS>
                <RESULT eventid="1184" points="488" swimtime="00:00:31.69" resultid="1436" heatid="1916" lane="4" entrytime="00:00:33.27" entrycourse="SCM" />
                <RESULT eventid="1140" points="392" swimtime="00:00:30.20" resultid="1437" heatid="1899" lane="4" entrytime="00:00:31.26" entrycourse="SCM" />
                <RESULT eventid="1074" points="428" swimtime="00:02:25.40" resultid="1438" heatid="1876" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:07.84" />
                    <SPLIT distance="150" swimtime="00:01:48.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="418" swimtime="00:00:26.95" resultid="1439" heatid="1956" lane="3" />
                <RESULT eventid="1288" points="395" swimtime="00:01:05.85" resultid="1440" heatid="1948" lane="5" entrytime="00:01:08.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mendes Costa" birthdate="2014-04-03" gender="F" nation="BRA" license="378341" swrid="5603873" athleteid="1628" externalid="378341">
              <RESULTS>
                <RESULT eventid="1296" points="128" swimtime="00:00:45.47" resultid="1629" heatid="1950" lane="2" entrytime="00:00:47.55" entrycourse="SCM" />
                <RESULT eventid="1274" points="115" swimtime="00:00:58.27" resultid="1630" heatid="1942" lane="2" entrytime="00:01:03.04" entrycourse="SCM" />
                <RESULT eventid="1222" points="82" swimtime="00:00:56.06" resultid="1631" heatid="1926" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Bernardo Padua" birthdate="2013-07-15" gender="M" nation="BRA" license="392108" swrid="5305422" athleteid="1570" externalid="392108">
              <RESULTS>
                <RESULT eventid="1173" points="130" swimtime="00:00:39.76" resultid="1571" heatid="1912" lane="2" entrytime="00:00:39.45" entrycourse="SCM" />
                <RESULT eventid="1151" points="132" swimtime="00:01:36.60" resultid="1572" heatid="1904" lane="4" entrytime="00:01:48.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="144" swimtime="00:01:45.31" resultid="1573" heatid="1881" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Biason Santana" birthdate="2009-01-21" gender="M" nation="BRA" license="366969" swrid="5317765" athleteid="1441" externalid="366969">
              <RESULTS>
                <RESULT eventid="1162" points="390" swimtime="00:01:05.36" resultid="1442" heatid="1908" lane="1" entrytime="00:01:04.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="394" swimtime="00:00:27.49" resultid="1443" heatid="1959" lane="6" entrytime="00:00:28.15" entrycourse="SCM" />
                <RESULT eventid="1262" points="416" swimtime="00:00:29.12" resultid="1444" heatid="1938" lane="2" entrytime="00:00:29.07" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Pavão" birthdate="2012-04-04" gender="F" nation="BRA" license="377259" swrid="5603888" athleteid="1487" externalid="377259">
              <RESULTS>
                <RESULT eventid="1148" points="212" swimtime="00:01:34.70" resultid="1488" heatid="1901" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="191" swimtime="00:00:43.82" resultid="1489" heatid="1889" lane="4" entrytime="00:00:44.30" entrycourse="SCM" />
                <RESULT eventid="1060" points="181" swimtime="00:03:14.72" resultid="1490" heatid="1871" lane="4" entrytime="00:03:39.26" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauan" lastname="Gabriel Pereira" birthdate="2014-05-14" gender="M" nation="BRA" license="407181" athleteid="1644" externalid="407181">
              <RESULTS>
                <RESULT eventid="1299" points="58" swimtime="00:00:52.03" resultid="1645" heatid="1951" lane="2" />
                <RESULT eventid="1251" points="39" swimtime="00:01:05.08" resultid="1646" heatid="1934" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Campelo" birthdate="2011-09-12" gender="M" nation="BRA" license="366963" swrid="5588742" athleteid="1457" externalid="366963">
              <RESULTS>
                <RESULT eventid="1162" points="260" swimtime="00:01:14.85" resultid="1458" heatid="1907" lane="3" entrytime="00:01:22.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="350" swimtime="00:01:03.59" resultid="1459" heatid="1885" lane="3" entrytime="00:01:04.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="280" swimtime="00:01:13.87" resultid="1460" heatid="1948" lane="6" entrytime="00:01:16.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Tomazeli" birthdate="2013-02-05" gender="M" nation="BRA" license="392109" swrid="5614097" athleteid="1574" externalid="392109">
              <RESULTS>
                <RESULT eventid="1151" points="133" swimtime="00:01:36.37" resultid="1575" heatid="1904" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="126" swimtime="00:00:44.00" resultid="1576" heatid="1891" lane="5" entrytime="00:00:45.72" entrycourse="SCM" />
                <RESULT eventid="1063" points="159" swimtime="00:03:03.26" resultid="1577" heatid="1873" lane="2" entrytime="00:03:11.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                    <SPLIT distance="100" swimtime="00:01:25.80" />
                    <SPLIT distance="150" swimtime="00:02:14.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Inoue" birthdate="2008-10-31" gender="F" nation="BRA" license="378348" swrid="5603856" athleteid="1445" externalid="378348">
              <RESULTS>
                <RESULT eventid="1154" points="205" swimtime="00:01:31.65" resultid="1446" heatid="1906" lane="5" entrytime="00:01:25.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="326" swimtime="00:01:12.95" resultid="1447" heatid="1882" lane="5" entrytime="00:01:14.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" status="DSQ" swimtime="00:00:32.61" resultid="1448" heatid="1954" lane="4" entrytime="00:00:32.38" entrycourse="SCM" />
                <RESULT eventid="1202" points="241" swimtime="00:06:11.45" resultid="1449" heatid="1922" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.85" />
                    <SPLIT distance="100" swimtime="00:01:29.06" />
                    <SPLIT distance="150" swimtime="00:02:16.79" />
                    <SPLIT distance="200" swimtime="00:03:05.11" />
                    <SPLIT distance="250" swimtime="00:03:52.54" />
                    <SPLIT distance="300" swimtime="00:04:39.84" />
                    <SPLIT distance="350" swimtime="00:05:27.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Catarina" lastname="Wendt Jesus" birthdate="2013-07-09" gender="F" nation="BRA" license="393778" swrid="5641780" athleteid="1599" externalid="393778">
              <RESULTS>
                <RESULT eventid="1170" points="317" swimtime="00:00:33.62" resultid="1600" heatid="1911" lane="4" entrytime="00:00:35.30" entrycourse="SCM" />
                <RESULT eventid="1126" points="165" swimtime="00:01:38.41" resultid="1601" heatid="1895" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1082" points="278" swimtime="00:01:35.45" resultid="1602" heatid="1879" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Ayres" birthdate="2012-05-05" gender="M" nation="BRA" license="378035" swrid="5208079" athleteid="1503" externalid="378035">
              <RESULTS>
                <RESULT eventid="1151" points="212" swimtime="00:01:22.54" resultid="1504" heatid="1903" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="195" swimtime="00:01:35.24" resultid="1505" heatid="1881" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="286" swimtime="00:02:30.70" resultid="1506" heatid="1874" lane="3" entrytime="00:02:34.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="100" swimtime="00:01:11.40" />
                    <SPLIT distance="150" swimtime="00:01:52.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Danilo" lastname="Seganfredo Boscolo" birthdate="2012-09-15" gender="M" nation="BRA" license="399737" swrid="5651351" athleteid="1607" externalid="399737">
              <RESULTS>
                <RESULT eventid="1173" points="100" swimtime="00:00:43.31" resultid="1608" heatid="1912" lane="1" entrytime="00:00:52.97" entrycourse="SCM" />
                <RESULT eventid="1151" points="85" swimtime="00:01:51.88" resultid="1609" heatid="1904" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="117" swimtime="00:01:52.98" resultid="1610" heatid="1881" lane="4" entrytime="00:02:22.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Furuchi Martins" birthdate="2011-10-05" gender="F" nation="BRA" swrid="5602616" athleteid="1961" />
            <ATHLETE firstname="Rafael" lastname="Felipe Sakaguti" birthdate="2007-06-22" gender="M" nation="BRA" license="407187" athleteid="1657" externalid="407187">
              <RESULTS>
                <RESULT eventid="1140" points="64" swimtime="00:00:55.25" resultid="1658" heatid="1898" lane="2" />
                <RESULT eventid="1096" points="74" swimtime="00:01:46.46" resultid="1659" heatid="1884" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="80" swimtime="00:00:46.71" resultid="1660" heatid="1956" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietro" lastname="Nabas De Assis" birthdate="2011-07-09" gender="M" nation="BRA" license="366968" swrid="5603878" athleteid="1461" externalid="366968">
              <RESULTS>
                <RESULT eventid="1184" points="285" swimtime="00:00:37.90" resultid="1462" heatid="1916" lane="5" entrytime="00:00:37.30" entrycourse="SCM" />
                <RESULT eventid="1074" points="252" swimtime="00:02:53.46" resultid="1463" heatid="1878" lane="6" entrytime="00:03:02.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.91" />
                    <SPLIT distance="100" swimtime="00:01:28.06" />
                    <SPLIT distance="150" swimtime="00:02:14.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="274" swimtime="00:00:31.03" resultid="1464" heatid="1957" lane="3" entrytime="00:00:31.48" entrycourse="SCM" />
                <RESULT eventid="1236" points="331" swimtime="00:01:19.87" resultid="1465" heatid="1929" lane="3" entrytime="00:01:24.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Gabriel Oliveira" birthdate="2006-05-31" gender="M" nation="BRA" license="345589" swrid="5603838" athleteid="1450" externalid="345589">
              <RESULTS>
                <RESULT eventid="1162" points="278" swimtime="00:01:13.20" resultid="1451" heatid="1908" lane="6" entrytime="00:01:10.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="427" swimtime="00:00:59.52" resultid="1452" heatid="1886" lane="5" entrytime="00:00:59.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="412" swimtime="00:00:27.08" resultid="1453" heatid="1959" lane="5" entrytime="00:00:27.20" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrielle" lastname="Borba" birthdate="2014-06-15" gender="F" nation="BRA" license="385705" swrid="5323267" athleteid="1519" externalid="385705">
              <RESULTS>
                <RESULT eventid="1296" points="111" swimtime="00:00:47.61" resultid="1520" heatid="1950" lane="4" entrytime="00:00:45.19" entrycourse="SCM" />
                <RESULT eventid="1274" points="100" swimtime="00:01:01.07" resultid="1521" heatid="1942" lane="4" entrytime="00:00:57.94" entrycourse="SCM" />
                <RESULT eventid="1248" points="94" swimtime="00:00:55.49" resultid="1522" heatid="1933" lane="2" entrytime="00:00:56.05" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Baldo De França" birthdate="2014-04-21" gender="M" nation="BRA" license="393773" swrid="5507467" athleteid="1587" externalid="393773">
              <RESULTS>
                <RESULT eventid="1299" points="60" swimtime="00:00:51.30" resultid="1588" heatid="1952" lane="2" entrytime="00:00:45.96" entrycourse="SCM" />
                <RESULT eventid="1277" points="74" swimtime="00:00:59.20" resultid="1589" heatid="1944" lane="2" entrytime="00:00:58.84" entrycourse="SCM" />
                <RESULT eventid="1225" points="90" swimtime="00:00:48.49" resultid="1590" heatid="1927" lane="4" entrytime="00:00:58.49" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lavinia" lastname="Bossoni" birthdate="2013-11-03" gender="F" nation="BRA" license="377260" swrid="5343093" athleteid="1491" externalid="377260">
              <RESULTS>
                <RESULT eventid="1148" points="138" swimtime="00:01:49.20" resultid="1492" heatid="1902" lane="5" entrytime="00:01:46.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="142" swimtime="00:00:48.30" resultid="1493" heatid="1889" lane="6" entrytime="00:00:47.25" entrycourse="SCM" />
                <RESULT eventid="1060" points="165" swimtime="00:03:21.01" resultid="1494" heatid="1872" lane="5" entrytime="00:03:25.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.22" />
                    <SPLIT distance="100" swimtime="00:01:37.95" />
                    <SPLIT distance="150" swimtime="00:02:31.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Garcia Cavalcante" birthdate="2008-08-11" gender="M" nation="BRA" license="369676" swrid="5603841" athleteid="1399" externalid="369676">
              <RESULTS>
                <RESULT eventid="1074" points="377" swimtime="00:02:31.72" resultid="1400" heatid="1878" lane="5" entrytime="00:02:36.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="100" swimtime="00:01:16.83" />
                    <SPLIT distance="150" swimtime="00:01:57.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="358" swimtime="00:00:28.39" resultid="1401" heatid="1956" lane="5" />
                <RESULT eventid="1236" points="424" swimtime="00:01:13.55" resultid="1402" heatid="1930" lane="5" entrytime="00:01:16.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Santos Carraro" birthdate="2014-06-04" gender="M" nation="BRA" license="392097" swrid="5603908" athleteid="1545" externalid="392097">
              <RESULTS>
                <RESULT eventid="1299" points="162" swimtime="00:00:36.98" resultid="1546" heatid="1952" lane="3" entrytime="00:00:39.08" entrycourse="SCM" />
                <RESULT eventid="1277" points="69" swimtime="00:01:00.65" resultid="1547" heatid="1944" lane="6" />
                <RESULT eventid="1225" points="96" swimtime="00:00:47.47" resultid="1548" heatid="1927" lane="3" entrytime="00:00:50.46" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ghelere" birthdate="2011-04-03" gender="F" nation="BRA" license="368146" swrid="5603843" athleteid="1466" externalid="368146">
              <RESULTS>
                <RESULT eventid="1154" points="177" swimtime="00:01:36.24" resultid="1467" heatid="1906" lane="1" entrytime="00:01:45.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="294" swimtime="00:01:15.53" resultid="1468" heatid="1882" lane="2" entrytime="00:01:13.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="254" swimtime="00:03:12.23" resultid="1469" heatid="1960" lane="2" entrytime="00:03:15.10" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Schuch Pimpao" birthdate="2010-12-31" gender="M" nation="BRA" license="355586" swrid="5588908" athleteid="1454" externalid="355586">
              <RESULTS>
                <RESULT eventid="1288" points="289" swimtime="00:01:13.05" resultid="1455" heatid="1947" lane="3" entrytime="00:01:20.43" entrycourse="SCM" />
                <RESULT eventid="1210" points="294" swimtime="00:05:19.20" resultid="1456" heatid="1924" lane="5" entrytime="00:05:23.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:15.21" />
                    <SPLIT distance="150" swimtime="00:01:54.75" />
                    <SPLIT distance="200" swimtime="00:02:35.79" />
                    <SPLIT distance="250" swimtime="00:03:18.10" />
                    <SPLIT distance="300" swimtime="00:03:59.79" />
                    <SPLIT distance="350" swimtime="00:04:41.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="De Correa" birthdate="2014-12-03" gender="M" nation="BRA" license="403387" swrid="5676286" athleteid="1614" externalid="403387">
              <RESULTS>
                <RESULT eventid="1299" points="96" swimtime="00:00:44.02" resultid="1615" heatid="1952" lane="5" entrytime="00:00:46.13" entrycourse="SCM" />
                <RESULT eventid="1277" points="62" swimtime="00:01:02.81" resultid="1616" heatid="1943" lane="2" />
                <RESULT eventid="1199" points="93" swimtime="00:01:38.62" resultid="1617" heatid="1920" lane="2" entrytime="00:01:45.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Novak Pinho" birthdate="2012-11-14" gender="M" nation="BRA" license="378199" swrid="5603879" athleteid="1507" externalid="378199">
              <RESULTS>
                <RESULT eventid="1173" points="163" swimtime="00:00:36.88" resultid="1508" heatid="1913" lane="1" entrytime="00:00:35.96" entrycourse="SCM" />
                <RESULT eventid="1107" points="134" swimtime="00:00:43.19" resultid="1509" heatid="1891" lane="2" entrytime="00:00:45.48" entrycourse="SCM" />
                <RESULT eventid="1063" points="194" swimtime="00:02:51.49" resultid="1510" heatid="1873" lane="3" entrytime="00:03:03.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                    <SPLIT distance="100" swimtime="00:01:21.83" />
                    <SPLIT distance="150" swimtime="00:02:08.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="1661" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Enrico" lastname="Santin Rezende" birthdate="2016-02-15" gender="M" nation="BRA" license="407196" athleteid="1865" externalid="407196">
              <RESULTS>
                <RESULT eventid="1272" points="25" swimtime="00:00:30.75" resultid="1866" heatid="1940" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Silverio Duarte" birthdate="2011-08-08" gender="M" nation="BRA" license="392138" swrid="5603913" athleteid="1795" externalid="392138">
              <RESULTS>
                <RESULT eventid="1140" points="43" swimtime="00:01:02.80" resultid="1796" heatid="1898" lane="3" />
                <RESULT eventid="1096" points="68" swimtime="00:01:49.84" resultid="1797" heatid="1884" lane="5" entrytime="00:02:09.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" status="DNS" swimtime="00:00:00.00" resultid="1798" heatid="1957" lane="1" entrytime="00:01:00.65" entrycourse="SCM" />
                <RESULT eventid="1262" status="DSQ" swimtime="00:01:00.59" resultid="1799" heatid="1937" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Valentina Gozaga" birthdate="2014-06-28" gender="F" nation="BRA" license="385709" swrid="5603924" athleteid="1766" externalid="385709">
              <RESULTS>
                <RESULT eventid="1296" points="178" swimtime="00:00:40.76" resultid="1767" heatid="1950" lane="3" entrytime="00:00:43.69" entrycourse="SCM" />
                <RESULT eventid="1248" points="132" swimtime="00:00:49.59" resultid="1768" heatid="1933" lane="4" entrytime="00:00:54.63" entrycourse="SCM" />
                <RESULT eventid="1196" points="133" swimtime="00:01:38.21" resultid="1769" heatid="1918" lane="4" entrytime="00:01:40.08" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Rossi" birthdate="2012-05-21" gender="M" nation="BRA" license="378346" swrid="5603901" athleteid="1716" externalid="378346">
              <RESULTS>
                <RESULT eventid="1173" points="225" swimtime="00:00:33.12" resultid="1717" heatid="1913" lane="4" entrytime="00:00:33.44" entrycourse="SCM" />
                <RESULT eventid="1107" points="189" swimtime="00:00:38.49" resultid="1718" heatid="1891" lane="1" entrytime="00:00:48.70" entrycourse="SCM" />
                <RESULT eventid="1085" points="143" swimtime="00:01:45.60" resultid="1719" heatid="1881" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Guinoza" birthdate="2013-01-06" gender="F" nation="BRA" license="392012" swrid="5510698" athleteid="1791" externalid="392012">
              <RESULTS>
                <RESULT eventid="1170" points="189" swimtime="00:00:39.92" resultid="1792" heatid="1910" lane="6" entrytime="00:00:44.42" entrycourse="SCM" />
                <RESULT eventid="1148" points="162" swimtime="00:01:43.57" resultid="1793" heatid="1901" lane="4" entrytime="00:01:57.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1082" points="197" swimtime="00:01:47.01" resultid="1794" heatid="1879" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elen" lastname="Torres Gomes" birthdate="2015-10-15" gender="F" nation="BRA" license="396850" swrid="5641777" athleteid="1808" externalid="396850">
              <RESULTS>
                <RESULT eventid="1296" status="DNS" swimtime="00:00:00.00" resultid="1809" heatid="1950" lane="1" entrytime="00:00:57.87" entrycourse="SCM" />
                <RESULT eventid="1274" status="DNS" swimtime="00:00:00.00" resultid="1810" heatid="1941" lane="3" />
                <RESULT eventid="1248" status="DNS" swimtime="00:00:00.00" resultid="1811" heatid="1933" lane="5" entrytime="00:01:02.37" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Pazinato" birthdate="2011-01-05" gender="M" nation="BRA" license="368149" swrid="5603889" athleteid="1736" externalid="368149">
              <RESULTS>
                <RESULT eventid="1096" points="282" swimtime="00:01:08.33" resultid="1737" heatid="1885" lane="1" entrytime="00:01:09.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="220" swimtime="00:03:01.48" resultid="1738" heatid="1877" lane="3" entrytime="00:03:03.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:22.61" />
                    <SPLIT distance="150" swimtime="00:02:21.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="277" swimtime="00:00:30.92" resultid="1739" heatid="1958" lane="1" entrytime="00:00:30.40" entrycourse="SCM" />
                <RESULT eventid="1288" points="230" swimtime="00:01:18.84" resultid="1740" heatid="1947" lane="4" entrytime="00:01:22.27" entrycourse="SCM" />
                <RESULT eventid="1210" points="264" swimtime="00:05:30.57" resultid="1741" heatid="1924" lane="6" entrytime="00:05:38.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                    <SPLIT distance="100" swimtime="00:01:18.94" />
                    <SPLIT distance="150" swimtime="00:02:01.07" />
                    <SPLIT distance="200" swimtime="00:02:43.21" />
                    <SPLIT distance="250" swimtime="00:03:26.57" />
                    <SPLIT distance="300" swimtime="00:04:09.21" />
                    <SPLIT distance="350" swimtime="00:04:51.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robsson" lastname="Tows Oliveira" birthdate="2014-03-05" gender="M" nation="BRA" license="392107" swrid="5603922" athleteid="1824" externalid="392107">
              <RESULTS>
                <RESULT eventid="1299" points="139" swimtime="00:00:38.87" resultid="1825" heatid="1952" lane="4" entrytime="00:00:40.49" entrycourse="SCM" />
                <RESULT eventid="1277" points="122" swimtime="00:00:50.22" resultid="1826" heatid="1944" lane="4" entrytime="00:00:49.66" entrycourse="SCM" />
                <RESULT eventid="1199" points="139" swimtime="00:01:26.48" resultid="1827" heatid="1920" lane="4" entrytime="00:01:26.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Gevaerd Verssutti Garcia" birthdate="2013-10-15" gender="F" nation="BRA" license="378404" swrid="5588723" athleteid="1752" externalid="378404">
              <RESULTS>
                <RESULT eventid="1148" points="162" swimtime="00:01:43.57" resultid="1753" heatid="1901" lane="3" entrytime="00:01:52.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="212" swimtime="00:00:42.32" resultid="1754" heatid="1889" lane="2" entrytime="00:00:44.74" entrycourse="SCM" />
                <RESULT eventid="1082" points="148" swimtime="00:01:57.83" resultid="1755" heatid="1880" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Livia" lastname="Eloisa Silva" birthdate="2012-03-03" gender="F" nation="BRA" license="399725" swrid="5651341" athleteid="1812" externalid="399725">
              <RESULTS>
                <RESULT eventid="1170" points="104" swimtime="00:00:48.70" resultid="1813" heatid="1909" lane="3" entrytime="00:00:45.25" entrycourse="SCM" />
                <RESULT eventid="1148" status="DSQ" swimtime="00:02:10.25" resultid="1814" heatid="1901" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="123" swimtime="00:00:50.69" resultid="1815" heatid="1888" lane="5" entrytime="00:00:56.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andressa" lastname="Zamarian Gouvea" birthdate="2007-09-18" gender="F" nation="BRA" license="318503" swrid="5603929" athleteid="1662" externalid="318503">
              <RESULTS>
                <RESULT eventid="1132" points="359" swimtime="00:00:35.52" resultid="1663" heatid="1897" lane="3" entrytime="00:00:35.29" entrycourse="SCM" />
                <RESULT eventid="1110" points="335" swimtime="00:21:46.88" resultid="1664" heatid="1892" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="354" swimtime="00:01:17.57" resultid="1665" heatid="1946" lane="4" entrytime="00:01:15.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="371" swimtime="00:00:33.90" resultid="1666" heatid="1935" lane="2" />
                <RESULT eventid="1202" points="369" swimtime="00:05:22.25" resultid="1667" heatid="1922" lane="4" entrytime="00:05:19.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                    <SPLIT distance="100" swimtime="00:01:15.13" />
                    <SPLIT distance="150" swimtime="00:01:56.33" />
                    <SPLIT distance="200" swimtime="00:02:36.60" />
                    <SPLIT distance="250" swimtime="00:03:18.13" />
                    <SPLIT distance="300" swimtime="00:03:59.56" />
                    <SPLIT distance="350" swimtime="00:04:42.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Fernandes Dantas" birthdate="2016-12-14" gender="M" nation="BRA" license="406932" athleteid="1863" externalid="406932">
              <RESULTS>
                <RESULT eventid="1272" points="29" swimtime="00:00:29.28" resultid="1864" heatid="1940" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Bilemjian Leszczynski" birthdate="2014-02-22" gender="M" nation="BRA" license="406924" athleteid="1843" externalid="406924">
              <RESULTS>
                <RESULT eventid="1277" points="72" swimtime="00:00:59.86" resultid="1844" heatid="1943" lane="5" />
                <RESULT eventid="1199" points="65" swimtime="00:01:51.25" resultid="1845" heatid="1920" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Ognibeni Paupitz" birthdate="2014-08-08" gender="F" nation="BRA" license="406923" athleteid="1840" externalid="406923">
              <RESULTS>
                <RESULT eventid="1296" points="113" swimtime="00:00:47.38" resultid="1841" heatid="1949" lane="4" />
                <RESULT eventid="1274" points="86" swimtime="00:01:04.07" resultid="1842" heatid="1941" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Lima Coelho" birthdate="2012-12-12" gender="M" nation="BRA" license="393775" swrid="5615959" athleteid="1828" externalid="393775">
              <RESULTS>
                <RESULT eventid="1173" points="145" swimtime="00:00:38.30" resultid="1829" heatid="1912" lane="4" entrytime="00:00:39.41" entrycourse="SCM" />
                <RESULT eventid="1151" status="DSQ" swimtime="00:01:42.30" resultid="1830" heatid="1903" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="142" swimtime="00:00:42.35" resultid="1831" heatid="1891" lane="6" entrytime="00:00:49.16" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Tiemi Yamaguchi" birthdate="2013-02-28" gender="F" nation="BRA" license="385707" swrid="5603920" athleteid="1756" externalid="385707">
              <RESULTS>
                <RESULT eventid="1148" points="242" swimtime="00:01:30.64" resultid="1757" heatid="1902" lane="4" entrytime="00:01:41.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1126" points="208" swimtime="00:01:31.14" resultid="1758" heatid="1894" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1082" points="245" swimtime="00:01:39.61" resultid="1759" heatid="1879" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Taparo" birthdate="2012-04-20" gender="F" nation="BRA" license="407283" athleteid="1867" externalid="407283">
              <RESULTS>
                <RESULT eventid="1170" points="198" swimtime="00:00:39.33" resultid="1868" heatid="1909" lane="5" />
                <RESULT eventid="1104" points="169" swimtime="00:00:45.66" resultid="1869" heatid="1887" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eloah" lastname="Frasson" birthdate="2012-06-14" gender="F" nation="BRA" license="378338" swrid="5577016" athleteid="1702" externalid="378338">
              <RESULTS>
                <RESULT eventid="1170" points="254" swimtime="00:00:36.19" resultid="1703" heatid="1911" lane="5" entrytime="00:00:36.93" entrycourse="SCM" />
                <RESULT eventid="1148" points="183" swimtime="00:01:39.50" resultid="1704" heatid="1900" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1082" points="259" swimtime="00:01:37.76" resultid="1705" heatid="1880" lane="4" entrytime="00:01:38.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Jacobsen Donati" birthdate="2011-07-14" gender="M" nation="BRA" license="391851" swrid="5615735" athleteid="1785" externalid="391851">
              <RESULTS>
                <RESULT eventid="1096" status="DNS" swimtime="00:00:00.00" resultid="1786" heatid="1885" lane="2" entrytime="00:01:06.76" entrycourse="SCM" />
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="1787" heatid="1877" lane="2" entrytime="00:03:05.14" entrycourse="SCM" />
                <RESULT eventid="1310" status="DNS" swimtime="00:00:00.00" resultid="1788" heatid="1958" lane="4" entrytime="00:00:29.84" entrycourse="SCM" />
                <RESULT eventid="1288" status="DNS" swimtime="00:00:00.00" resultid="1789" heatid="1947" lane="5" entrytime="00:01:24.87" entrycourse="SCM" />
                <RESULT eventid="1210" status="DNS" swimtime="00:00:00.00" resultid="1790" heatid="1923" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Moreschi" birthdate="2012-08-09" gender="M" nation="BRA" license="385715" swrid="5603876" athleteid="1773" externalid="385715">
              <RESULTS>
                <RESULT eventid="1151" points="166" swimtime="00:01:29.61" resultid="1774" heatid="1904" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="198" swimtime="00:01:34.81" resultid="1775" heatid="1881" lane="3" entrytime="00:01:46.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="205" swimtime="00:02:48.48" resultid="1776" heatid="1874" lane="2" entrytime="00:02:47.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:19.58" />
                    <SPLIT distance="150" swimtime="00:02:04.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theodoro" lastname="Marques Serra" birthdate="2009-11-24" gender="M" nation="BRA" license="370661" swrid="5603870" athleteid="1742" externalid="370661">
              <RESULTS>
                <RESULT eventid="1140" points="281" swimtime="00:00:33.73" resultid="1743" heatid="1899" lane="5" entrytime="00:00:37.61" entrycourse="SCM" />
                <RESULT eventid="1096" points="311" swimtime="00:01:06.17" resultid="1744" heatid="1886" lane="6" entrytime="00:01:04.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="348" swimtime="00:02:35.84" resultid="1745" heatid="1878" lane="2" entrytime="00:02:36.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                    <SPLIT distance="100" swimtime="00:01:11.59" />
                    <SPLIT distance="150" swimtime="00:01:59.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="324" swimtime="00:01:10.36" resultid="1746" heatid="1948" lane="1" entrytime="00:01:09.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1210" points="347" swimtime="00:05:01.90" resultid="1747" heatid="1923" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                    <SPLIT distance="100" swimtime="00:01:11.69" />
                    <SPLIT distance="150" swimtime="00:01:51.02" />
                    <SPLIT distance="200" swimtime="00:02:30.07" />
                    <SPLIT distance="250" swimtime="00:03:09.24" />
                    <SPLIT distance="300" swimtime="00:03:47.61" />
                    <SPLIT distance="350" swimtime="00:04:26.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alex" lastname="Junior" birthdate="2013-03-11" gender="M" nation="BRA" license="385710" swrid="5603860" athleteid="1770" externalid="385710">
              <RESULTS>
                <RESULT eventid="1173" points="79" swimtime="00:00:46.98" resultid="1771" heatid="1912" lane="6" entrytime="00:00:54.38" entrycourse="SCM" />
                <RESULT eventid="1107" status="DSQ" swimtime="00:00:54.38" resultid="1772" heatid="1890" lane="4" entrytime="00:01:00.82" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Scalise Drapzichinski" birthdate="2012-03-07" gender="F" nation="BRA" license="378349" swrid="5603909" athleteid="1720" externalid="378349">
              <RESULTS>
                <RESULT eventid="1170" points="353" swimtime="00:00:32.43" resultid="1721" heatid="1911" lane="3" entrytime="00:00:32.82" entrycourse="SCM" />
                <RESULT eventid="1104" points="263" swimtime="00:00:39.38" resultid="1722" heatid="1889" lane="3" entrytime="00:00:40.08" entrycourse="SCM" />
                <RESULT eventid="1082" status="DSQ" swimtime="00:01:25.31" resultid="1723" heatid="1880" lane="3" entrytime="00:01:35.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Dias Rezende" birthdate="2016-03-04" gender="F" nation="BRA" license="406930" athleteid="1861" externalid="406930">
              <RESULTS>
                <RESULT eventid="1270" points="22" swimtime="00:00:37.04" resultid="1862" heatid="1939" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eloah" lastname="Juvedi Trindade" birthdate="2011-03-05" gender="F" nation="BRA" license="396829" swrid="5641768" athleteid="1800" externalid="396829">
              <RESULTS>
                <RESULT eventid="1154" points="88" swimtime="00:02:01.15" resultid="1801" heatid="1906" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" status="DSQ" swimtime="00:03:34.53" resultid="1802" heatid="1875" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.77" />
                    <SPLIT distance="100" swimtime="00:01:46.57" />
                    <SPLIT distance="150" swimtime="00:02:45.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="221" swimtime="00:00:37.88" resultid="1803" heatid="1953" lane="3" entrytime="00:00:38.80" entrycourse="SCM" />
                <RESULT eventid="1280" points="183" swimtime="00:01:36.68" resultid="1804" heatid="1945" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="199" swimtime="00:01:46.73" resultid="1805" heatid="1973" lane="5" entrytime="00:01:49.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Bagatim" birthdate="2014-05-27" gender="F" nation="BRA" license="378353" swrid="5236649" athleteid="1728" externalid="378353">
              <RESULTS>
                <RESULT eventid="1274" points="181" swimtime="00:00:50.09" resultid="1729" heatid="1942" lane="3" entrytime="00:00:49.48" entrycourse="SCM" />
                <RESULT eventid="1222" points="211" swimtime="00:00:40.89" resultid="1730" heatid="1926" lane="3" entrytime="00:00:40.48" entrycourse="SCM" />
                <RESULT eventid="1196" points="216" swimtime="00:01:23.66" resultid="1731" heatid="1918" lane="3" entrytime="00:01:25.58" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Bilemjian Leszczynski" birthdate="2011-08-06" gender="M" nation="BRA" license="406925" athleteid="1846" externalid="406925">
              <RESULTS>
                <RESULT eventid="1184" status="DSQ" swimtime="00:00:50.25" resultid="1847" heatid="1915" lane="5" />
                <RESULT eventid="1096" points="135" swimtime="00:01:27.33" resultid="1848" heatid="1884" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="138" swimtime="00:00:38.92" resultid="1849" heatid="1957" lane="6" />
                <RESULT eventid="1262" status="DSQ" swimtime="00:00:48.19" resultid="1850" heatid="1937" lane="5" />
                <RESULT eventid="1236" status="DSQ" swimtime="00:01:51.03" resultid="1851" heatid="1929" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Britto" birthdate="2012-10-04" gender="M" nation="BRA" license="378350" swrid="5588566" athleteid="1724" externalid="378350">
              <RESULTS>
                <RESULT eventid="1173" points="274" swimtime="00:00:31.01" resultid="1725" heatid="1913" lane="5" entrytime="00:00:33.63" entrycourse="SCM" />
                <RESULT eventid="1107" points="227" swimtime="00:00:36.22" resultid="1726" heatid="1891" lane="3" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="1085" points="165" swimtime="00:01:40.71" resultid="1727" heatid="1881" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Azevedo Martins" birthdate="2014-07-05" gender="F" nation="BRA" license="401859" swrid="5661340" athleteid="1816" externalid="401859">
              <RESULTS>
                <RESULT eventid="1296" points="64" swimtime="00:00:57.20" resultid="1817" heatid="1949" lane="2" />
                <RESULT eventid="1274" points="88" swimtime="00:01:03.64" resultid="1818" heatid="1941" lane="4" />
                <RESULT eventid="1222" points="49" swimtime="00:01:06.21" resultid="1819" heatid="1926" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monique" lastname="Istake" birthdate="2012-04-03" gender="F" nation="BRA" license="372023" swrid="5603857" athleteid="1732" externalid="372023">
              <RESULTS>
                <RESULT eventid="1148" points="272" swimtime="00:01:27.14" resultid="1733" heatid="1902" lane="3" entrytime="00:01:31.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1126" points="255" swimtime="00:01:25.15" resultid="1734" heatid="1895" lane="3" entrytime="00:01:29.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="318" swimtime="00:02:41.60" resultid="1735" heatid="1872" lane="3" entrytime="00:02:43.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                    <SPLIT distance="100" swimtime="00:01:14.78" />
                    <SPLIT distance="150" swimtime="00:01:58.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabel" lastname="Rezende" birthdate="2013-12-13" gender="F" nation="BRA" license="370657" swrid="5603900" athleteid="1674" externalid="370657">
              <RESULTS>
                <RESULT eventid="1104" points="166" swimtime="00:00:45.88" resultid="1675" heatid="1888" lane="2" entrytime="00:00:51.33" entrycourse="SCM" />
                <RESULT eventid="1082" points="101" swimtime="00:02:13.62" resultid="1676" heatid="1879" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="181" swimtime="00:03:14.97" resultid="1677" heatid="1872" lane="2" entrytime="00:03:15.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                    <SPLIT distance="100" swimtime="00:01:30.28" />
                    <SPLIT distance="150" swimtime="00:02:23.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Souza" birthdate="2013-09-11" gender="M" nation="BRA" license="382211" swrid="5603916" athleteid="1832" externalid="382211">
              <RESULTS>
                <RESULT eventid="1173" points="171" swimtime="00:00:36.26" resultid="1833" heatid="1912" lane="3" entrytime="00:00:37.99" entrycourse="SCM" />
                <RESULT eventid="1151" points="143" swimtime="00:01:34.06" resultid="1834" heatid="1904" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="186" swimtime="00:02:54.02" resultid="1835" heatid="1873" lane="4" entrytime="00:03:09.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:21.90" />
                    <SPLIT distance="150" swimtime="00:02:09.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Kenji Yamaguchi" birthdate="2011-08-25" gender="M" nation="BRA" license="385708" swrid="5603862" athleteid="1760" externalid="385708">
              <RESULTS>
                <RESULT eventid="1162" points="174" swimtime="00:01:25.55" resultid="1761" heatid="1907" lane="4" entrytime="00:01:42.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="238" swimtime="00:02:56.77" resultid="1762" heatid="1877" lane="4" entrytime="00:03:04.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:20.91" />
                    <SPLIT distance="150" swimtime="00:02:14.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="223" swimtime="00:00:33.20" resultid="1763" heatid="1957" lane="2" entrytime="00:00:33.78" entrycourse="SCM" />
                <RESULT eventid="1262" points="243" swimtime="00:00:34.85" resultid="1764" heatid="1938" lane="6" entrytime="00:00:40.14" entrycourse="SCM" />
                <RESULT eventid="1236" points="220" swimtime="00:01:31.56" resultid="1765" heatid="1929" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Schmeiske Ruivo" birthdate="2013-10-21" gender="F" nation="BRA" license="402006" swrid="5661354" athleteid="1820" externalid="402006">
              <RESULTS>
                <RESULT eventid="1170" points="190" swimtime="00:00:39.85" resultid="1821" heatid="1910" lane="1" entrytime="00:00:43.39" entrycourse="SCM" />
                <RESULT eventid="1104" points="178" swimtime="00:00:44.88" resultid="1822" heatid="1888" lane="3" entrytime="00:00:48.59" entrycourse="SCM" />
                <RESULT eventid="1082" status="DSQ" swimtime="00:01:46.15" resultid="1823" heatid="1879" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Rezende" birthdate="2012-01-23" gender="F" nation="BRA" license="370669" swrid="5603899" athleteid="1748" externalid="370669">
              <RESULTS>
                <RESULT eventid="1170" points="186" swimtime="00:00:40.15" resultid="1749" heatid="1911" lane="1" entrytime="00:00:38.69" entrycourse="SCM" />
                <RESULT eventid="1148" points="144" swimtime="00:01:47.66" resultid="1750" heatid="1902" lane="2" entrytime="00:01:44.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="205" swimtime="00:03:06.94" resultid="1751" heatid="1872" lane="4" entrytime="00:03:13.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                    <SPLIT distance="100" swimtime="00:01:30.43" />
                    <SPLIT distance="150" swimtime="00:02:19.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Berto" birthdate="2008-10-22" gender="M" nation="BRA" license="378342" swrid="5312223" athleteid="1690" externalid="378342">
              <RESULTS>
                <RESULT eventid="1184" points="327" swimtime="00:00:36.18" resultid="1691" heatid="1916" lane="1" entrytime="00:00:37.44" entrycourse="SCM" />
                <RESULT eventid="1096" points="309" swimtime="00:01:06.32" resultid="1692" heatid="1884" lane="3" entrytime="00:01:11.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="274" swimtime="00:00:31.03" resultid="1693" heatid="1958" lane="2" entrytime="00:00:30.27" entrycourse="SCM" />
                <RESULT eventid="1262" points="235" swimtime="00:00:35.22" resultid="1694" heatid="1937" lane="1" />
                <RESULT eventid="1236" points="346" swimtime="00:01:18.71" resultid="1695" heatid="1930" lane="1" entrytime="00:01:17.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Ortega" birthdate="1999-08-05" gender="M" nation="BRA" license="383118" swrid="5603852" athleteid="1678" externalid="383118">
              <RESULTS>
                <RESULT eventid="1184" points="257" swimtime="00:00:39.23" resultid="1679" heatid="1914" lane="2" />
                <RESULT eventid="1140" points="363" swimtime="00:00:30.98" resultid="1680" heatid="1899" lane="2" entrytime="00:00:33.03" entrycourse="SCM" />
                <RESULT eventid="1074" points="317" swimtime="00:02:40.71" resultid="1681" heatid="1878" lane="1" entrytime="00:02:49.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                    <SPLIT distance="100" swimtime="00:01:10.20" />
                    <SPLIT distance="150" swimtime="00:01:59.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="396" swimtime="00:00:27.44" resultid="1682" heatid="1959" lane="1" entrytime="00:00:27.42" entrycourse="SCM" />
                <RESULT eventid="1210" points="301" swimtime="00:05:16.64" resultid="1683" heatid="1924" lane="1" entrytime="00:05:27.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                    <SPLIT distance="100" swimtime="00:01:09.03" />
                    <SPLIT distance="150" swimtime="00:01:48.72" />
                    <SPLIT distance="200" swimtime="00:02:29.37" />
                    <SPLIT distance="250" swimtime="00:03:10.16" />
                    <SPLIT distance="300" swimtime="00:03:52.59" />
                    <SPLIT distance="350" swimtime="00:04:35.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Stephany" birthdate="2012-07-27" gender="F" nation="BRA" license="382210" swrid="5603917" athleteid="1836" externalid="382210">
              <RESULTS>
                <RESULT eventid="1170" points="220" swimtime="00:00:37.96" resultid="1837" heatid="1911" lane="6" entrytime="00:00:39.26" entrycourse="SCM" />
                <RESULT eventid="1126" points="97" swimtime="00:01:57.62" resultid="1838" heatid="1895" lane="4" entrytime="00:01:52.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="173" swimtime="00:00:45.29" resultid="1839" heatid="1888" lane="4" entrytime="00:00:50.69" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Dias Rezende" birthdate="2016-03-04" gender="F" nation="BRA" license="406929" athleteid="1859" externalid="406929">
              <RESULTS>
                <RESULT eventid="1270" points="18" swimtime="00:00:39.90" resultid="1860" heatid="1939" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dante" lastname="Gabriel Rossi" birthdate="2016-01-19" gender="M" nation="BRA" license="406928" athleteid="1856" externalid="406928">
              <RESULTS>
                <RESULT eventid="1272" points="58" swimtime="00:00:23.35" resultid="1857" heatid="1940" lane="5" />
                <RESULT eventid="1194" points="46" swimtime="00:00:27.36" resultid="1858" heatid="1917" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Posser" birthdate="2013-02-07" gender="F" nation="BRA" license="378343" swrid="5603896" athleteid="1706" externalid="378343">
              <RESULTS>
                <RESULT eventid="1170" status="DNS" swimtime="00:00:00.00" resultid="1707" heatid="1910" lane="2" entrytime="00:00:42.80" entrycourse="SCM" />
                <RESULT eventid="1148" status="DNS" swimtime="00:00:00.00" resultid="1708" heatid="1901" lane="2" entrytime="00:02:05.76" entrycourse="SCM" />
                <RESULT eventid="1126" status="DNS" swimtime="00:00:00.00" resultid="1709" heatid="1895" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Traci Rodrigues" birthdate="2011-03-06" gender="M" nation="BRA" license="406927" athleteid="1852" externalid="406927">
              <RESULTS>
                <RESULT eventid="1184" status="DSQ" swimtime="00:00:49.60" resultid="1853" heatid="1914" lane="4" />
                <RESULT eventid="1140" points="103" swimtime="00:00:47.06" resultid="1854" heatid="1898" lane="5" />
                <RESULT eventid="1310" points="157" swimtime="00:00:37.34" resultid="1855" heatid="1956" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Braga" birthdate="2010-05-07" gender="M" nation="BRA" license="378345" swrid="5343953" athleteid="1710" externalid="378345">
              <RESULTS>
                <RESULT eventid="1184" points="358" swimtime="00:00:35.12" resultid="1711" heatid="1916" lane="6" entrytime="00:00:41.24" entrycourse="SCM" />
                <RESULT eventid="1096" points="306" swimtime="00:01:06.54" resultid="1712" heatid="1884" lane="4" entrytime="00:01:16.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="266" swimtime="00:00:31.33" resultid="1713" heatid="1958" lane="6" entrytime="00:00:30.73" entrycourse="SCM" />
                <RESULT eventid="1236" points="398" swimtime="00:01:15.11" resultid="1714" heatid="1930" lane="2" entrytime="00:01:16.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1210" points="327" swimtime="00:05:07.86" resultid="1715" heatid="1923" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                    <SPLIT distance="100" swimtime="00:01:12.04" />
                    <SPLIT distance="150" swimtime="00:01:51.46" />
                    <SPLIT distance="200" swimtime="00:02:31.10" />
                    <SPLIT distance="250" swimtime="00:03:10.92" />
                    <SPLIT distance="300" swimtime="00:03:50.51" />
                    <SPLIT distance="350" swimtime="00:04:29.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Jupi Takaki" birthdate="2013-03-26" gender="F" nation="BRA" license="391845" swrid="5603861" athleteid="1777" externalid="391845">
              <RESULTS>
                <RESULT eventid="1170" points="239" swimtime="00:00:36.91" resultid="1778" heatid="1910" lane="4" entrytime="00:00:40.56" entrycourse="SCM" />
                <RESULT eventid="1126" points="182" swimtime="00:01:35.27" resultid="1779" heatid="1894" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="214" swimtime="00:03:04.37" resultid="1780" heatid="1872" lane="1" entrytime="00:03:29.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                    <SPLIT distance="100" swimtime="00:01:29.13" />
                    <SPLIT distance="150" swimtime="00:02:18.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benicio" lastname="Garcia" birthdate="2011-09-09" gender="M" nation="BRA" license="378347" swrid="5603842" athleteid="1668" externalid="378347">
              <RESULTS>
                <RESULT eventid="1184" points="120" swimtime="00:00:50.57" resultid="1669" heatid="1915" lane="1" />
                <RESULT eventid="1162" points="113" swimtime="00:01:38.72" resultid="1670" heatid="1907" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="249" swimtime="00:00:35.10" resultid="1671" heatid="1899" lane="1" entrytime="00:00:38.66" entrycourse="SCM" />
                <RESULT eventid="1288" points="216" swimtime="00:01:20.44" resultid="1672" heatid="1947" lane="2" entrytime="00:01:23.52" entrycourse="SCM" />
                <RESULT eventid="1262" points="192" swimtime="00:00:37.70" resultid="1673" heatid="1937" lane="3" entrytime="00:00:47.01" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Drapzichinski" birthdate="2015-08-21" gender="M" nation="BRA" license="391848" swrid="5603890" athleteid="1781" externalid="391848">
              <RESULTS>
                <RESULT eventid="1299" points="103" swimtime="00:00:42.94" resultid="1782" heatid="1952" lane="1" entrytime="00:00:48.85" entrycourse="SCM" />
                <RESULT eventid="1251" points="71" swimtime="00:00:53.31" resultid="1783" heatid="1934" lane="3" entrytime="00:01:00.64" entrycourse="SCM" />
                <RESULT eventid="1199" points="95" swimtime="00:01:38.18" resultid="1784" heatid="1919" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Silveira De Almeida" birthdate="2008-07-08" gender="M" nation="BRA" license="368152" swrid="5603912" athleteid="1696" externalid="368152">
              <RESULTS>
                <RESULT eventid="1162" points="479" swimtime="00:01:01.06" resultid="1697" heatid="1908" lane="5" entrytime="00:01:03.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="332" swimtime="00:01:04.71" resultid="1698" heatid="1886" lane="1" entrytime="00:01:02.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="423" swimtime="00:02:26.03" resultid="1699" heatid="1878" lane="4" entrytime="00:02:33.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.58" />
                    <SPLIT distance="100" swimtime="00:01:07.78" />
                    <SPLIT distance="150" swimtime="00:01:52.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1262" points="471" swimtime="00:00:27.94" resultid="1700" heatid="1938" lane="5" entrytime="00:00:32.49" entrycourse="SCM" />
                <RESULT eventid="1210" points="357" swimtime="00:04:59.04" resultid="1701" heatid="1923" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:10.59" />
                    <SPLIT distance="150" swimtime="00:01:48.05" />
                    <SPLIT distance="200" swimtime="00:02:27.79" />
                    <SPLIT distance="250" swimtime="00:03:05.85" />
                    <SPLIT distance="300" swimtime="00:03:44.59" />
                    <SPLIT distance="350" swimtime="00:04:22.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marco" lastname="Manzotti Marchi" birthdate="2015-06-26" gender="M" nation="BRA" license="396849" swrid="5641769" athleteid="1806" externalid="396849">
              <RESULTS>
                <RESULT eventid="1225" status="DNS" swimtime="00:00:00.00" resultid="1807" heatid="1927" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Magalhães Rezende" birthdate="2010-05-29" gender="F" nation="BRA" license="366960" swrid="5588793" athleteid="1684" externalid="366960">
              <RESULTS>
                <RESULT eventid="1110" points="303" swimtime="00:22:31.63" resultid="1685" heatid="1892" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="331" swimtime="00:02:56.10" resultid="1686" heatid="1960" lane="3" entrytime="00:02:51.11" entrycourse="SCM" />
                <RESULT eventid="1302" points="329" swimtime="00:00:33.19" resultid="1687" heatid="1954" lane="3" entrytime="00:00:31.73" entrycourse="SCM" />
                <RESULT eventid="1228" points="299" swimtime="00:01:33.21" resultid="1688" heatid="1973" lane="4" entrytime="00:01:27.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="329" swimtime="00:05:34.86" resultid="1689" heatid="1922" lane="1" entrytime="00:05:27.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                    <SPLIT distance="100" swimtime="00:01:17.39" />
                    <SPLIT distance="150" swimtime="00:01:59.79" />
                    <SPLIT distance="200" swimtime="00:02:42.33" />
                    <SPLIT distance="250" swimtime="00:03:25.40" />
                    <SPLIT distance="300" swimtime="00:04:08.93" />
                    <SPLIT distance="350" swimtime="00:04:52.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15981" nation="BRA" region="PR" clubid="1318" swrid="93783" name="Quinto Nado" shortname="5º Nado">
          <ATHLETES>
            <ATHLETE firstname="Guilherme" lastname="Kikuchi Fujii" birthdate="2007-01-04" gender="M" nation="BRA" license="297805" swrid="5603863" athleteid="1319" externalid="297805" level="G-OLIMPICA">
              <RESULTS>
                <RESULT eventid="1162" points="536" swimtime="00:00:58.81" resultid="1320" heatid="1908" lane="3" entrytime="00:01:00.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="506" swimtime="00:00:56.25" resultid="1321" heatid="1886" lane="4" entrytime="00:00:54.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="491" swimtime="00:00:25.54" resultid="1322" heatid="1956" lane="2" />
                <RESULT eventid="1288" points="485" swimtime="00:01:01.50" resultid="1323" heatid="1948" lane="3" entrytime="00:01:01.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1236" points="596" swimtime="00:01:05.68" resultid="1324" heatid="1930" lane="4" entrytime="00:01:05.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Takemura Couto" birthdate="2010-02-08" gender="F" nation="BRA" license="376950" swrid="5603919" athleteid="1343" externalid="376950">
              <RESULTS>
                <RESULT eventid="1154" points="317" swimtime="00:01:19.27" resultid="1344" heatid="1905" lane="4" />
                <RESULT eventid="1088" points="458" swimtime="00:01:05.15" resultid="1345" heatid="1882" lane="4" entrytime="00:01:13.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="470" swimtime="00:00:29.49" resultid="1346" heatid="1955" lane="6" entrytime="00:00:30.90" entrycourse="SCM" />
                <RESULT eventid="1280" points="330" swimtime="00:01:19.39" resultid="1347" heatid="1946" lane="1" entrytime="00:01:18.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="276" swimtime="00:01:35.68" resultid="1348" heatid="1928" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Betina" lastname="Tramontini Queiroz" birthdate="2007-09-11" gender="F" nation="BRA" license="357155" swrid="5658063" athleteid="1331" externalid="357155" level="VIBE">
              <RESULTS>
                <RESULT eventid="1154" points="333" swimtime="00:01:17.92" resultid="1332" heatid="1906" lane="4" entrytime="00:01:21.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="495" swimtime="00:01:03.52" resultid="1333" heatid="1883" lane="3" entrytime="00:01:02.50" entrycourse="SCM" />
                <RESULT eventid="1302" points="478" swimtime="00:00:29.31" resultid="1334" heatid="1955" lane="5" entrytime="00:00:30.53" entrycourse="SCM" />
                <RESULT eventid="1228" points="379" swimtime="00:01:26.14" resultid="1335" heatid="1973" lane="3" entrytime="00:01:23.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="513" swimtime="00:04:48.88" resultid="1336" heatid="1922" lane="3" entrytime="00:04:43.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                    <SPLIT distance="100" swimtime="00:01:09.49" />
                    <SPLIT distance="150" swimtime="00:01:45.76" />
                    <SPLIT distance="200" swimtime="00:02:23.00" />
                    <SPLIT distance="250" swimtime="00:02:59.45" />
                    <SPLIT distance="300" swimtime="00:03:36.14" />
                    <SPLIT distance="350" swimtime="00:04:12.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Poletti Veiga" birthdate="2010-10-01" gender="F" nation="BRA" license="376951" swrid="5603895" athleteid="1337" externalid="376951">
              <RESULTS>
                <RESULT eventid="1154" points="309" swimtime="00:01:19.90" resultid="1338" heatid="1906" lane="2" entrytime="00:01:24.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="441" swimtime="00:01:05.98" resultid="1339" heatid="1883" lane="5" entrytime="00:01:07.45" entrycourse="SCM" />
                <RESULT eventid="1302" points="437" swimtime="00:00:30.20" resultid="1340" heatid="1955" lane="4" entrytime="00:00:30.36" entrycourse="SCM" />
                <RESULT eventid="1280" points="367" swimtime="00:01:16.62" resultid="1341" heatid="1946" lane="5" entrytime="00:01:18.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1254" points="385" swimtime="00:00:33.50" resultid="1342" heatid="1936" lane="2" entrytime="00:00:35.19" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Bordini Zocco" birthdate="2008-08-04" gender="F" nation="BRA" license="385677" swrid="5332871" athleteid="1325" externalid="385677">
              <RESULTS>
                <RESULT eventid="1154" points="301" swimtime="00:01:20.64" resultid="1326" heatid="1905" lane="2" />
                <RESULT eventid="1088" points="382" swimtime="00:01:09.23" resultid="1327" heatid="1882" lane="3" entrytime="00:01:12.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="370" swimtime="00:00:31.92" resultid="1328" heatid="1954" lane="5" entrytime="00:00:34.04" entrycourse="SCM" />
                <RESULT eventid="1280" points="314" swimtime="00:01:20.72" resultid="1329" heatid="1946" lane="6" entrytime="00:01:22.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="331" swimtime="00:01:30.10" resultid="1330" heatid="1973" lane="2" entrytime="00:01:32.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Gomes" birthdate="2011-12-03" gender="F" nation="BRA" license="382051" swrid="5603846" athleteid="1355" externalid="382051">
              <RESULTS>
                <RESULT eventid="1132" points="173" swimtime="00:00:45.25" resultid="1356" heatid="1897" lane="6" entrytime="00:00:47.17" entrycourse="SCM" />
                <RESULT eventid="1088" points="214" swimtime="00:01:23.97" resultid="1357" heatid="1882" lane="6" entrytime="00:01:31.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1302" points="212" swimtime="00:00:38.42" resultid="1358" heatid="1953" lane="4" entrytime="00:00:40.99" entrycourse="SCM" />
                <RESULT eventid="1254" points="127" swimtime="00:00:48.42" resultid="1359" heatid="1935" lane="4" />
                <RESULT eventid="1202" points="207" swimtime="00:06:30.70" resultid="1360" heatid="1921" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.77" />
                    <SPLIT distance="100" swimtime="00:01:32.68" />
                    <SPLIT distance="150" swimtime="00:02:22.54" />
                    <SPLIT distance="200" swimtime="00:03:11.81" />
                    <SPLIT distance="250" swimtime="00:04:01.89" />
                    <SPLIT distance="300" swimtime="00:04:52.76" />
                    <SPLIT distance="350" swimtime="00:05:41.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Clara Bobroff" birthdate="2013-02-09" gender="F" nation="BRA" license="391752" swrid="5419807" athleteid="1361" externalid="391752">
              <RESULTS>
                <RESULT eventid="1170" points="243" swimtime="00:00:36.74" resultid="1362" heatid="1910" lane="3" entrytime="00:00:39.49" entrycourse="SCM" />
                <RESULT eventid="1148" points="188" swimtime="00:01:38.53" resultid="1363" heatid="1902" lane="1" entrytime="00:01:50.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="213" swimtime="00:03:04.67" resultid="1364" heatid="1871" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Silva Telles" birthdate="2011-07-19" gender="M" nation="BRA" license="377311" swrid="5603911" athleteid="1349" externalid="377311">
              <RESULTS>
                <RESULT eventid="1184" points="190" swimtime="00:00:43.37" resultid="1350" heatid="1914" lane="3" />
                <RESULT eventid="1096" points="205" swimtime="00:01:15.97" resultid="1351" heatid="1884" lane="2" entrytime="00:01:27.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1310" points="195" swimtime="00:00:34.72" resultid="1352" heatid="1957" lane="5" entrytime="00:00:39.08" entrycourse="SCM" />
                <RESULT eventid="1262" points="111" swimtime="00:00:45.17" resultid="1353" heatid="1937" lane="6" />
                <RESULT eventid="1236" points="183" swimtime="00:01:37.25" resultid="1354" heatid="1929" lane="5" entrytime="00:01:49.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
