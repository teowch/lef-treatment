<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.79911">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Pato Branco" name="70º Jogos Escolares do Paraná (15/17 Anos) 2024" course="SCM" entrytype="INVITATION" hostclub="Secretaria do Esporte, Governo do Estado do Paraná" hostclub.url="https://www.esporte.pr.gov.br/" number="38312" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/newInterface/eventos/38312" startmethod="1" timing="AUTOMATIC" touchpad="ONESIDE" masters="F" state="PR" nation="BRA">
      <AGEDATE value="2024-01-01" type="YEAR" />
      <POOL lanemin="1" lanemax="8" />
      <FACILITY city="Pato Branco" nation="BRA" state="PR" street="Rua Bispo Dom Carlos Eduardo, 173" street2="La Salle" zip="85505-280" />
      <POINTTABLE pointtableid="3016" name="FINA Point Scoring" version="2023" />
      <QUALIFY from="2023-08-03" until="2024-08-02" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-08-03" daytime="09:10" endtime="12:21" number="1" officialmeeting="08:30" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1061" daytime="09:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1064" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1494" />
                    <RANKING order="2" place="2" resultid="1721" />
                    <RANKING order="3" place="3" resultid="1657" />
                    <RANKING order="4" place="4" resultid="1902" />
                    <RANKING order="5" place="5" resultid="1712" />
                    <RANKING order="6" place="6" resultid="1924" />
                    <RANKING order="7" place="7" resultid="1870" />
                    <RANKING order="8" place="8" resultid="1612" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1975" daytime="09:10" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1065" daytime="09:24" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1927" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1302" />
                    <RANKING order="2" place="2" resultid="1883" />
                    <RANKING order="3" place="3" resultid="1282" />
                    <RANKING order="4" place="4" resultid="1406" />
                    <RANKING order="5" place="5" resultid="1439" />
                    <RANKING order="6" place="-1" resultid="1523" />
                    <RANKING order="7" place="-1" resultid="1568" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1976" daytime="09:24" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1069" daytime="09:28" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1928" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1652" />
                    <RANKING order="2" place="2" resultid="1252" />
                    <RANKING order="3" place="3" resultid="1499" />
                    <RANKING order="4" place="4" resultid="1343" />
                    <RANKING order="5" place="-1" resultid="1669" />
                    <RANKING order="6" place="-1" resultid="1427" />
                    <RANKING order="7" place="-1" resultid="1593" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1977" daytime="09:28" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1073" daytime="09:46" gender="M" number="4" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1929" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1242" />
                    <RANKING order="2" place="2" resultid="1919" />
                    <RANKING order="3" place="3" resultid="1632" />
                    <RANKING order="4" place="4" resultid="1398" />
                    <RANKING order="5" place="5" resultid="1257" />
                    <RANKING order="6" place="6" resultid="1879" />
                    <RANKING order="7" place="7" resultid="1874" />
                    <RANKING order="8" place="8" resultid="1472" />
                    <RANKING order="9" place="9" resultid="1434" />
                    <RANKING order="10" place="10" resultid="1218" />
                    <RANKING order="11" place="11" resultid="1476" />
                    <RANKING order="12" place="-1" resultid="1825" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1978" daytime="09:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1979" daytime="09:48" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1077" daytime="09:52" gender="F" number="5" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1930" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1546" />
                    <RANKING order="2" place="2" resultid="1560" />
                    <RANKING order="3" place="2" resultid="1839" />
                    <RANKING order="4" place="4" resultid="1862" />
                    <RANKING order="5" place="5" resultid="1532" />
                    <RANKING order="6" place="6" resultid="1779" />
                    <RANKING order="7" place="7" resultid="1791" />
                    <RANKING order="8" place="8" resultid="1292" />
                    <RANKING order="9" place="9" resultid="1692" />
                    <RANKING order="10" place="10" resultid="1490" />
                    <RANKING order="11" place="11" resultid="1273" />
                    <RANKING order="12" place="12" resultid="1464" />
                    <RANKING order="13" place="13" resultid="1352" />
                    <RANKING order="14" place="14" resultid="1372" />
                    <RANKING order="15" place="15" resultid="1828" />
                    <RANKING order="16" place="16" resultid="1415" />
                    <RANKING order="17" place="17" resultid="1741" />
                    <RANKING order="18" place="18" resultid="1648" />
                    <RANKING order="19" place="19" resultid="1469" />
                    <RANKING order="20" place="20" resultid="1418" />
                    <RANKING order="21" place="21" resultid="1431" />
                    <RANKING order="22" place="-1" resultid="1390" />
                    <RANKING order="23" place="-1" resultid="1327" />
                    <RANKING order="24" place="-1" resultid="1359" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1980" daytime="09:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1981" daytime="09:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1982" daytime="09:58" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1081" daytime="10:22" gender="M" number="6" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1931" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1542" />
                    <RANKING order="2" place="2" resultid="1750" />
                    <RANKING order="3" place="3" resultid="1583" />
                    <RANKING order="4" place="4" resultid="1448" />
                    <RANKING order="5" place="5" resultid="1835" />
                    <RANKING order="6" place="6" resultid="1675" />
                    <RANKING order="7" place="7" resultid="1702" />
                    <RANKING order="8" place="8" resultid="1755" />
                    <RANKING order="9" place="9" resultid="1550" />
                    <RANKING order="10" place="10" resultid="1716" />
                    <RANKING order="11" place="11" resultid="1394" />
                    <RANKING order="12" place="12" resultid="1572" />
                    <RANKING order="13" place="13" resultid="1355" />
                    <RANKING order="14" place="14" resultid="1381" />
                    <RANKING order="15" place="15" resultid="1815" />
                    <RANKING order="16" place="16" resultid="1688" />
                    <RANKING order="17" place="17" resultid="1262" />
                    <RANKING order="18" place="18" resultid="1238" />
                    <RANKING order="19" place="19" resultid="1878" />
                    <RANKING order="20" place="20" resultid="1576" />
                    <RANKING order="21" place="21" resultid="1247" />
                    <RANKING order="22" place="22" resultid="1267" />
                    <RANKING order="23" place="23" resultid="1460" />
                    <RANKING order="24" place="24" resultid="1873" />
                    <RANKING order="25" place="25" resultid="1231" />
                    <RANKING order="26" place="26" resultid="1888" />
                    <RANKING order="27" place="27" resultid="1367" />
                    <RANKING order="28" place="28" resultid="1277" />
                    <RANKING order="29" place="29" resultid="1363" />
                    <RANKING order="30" place="30" resultid="1234" />
                    <RANKING order="31" place="31" resultid="1907" />
                    <RANKING order="32" place="32" resultid="1438" />
                    <RANKING order="33" place="-1" resultid="1210" />
                    <RANKING order="34" place="-1" resultid="1410" />
                    <RANKING order="35" place="-1" resultid="1810" />
                    <RANKING order="36" place="-1" resultid="1820" />
                    <RANKING order="37" place="-1" resultid="1588" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1983" daytime="10:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1984" daytime="10:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1985" daytime="10:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="1986" daytime="10:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="1987" daytime="10:32" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1085" daytime="10:36" gender="F" number="7" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1932" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1897" />
                    <RANKING order="2" place="2" resultid="1602" />
                    <RANKING order="3" place="3" resultid="1679" />
                    <RANKING order="4" place="4" resultid="1272" />
                    <RANKING order="5" place="5" resultid="1489" />
                    <RANKING order="6" place="6" resultid="1764" />
                    <RANKING order="7" place="7" resultid="1805" />
                    <RANKING order="8" place="8" resultid="1287" />
                    <RANKING order="9" place="9" resultid="1310" />
                    <RANKING order="10" place="10" resultid="1351" />
                    <RANKING order="11" place="11" resultid="1371" />
                    <RANKING order="12" place="12" resultid="1504" />
                    <RANKING order="13" place="13" resultid="1468" />
                    <RANKING order="14" place="14" resultid="1347" />
                    <RANKING order="15" place="15" resultid="1314" />
                    <RANKING order="16" place="16" resultid="1456" />
                    <RANKING order="17" place="17" resultid="1740" />
                    <RANKING order="18" place="18" resultid="1414" />
                    <RANKING order="19" place="19" resultid="1647" />
                    <RANKING order="20" place="20" resultid="1426" />
                    <RANKING order="21" place="21" resultid="1430" />
                    <RANKING order="22" place="-1" resultid="1389" />
                    <RANKING order="23" place="-1" resultid="1514" />
                    <RANKING order="24" place="-1" resultid="1735" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1988" daytime="10:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1989" daytime="10:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1990" daytime="10:42" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1089" daytime="10:58" gender="M" number="8" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1934" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1637" />
                    <RANKING order="2" place="2" resultid="1627" />
                    <RANKING order="3" place="3" resultid="1306" />
                    <RANKING order="4" place="4" resultid="1800" />
                    <RANKING order="5" place="-1" resultid="1402" />
                    <RANKING order="6" place="-1" resultid="1331" />
                    <RANKING order="7" place="-1" resultid="1769" />
                    <RANKING order="8" place="-1" resultid="1577" />
                    <RANKING order="9" place="-1" resultid="1597" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1991" daytime="10:58" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1093" daytime="11:04" gender="F" number="9" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1933" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1697" />
                    <RANKING order="2" place="2" resultid="1323" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1992" daytime="11:04" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1097" daytime="11:10" gender="M" number="10" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1935" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1731" />
                    <RANKING order="2" place="2" resultid="1759" />
                    <RANKING order="3" place="3" resultid="1543" />
                    <RANKING order="4" place="4" resultid="1519" />
                    <RANKING order="5" place="5" resultid="1858" />
                    <RANKING order="6" place="6" resultid="1555" />
                    <RANKING order="7" place="7" resultid="1283" />
                    <RANKING order="8" place="8" resultid="1783" />
                    <RANKING order="9" place="9" resultid="1509" />
                    <RANKING order="10" place="10" resultid="1382" />
                    <RANKING order="11" place="11" resultid="1339" />
                    <RANKING order="12" place="12" resultid="1527" />
                    <RANKING order="13" place="13" resultid="1551" />
                    <RANKING order="14" place="14" resultid="1318" />
                    <RANKING order="15" place="15" resultid="1461" />
                    <RANKING order="16" place="16" resultid="1385" />
                    <RANKING order="17" place="17" resultid="1479" />
                    <RANKING order="18" place="18" resultid="1617" />
                    <RANKING order="19" place="19" resultid="1910" />
                    <RANKING order="20" place="20" resultid="1227" />
                    <RANKING order="21" place="-1" resultid="1263" />
                    <RANKING order="22" place="-1" resultid="1215" />
                    <RANKING order="23" place="-1" resultid="1224" />
                    <RANKING order="24" place="-1" resultid="1221" />
                    <RANKING order="25" place="-1" resultid="1364" />
                    <RANKING order="26" place="-1" resultid="1821" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1993" daytime="11:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1994" daytime="11:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1995" daytime="11:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="1996" daytime="11:16" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1101" daytime="11:20" gender="F" number="11" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1936" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1774" />
                    <RANKING order="2" place="2" resultid="1297" />
                    <RANKING order="3" place="3" resultid="1607" />
                    <RANKING order="4" place="4" resultid="1622" />
                    <RANKING order="5" place="5" resultid="1796" />
                    <RANKING order="6" place="6" resultid="1843" />
                    <RANKING order="7" place="7" resultid="1344" />
                    <RANKING order="8" place="8" resultid="1373" />
                    <RANKING order="9" place="9" resultid="1315" />
                    <RANKING order="10" place="10" resultid="1452" />
                    <RANKING order="11" place="11" resultid="1422" />
                    <RANKING order="12" place="12" resultid="1457" />
                    <RANKING order="13" place="-1" resultid="1360" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1997" daytime="11:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1998" daytime="11:22" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1105" daytime="11:40" gender="M" number="12" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1938" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1661" />
                    <RANKING order="2" place="2" resultid="1707" />
                    <RANKING order="3" place="3" resultid="1335" />
                    <RANKING order="4" place="4" resultid="1642" />
                    <RANKING order="5" place="5" resultid="1853" />
                    <RANKING order="6" place="6" resultid="1684" />
                    <RANKING order="7" place="7" resultid="1787" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1999" daytime="11:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1109" daytime="12:02" gender="X" number="13" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1110" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1850" />
                    <RANKING order="2" place="2" resultid="1672" />
                    <RANKING order="3" place="3" resultid="1378" />
                    <RANKING order="4" place="4" resultid="1486" />
                    <RANKING order="5" place="5" resultid="1445" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2000" daytime="12:02" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-08-03" daytime="15:40" endtime="18:22" number="2" officialmeeting="15:00" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1111" daytime="15:40" gender="F" number="14" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1939" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1495" />
                    <RANKING order="2" place="2" resultid="1547" />
                    <RANKING order="3" place="3" resultid="1658" />
                    <RANKING order="4" place="4" resultid="1903" />
                    <RANKING order="5" place="5" resultid="1298" />
                    <RANKING order="6" place="6" resultid="1867" />
                    <RANKING order="7" place="7" resultid="1781" />
                    <RANKING order="8" place="8" resultid="1713" />
                    <RANKING order="9" place="9" resultid="1613" />
                    <RANKING order="10" place="-1" resultid="1515" />
                    <RANKING order="11" place="-1" resultid="1736" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2001" daytime="15:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2002" daytime="15:46" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1115" daytime="15:54" gender="M" number="15" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1940" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1584" />
                    <RANKING order="2" place="2" resultid="1564" />
                    <RANKING order="3" place="3" resultid="1662" />
                    <RANKING order="4" place="4" resultid="1884" />
                    <RANKING order="5" place="5" resultid="1854" />
                    <RANKING order="6" place="6" resultid="1685" />
                    <RANKING order="7" place="7" resultid="1689" />
                    <RANKING order="8" place="8" resultid="1368" />
                    <RANKING order="9" place="9" resultid="1537" />
                    <RANKING order="10" place="-1" resultid="1726" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2003" daytime="15:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2004" daytime="16:04" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1119" daytime="16:28" gender="F" number="16" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1941" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1670" />
                    <RANKING order="2" place="2" resultid="1608" />
                    <RANKING order="3" place="3" resultid="1775" />
                    <RANKING order="4" place="4" resultid="1500" />
                    <RANKING order="5" place="5" resultid="1844" />
                    <RANKING order="6" place="-1" resultid="1594" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2005" daytime="16:28" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1123" daytime="16:34" gender="M" number="17" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1942" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1732" />
                    <RANKING order="2" place="2" resultid="1760" />
                    <RANKING order="3" place="3" resultid="1859" />
                    <RANKING order="4" place="4" resultid="1665" />
                    <RANKING order="5" place="5" resultid="1556" />
                    <RANKING order="6" place="6" resultid="1784" />
                    <RANKING order="7" place="7" resultid="1788" />
                    <RANKING order="8" place="8" resultid="1407" />
                    <RANKING order="9" place="-1" resultid="1520" />
                    <RANKING order="10" place="-1" resultid="1643" />
                    <RANKING order="11" place="-1" resultid="1811" />
                    <RANKING order="12" place="-1" resultid="1569" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2006" daytime="16:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2007" daytime="16:38" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1127" daytime="16:44" gender="F" number="18" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1946" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1898" />
                    <RANKING order="2" place="2" resultid="1840" />
                    <RANKING order="3" place="3" resultid="1533" />
                    <RANKING order="4" place="4" resultid="1863" />
                    <RANKING order="5" place="5" resultid="1693" />
                    <RANKING order="6" place="6" resultid="1253" />
                    <RANKING order="7" place="7" resultid="1603" />
                    <RANKING order="8" place="8" resultid="1680" />
                    <RANKING order="9" place="9" resultid="1797" />
                    <RANKING order="10" place="10" resultid="1274" />
                    <RANKING order="11" place="11" resultid="1491" />
                    <RANKING order="12" place="12" resultid="1353" />
                    <RANKING order="13" place="13" resultid="1453" />
                    <RANKING order="14" place="14" resultid="1345" />
                    <RANKING order="15" place="15" resultid="1465" />
                    <RANKING order="16" place="16" resultid="1348" />
                    <RANKING order="17" place="17" resultid="1428" />
                    <RANKING order="18" place="18" resultid="1505" />
                    <RANKING order="19" place="19" resultid="1470" />
                    <RANKING order="20" place="20" resultid="1316" />
                    <RANKING order="21" place="21" resultid="1423" />
                    <RANKING order="22" place="22" resultid="1829" />
                    <RANKING order="23" place="23" resultid="1458" />
                    <RANKING order="24" place="24" resultid="1742" />
                    <RANKING order="25" place="25" resultid="1649" />
                    <RANKING order="26" place="26" resultid="1419" />
                    <RANKING order="27" place="-1" resultid="1806" />
                    <RANKING order="28" place="-1" resultid="1391" />
                    <RANKING order="29" place="-1" resultid="1516" />
                    <RANKING order="30" place="-1" resultid="1328" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2008" daytime="16:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2009" daytime="16:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2010" daytime="16:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2011" daytime="16:50" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1131" daytime="16:54" gender="M" number="19" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1945" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1544" />
                    <RANKING order="2" place="2" resultid="1449" />
                    <RANKING order="3" place="3" resultid="1836" />
                    <RANKING order="4" place="4" resultid="1510" />
                    <RANKING order="5" place="5" resultid="1756" />
                    <RANKING order="6" place="6" resultid="1676" />
                    <RANKING order="7" place="7" resultid="1703" />
                    <RANKING order="8" place="8" resultid="1308" />
                    <RANKING order="9" place="9" resultid="1552" />
                    <RANKING order="10" place="10" resultid="1243" />
                    <RANKING order="11" place="11" resultid="1396" />
                    <RANKING order="12" place="12" resultid="1336" />
                    <RANKING order="13" place="13" resultid="1717" />
                    <RANKING order="14" place="14" resultid="1264" />
                    <RANKING order="15" place="15" resultid="1239" />
                    <RANKING order="16" place="16" resultid="1340" />
                    <RANKING order="17" place="17" resultid="1383" />
                    <RANKING order="18" place="18" resultid="1880" />
                    <RANKING order="19" place="19" resultid="1356" />
                    <RANKING order="20" place="20" resultid="1746" />
                    <RANKING order="21" place="21" resultid="1268" />
                    <RANKING order="22" place="22" resultid="1473" />
                    <RANKING order="23" place="23" resultid="1399" />
                    <RANKING order="24" place="24" resultid="1875" />
                    <RANKING order="25" place="25" resultid="1211" />
                    <RANKING order="26" place="26" resultid="1232" />
                    <RANKING order="27" place="27" resultid="1278" />
                    <RANKING order="28" place="28" resultid="1258" />
                    <RANKING order="29" place="29" resultid="1480" />
                    <RANKING order="30" place="30" resultid="1618" />
                    <RANKING order="31" place="31" resultid="1386" />
                    <RANKING order="32" place="32" resultid="1319" />
                    <RANKING order="33" place="33" resultid="1911" />
                    <RANKING order="34" place="34" resultid="1889" />
                    <RANKING order="35" place="35" resultid="1477" />
                    <RANKING order="36" place="36" resultid="1219" />
                    <RANKING order="37" place="37" resultid="1216" />
                    <RANKING order="38" place="38" resultid="1235" />
                    <RANKING order="39" place="39" resultid="1435" />
                    <RANKING order="40" place="40" resultid="1832" />
                    <RANKING order="41" place="41" resultid="1225" />
                    <RANKING order="42" place="42" resultid="1222" />
                    <RANKING order="43" place="-1" resultid="1727" />
                    <RANKING order="44" place="-1" resultid="1822" />
                    <RANKING order="45" place="-1" resultid="1826" />
                    <RANKING order="46" place="-1" resultid="1848" />
                    <RANKING order="47" place="-1" resultid="1589" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2012" daytime="16:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2013" daytime="16:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2014" daytime="16:58" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2015" daytime="17:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2016" daytime="17:02" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2017" daytime="17:04" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1135" daytime="17:28" gender="F" number="20" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1944" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1561" />
                    <RANKING order="2" place="2" resultid="1653" />
                    <RANKING order="3" place="3" resultid="1623" />
                    <RANKING order="4" place="4" resultid="1792" />
                    <RANKING order="5" place="5" resultid="1780" />
                    <RANKING order="6" place="6" resultid="1293" />
                    <RANKING order="7" place="-1" resultid="1893" />
                    <RANKING order="8" place="-1" resultid="1925" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2018" daytime="17:28" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1139" daytime="17:34" gender="M" number="21" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1947" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1303" />
                    <RANKING order="2" place="2" resultid="1633" />
                    <RANKING order="3" place="3" resultid="1816" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2019" daytime="17:34" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1143" daytime="17:38" gender="F" number="22" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1948" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1324" />
                    <RANKING order="2" place="2" resultid="1765" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2020" daytime="17:38" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1147" daytime="17:42" gender="M" number="23" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1949" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1751" />
                    <RANKING order="2" place="2" resultid="1307" />
                    <RANKING order="3" place="3" resultid="1403" />
                    <RANKING order="4" place="4" resultid="1801" />
                    <RANKING order="5" place="5" resultid="1770" />
                    <RANKING order="6" place="6" resultid="1628" />
                    <RANKING order="7" place="7" resultid="1847" />
                    <RANKING order="8" place="8" resultid="1332" />
                    <RANKING order="9" place="9" resultid="1395" />
                    <RANKING order="10" place="10" resultid="1528" />
                    <RANKING order="11" place="11" resultid="1745" />
                    <RANKING order="12" place="12" resultid="1248" />
                    <RANKING order="13" place="13" resultid="1578" />
                    <RANKING order="14" place="-1" resultid="1573" />
                    <RANKING order="15" place="-1" resultid="1908" />
                    <RANKING order="16" place="-1" resultid="1411" />
                    <RANKING order="17" place="-1" resultid="1524" />
                    <RANKING order="18" place="-1" resultid="1598" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2021" daytime="17:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2022" daytime="17:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2023" daytime="17:48" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1151" daytime="17:58" gender="F" number="24" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1950" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1698" />
                    <RANKING order="2" place="2" resultid="1671" />
                    <RANKING order="3" place="3" resultid="1722" />
                    <RANKING order="4" place="-1" resultid="1288" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2024" daytime="17:58" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1155" daytime="18:06" gender="M" number="25" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1951" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1638" />
                    <RANKING order="2" place="2" resultid="1860" />
                    <RANKING order="3" place="3" resultid="1666" />
                    <RANKING order="4" place="4" resultid="1708" />
                    <RANKING order="5" place="-1" resultid="1599" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2025" daytime="18:06" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1159" daytime="18:30" gender="F" number="26" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1966" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1374" />
                    <RANKING order="2" place="2" resultid="1482" />
                    <RANKING order="3" place="3" resultid="1441" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2026" daytime="18:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1161" daytime="18:34" gender="M" number="27" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1965" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1443" />
                    <RANKING order="2" place="2" resultid="1376" />
                    <RANKING order="3" place="3" resultid="1484" />
                    <RANKING order="4" place="4" resultid="1228" />
                    <RANKING order="5" place="-1" resultid="1579" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2027" daytime="18:34" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-08-04" daytime="09:10" endtime="11:47" number="3" officialmeeting="08:30" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1163" daytime="09:10" gender="M" number="28" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1955" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1639" />
                    <RANKING order="2" place="2" resultid="1663" />
                    <RANKING order="3" place="3" resultid="1566" />
                    <RANKING order="4" place="4" resultid="1337" />
                    <RANKING order="5" place="5" resultid="1885" />
                    <RANKING order="6" place="6" resultid="1855" />
                    <RANKING order="7" place="7" resultid="1686" />
                    <RANKING order="8" place="8" resultid="1539" />
                    <RANKING order="9" place="-1" resultid="1320" />
                    <RANKING order="10" place="-1" resultid="1369" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2028" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2029" daytime="09:22" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1167" daytime="09:34" gender="F" number="29" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1954" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1548" />
                    <RANKING order="2" place="2" resultid="1562" />
                    <RANKING order="3" place="3" resultid="1841" />
                    <RANKING order="4" place="4" resultid="1864" />
                    <RANKING order="5" place="5" resultid="1654" />
                    <RANKING order="6" place="6" resultid="1793" />
                    <RANKING order="7" place="7" resultid="1904" />
                    <RANKING order="8" place="8" resultid="1294" />
                    <RANKING order="9" place="9" resultid="1845" />
                    <RANKING order="10" place="10" resultid="1311" />
                    <RANKING order="11" place="11" resultid="1466" />
                    <RANKING order="12" place="12" resultid="1420" />
                    <RANKING order="13" place="-1" resultid="1424" />
                    <RANKING order="14" place="-1" resultid="1432" />
                    <RANKING order="15" place="-1" resultid="1329" />
                    <RANKING order="16" place="-1" resultid="1766" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2030" daytime="09:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2031" daytime="09:38" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1171" daytime="09:42" gender="M" number="30" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1956" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1304" />
                    <RANKING order="2" place="2" resultid="1837" />
                    <RANKING order="3" place="3" resultid="1634" />
                    <RANKING order="4" place="4" resultid="1920" />
                    <RANKING order="5" place="5" resultid="1244" />
                    <RANKING order="6" place="6" resultid="1817" />
                    <RANKING order="7" place="7" resultid="1249" />
                    <RANKING order="8" place="8" resultid="1677" />
                    <RANKING order="9" place="9" resultid="1400" />
                    <RANKING order="10" place="10" resultid="1259" />
                    <RANKING order="11" place="11" resultid="1474" />
                    <RANKING order="12" place="12" resultid="1538" />
                    <RANKING order="13" place="-1" resultid="1436" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2032" daytime="09:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2033" daytime="09:46" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1175" daytime="09:58" gender="F" number="31" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1957" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1699" />
                    <RANKING order="2" place="2" resultid="1899" />
                    <RANKING order="3" place="3" resultid="1694" />
                    <RANKING order="4" place="4" resultid="1681" />
                    <RANKING order="5" place="5" resultid="1312" />
                    <RANKING order="6" place="6" resultid="1916" />
                    <RANKING order="7" place="7" resultid="1416" />
                    <RANKING order="8" place="-1" resultid="1894" />
                    <RANKING order="9" place="-1" resultid="1737" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2034" daytime="09:58" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1179" daytime="10:04" gender="M" number="32" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1953" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1585" />
                    <RANKING order="2" place="2" resultid="1752" />
                    <RANKING order="3" place="3" resultid="1565" />
                    <RANKING order="4" place="4" resultid="1450" />
                    <RANKING order="5" place="5" resultid="1709" />
                    <RANKING order="6" place="6" resultid="1629" />
                    <RANKING order="7" place="7" resultid="1644" />
                    <RANKING order="8" place="8" resultid="1690" />
                    <RANKING order="9" place="9" resultid="1747" />
                    <RANKING order="10" place="10" resultid="1890" />
                    <RANKING order="11" place="-1" resultid="1757" />
                    <RANKING order="12" place="-1" resultid="1590" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2035" daytime="10:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2036" daytime="10:08" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1183" daytime="10:34" gender="F" number="33" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1959" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1325" />
                    <RANKING order="2" place="2" resultid="1534" />
                    <RANKING order="3" place="3" resultid="1254" />
                    <RANKING order="4" place="4" resultid="1604" />
                    <RANKING order="5" place="5" resultid="1798" />
                    <RANKING order="6" place="6" resultid="1289" />
                    <RANKING order="7" place="7" resultid="1349" />
                    <RANKING order="8" place="8" resultid="1506" />
                    <RANKING order="9" place="-1" resultid="1807" />
                    <RANKING order="10" place="-1" resultid="1454" />
                    <RANKING order="11" place="-1" resultid="1595" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2037" daytime="10:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2038" daytime="10:38" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1187" daytime="10:40" gender="M" number="34" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1961" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1802" />
                    <RANKING order="2" place="2" resultid="1333" />
                    <RANKING order="3" place="3" resultid="1849" />
                    <RANKING order="4" place="4" resultid="1771" />
                    <RANKING order="5" place="5" resultid="1704" />
                    <RANKING order="6" place="6" resultid="1529" />
                    <RANKING order="7" place="7" resultid="1921" />
                    <RANKING order="8" place="8" resultid="1240" />
                    <RANKING order="9" place="9" resultid="1269" />
                    <RANKING order="10" place="10" resultid="1212" />
                    <RANKING order="11" place="11" resultid="1440" />
                    <RANKING order="12" place="12" resultid="1279" />
                    <RANKING order="13" place="-1" resultid="1357" />
                    <RANKING order="14" place="-1" resultid="1912" />
                    <RANKING order="15" place="-1" resultid="1404" />
                    <RANKING order="16" place="-1" resultid="1412" />
                    <RANKING order="17" place="-1" resultid="1525" />
                    <RANKING order="18" place="-1" resultid="1728" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2039" daytime="10:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2040" daytime="10:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2041" daytime="10:44" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1191" daytime="10:52" gender="F" number="35" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1960" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1776" />
                    <RANKING order="2" place="2" resultid="1299" />
                    <RANKING order="3" place="3" resultid="1609" />
                    <RANKING order="4" place="4" resultid="1501" />
                    <RANKING order="5" place="5" resultid="1624" />
                    <RANKING order="6" place="-1" resultid="1361" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2042" daytime="10:52" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1195" daytime="10:56" gender="M" number="36" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1962" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1733" />
                    <RANKING order="2" place="2" resultid="1761" />
                    <RANKING order="3" place="3" resultid="1521" />
                    <RANKING order="4" place="4" resultid="1557" />
                    <RANKING order="5" place="5" resultid="1667" />
                    <RANKING order="6" place="6" resultid="1284" />
                    <RANKING order="7" place="7" resultid="1785" />
                    <RANKING order="8" place="8" resultid="1574" />
                    <RANKING order="9" place="9" resultid="1511" />
                    <RANKING order="10" place="10" resultid="1341" />
                    <RANKING order="11" place="11" resultid="1718" />
                    <RANKING order="12" place="12" resultid="1408" />
                    <RANKING order="13" place="13" resultid="1365" />
                    <RANKING order="14" place="14" resultid="1462" />
                    <RANKING order="15" place="15" resultid="1619" />
                    <RANKING order="16" place="16" resultid="1481" />
                    <RANKING order="17" place="-1" resultid="1387" />
                    <RANKING order="18" place="-1" resultid="1812" />
                    <RANKING order="19" place="-1" resultid="1570" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2043" daytime="10:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2044" daytime="11:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2045" daytime="11:02" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1199" daytime="11:10" gender="F" number="37" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1963" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1496" />
                    <RANKING order="2" place="2" resultid="1723" />
                    <RANKING order="3" place="3" resultid="1659" />
                    <RANKING order="4" place="4" resultid="1868" />
                    <RANKING order="5" place="5" resultid="1926" />
                    <RANKING order="6" place="6" resultid="1871" />
                    <RANKING order="7" place="7" resultid="1614" />
                    <RANKING order="8" place="-1" resultid="1915" />
                    <RANKING order="9" place="-1" resultid="1714" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2046" daytime="11:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2047" daytime="11:32" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1203" daytime="12:12" gender="M" number="38" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1964" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1377" />
                    <RANKING order="2" place="2" resultid="1485" />
                    <RANKING order="3" place="3" resultid="1444" />
                    <RANKING order="4" place="-1" resultid="1580" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2048" daytime="12:12" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1205" daytime="12:18" gender="F" number="39" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1206" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1375" />
                    <RANKING order="2" place="2" resultid="1483" />
                    <RANKING order="3" place="-1" resultid="1442" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2049" daytime="12:18" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="17659" nation="BRA" region="PR" clubid="1507" name="International School Of Curitiba" shortname="Ctba-International,E">
          <ATHLETES>
            <ATHLETE firstname="Miguel" lastname="Faria Del Valle" birthdate="2009-08-28" gender="M" nation="BRA" license="376328" swrid="5600155" athleteid="1508" externalid="376328">
              <RESULTS>
                <RESULT eventid="1097" points="382" swimtime="00:00:34.36" resultid="1509" heatid="1996" lane="8" entrytime="00:00:33.04" entrycourse="SCM" />
                <RESULT eventid="1131" points="478" swimtime="00:00:25.77" resultid="1510" heatid="2017" lane="3" entrytime="00:00:25.18" entrycourse="SCM" />
                <RESULT eventid="1195" points="350" swimtime="00:01:18.39" resultid="1511" heatid="2043" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="10599" nation="BRA" region="PR" clubid="1767" name="Colégio Integral, Maringá" shortname="Mrga-Integral,C">
          <ATHLETES>
            <ATHLETE firstname="Lucas" lastname="Silveira De Almeida" birthdate="2008-07-08" gender="M" nation="BRA" license="368152" swrid="5603912" athleteid="1768" externalid="368152">
              <RESULTS>
                <RESULT eventid="1089" status="DSQ" swimtime="00:02:39.55" resultid="1769" heatid="1991" lane="5" entrytime="00:02:17.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                    <SPLIT distance="100" swimtime="00:01:09.96" />
                    <SPLIT distance="150" swimtime="00:01:54.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="397" swimtime="00:01:04.97" resultid="1770" heatid="2023" lane="5" entrytime="00:01:01.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="445" swimtime="00:00:28.48" resultid="1771" heatid="2041" lane="6" entrytime="00:00:27.94" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6577" nation="BRA" region="PR" clubid="1762" name="Colégio Dom Bosco, Maringá" shortname="Mrga-Dom Bosco,C">
          <ATHLETES>
            <ATHLETE firstname="Daniela" lastname="Inoue" birthdate="2008-10-31" gender="F" nation="BRA" license="378348" swrid="5603856" athleteid="1763" externalid="378348">
              <RESULTS>
                <RESULT eventid="1085" points="343" swimtime="00:01:11.76" resultid="1764" heatid="1990" lane="1" entrytime="00:01:10.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="233" swimtime="00:01:27.78" resultid="1765" heatid="2020" lane="5" entrytime="00:01:25.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" status="WDR" swimtime="00:00:00.00" resultid="1766" heatid="2030" lane="4" entrytime="00:01:23.34" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18907" nation="BRA" region="PR" clubid="1492" name="Colégio Dynâmico, Curitiba" shortname="Ctba-Dynâmico,C">
          <ATHLETES>
            <ATHLETE firstname="Isabelly" lastname="Sinnott" birthdate="2009-03-14" gender="F" nation="BRA" license="367255" swrid="5600258" athleteid="1493" externalid="367255">
              <RESULTS>
                <RESULT eventid="1061" points="551" swimtime="00:09:42.01" resultid="1494" heatid="1975" lane="4" entrytime="00:09:44.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="100" swimtime="00:01:08.21" />
                    <SPLIT distance="150" swimtime="00:01:44.15" />
                    <SPLIT distance="200" swimtime="00:02:20.57" />
                    <SPLIT distance="250" swimtime="00:02:57.42" />
                    <SPLIT distance="300" swimtime="00:03:34.21" />
                    <SPLIT distance="350" swimtime="00:04:11.13" />
                    <SPLIT distance="400" swimtime="00:04:48.18" />
                    <SPLIT distance="450" swimtime="00:05:24.86" />
                    <SPLIT distance="500" swimtime="00:06:01.70" />
                    <SPLIT distance="550" swimtime="00:06:38.46" />
                    <SPLIT distance="600" swimtime="00:07:15.51" />
                    <SPLIT distance="650" swimtime="00:07:52.18" />
                    <SPLIT distance="700" swimtime="00:08:29.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="560" swimtime="00:04:40.54" resultid="1495" heatid="2002" lane="5" entrytime="00:04:40.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:08.06" />
                    <SPLIT distance="150" swimtime="00:01:43.32" />
                    <SPLIT distance="200" swimtime="00:02:18.78" />
                    <SPLIT distance="250" swimtime="00:02:54.12" />
                    <SPLIT distance="300" swimtime="00:03:29.25" />
                    <SPLIT distance="350" swimtime="00:04:04.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" points="535" swimtime="00:18:38.54" resultid="1496" heatid="2047" lane="4" entrytime="00:18:34.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                    <SPLIT distance="100" swimtime="00:01:11.57" />
                    <SPLIT distance="150" swimtime="00:01:48.95" />
                    <SPLIT distance="200" swimtime="00:02:26.22" />
                    <SPLIT distance="250" swimtime="00:03:03.19" />
                    <SPLIT distance="300" swimtime="00:03:40.60" />
                    <SPLIT distance="350" swimtime="00:04:18.22" />
                    <SPLIT distance="400" swimtime="00:04:56.00" />
                    <SPLIT distance="450" swimtime="00:05:34.21" />
                    <SPLIT distance="500" swimtime="00:06:12.11" />
                    <SPLIT distance="550" swimtime="00:06:49.91" />
                    <SPLIT distance="600" swimtime="00:07:27.99" />
                    <SPLIT distance="650" swimtime="00:08:06.15" />
                    <SPLIT distance="700" swimtime="00:08:43.33" />
                    <SPLIT distance="750" swimtime="00:09:21.04" />
                    <SPLIT distance="800" swimtime="00:09:58.38" />
                    <SPLIT distance="850" swimtime="00:10:36.14" />
                    <SPLIT distance="900" swimtime="00:11:13.26" />
                    <SPLIT distance="950" swimtime="00:11:50.72" />
                    <SPLIT distance="1000" swimtime="00:12:27.86" />
                    <SPLIT distance="1050" swimtime="00:13:04.88" />
                    <SPLIT distance="1100" swimtime="00:13:41.85" />
                    <SPLIT distance="1150" swimtime="00:14:18.97" />
                    <SPLIT distance="1200" swimtime="00:14:56.23" />
                    <SPLIT distance="1250" swimtime="00:15:33.72" />
                    <SPLIT distance="1300" swimtime="00:16:11.33" />
                    <SPLIT distance="1350" swimtime="00:16:48.56" />
                    <SPLIT distance="1400" swimtime="00:17:26.21" />
                    <SPLIT distance="1450" swimtime="00:18:02.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17690" nation="BRA" region="PR" clubid="1823" name="6º Colégio Da Polícia Militar, Pato Branco" shortname="Pcbo-6ºcpm,C">
          <ATHLETES>
            <ATHLETE firstname="Arthur" lastname="Silva Figueiredo" birthdate="2009-03-30" gender="M" nation="BRA" license="V383381" athleteid="1824" externalid="V383381">
              <RESULTS>
                <RESULT eventid="1073" status="DNS" swimtime="00:00:00.00" resultid="1825" heatid="1978" lane="6" />
                <RESULT eventid="1131" status="DNS" swimtime="00:00:00.00" resultid="1826" heatid="2014" lane="5" entrytime="00:00:33.34" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sara" lastname="Piassa" birthdate="2009-08-07" gender="F" nation="BRA" license="V383175" athleteid="1827" externalid="V383175">
              <RESULTS>
                <RESULT eventid="1077" points="142" swimtime="00:00:48.33" resultid="1828" heatid="1981" lane="6" entrytime="00:00:45.26" entrycourse="SCM" />
                <RESULT eventid="1127" points="184" swimtime="00:00:40.30" resultid="1829" heatid="2010" lane="1" entrytime="00:00:38.61" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6536" nation="BRA" region="PR" clubid="1865" name="Colégio Diocesano Leão XIII, Paranaguá" shortname="Pgua-Leão XIII,C">
          <ATHLETES>
            <ATHLETE firstname="Gabriela" lastname="Marcelino De Souza" birthdate="2009-05-28" gender="F" nation="BRA" license="V414480" athleteid="1869" externalid="V414480">
              <RESULTS>
                <RESULT eventid="1061" points="317" swimtime="00:11:39.62" resultid="1870" heatid="1975" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.54" />
                    <SPLIT distance="100" swimtime="00:01:22.39" />
                    <SPLIT distance="150" swimtime="00:02:05.82" />
                    <SPLIT distance="200" swimtime="00:02:50.48" />
                    <SPLIT distance="250" swimtime="00:03:34.99" />
                    <SPLIT distance="300" swimtime="00:04:18.41" />
                    <SPLIT distance="350" swimtime="00:05:03.42" />
                    <SPLIT distance="400" swimtime="00:05:46.99" />
                    <SPLIT distance="450" swimtime="00:06:31.76" />
                    <SPLIT distance="500" swimtime="00:07:16.32" />
                    <SPLIT distance="550" swimtime="00:08:00.96" />
                    <SPLIT distance="600" swimtime="00:08:44.77" />
                    <SPLIT distance="650" swimtime="00:09:29.45" />
                    <SPLIT distance="700" swimtime="00:10:13.16" />
                    <SPLIT distance="750" swimtime="00:10:57.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" points="302" swimtime="00:22:33.24" resultid="1871" heatid="2047" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.09" />
                    <SPLIT distance="100" swimtime="00:01:22.48" />
                    <SPLIT distance="150" swimtime="00:02:07.47" />
                    <SPLIT distance="200" swimtime="00:02:52.84" />
                    <SPLIT distance="250" swimtime="00:03:38.35" />
                    <SPLIT distance="300" swimtime="00:04:24.13" />
                    <SPLIT distance="350" swimtime="00:05:10.39" />
                    <SPLIT distance="400" swimtime="00:05:56.05" />
                    <SPLIT distance="450" swimtime="00:06:42.01" />
                    <SPLIT distance="500" swimtime="00:07:27.79" />
                    <SPLIT distance="550" swimtime="00:08:13.15" />
                    <SPLIT distance="600" swimtime="00:08:58.49" />
                    <SPLIT distance="650" swimtime="00:09:43.82" />
                    <SPLIT distance="700" swimtime="00:10:29.19" />
                    <SPLIT distance="750" swimtime="00:11:14.61" />
                    <SPLIT distance="800" swimtime="00:12:00.00" />
                    <SPLIT distance="850" swimtime="00:12:45.51" />
                    <SPLIT distance="900" swimtime="00:13:31.26" />
                    <SPLIT distance="950" swimtime="00:14:17.04" />
                    <SPLIT distance="1000" swimtime="00:15:02.78" />
                    <SPLIT distance="1050" swimtime="00:15:48.37" />
                    <SPLIT distance="1100" swimtime="00:16:34.44" />
                    <SPLIT distance="1150" swimtime="00:17:20.63" />
                    <SPLIT distance="1200" swimtime="00:18:06.81" />
                    <SPLIT distance="1250" swimtime="00:18:52.22" />
                    <SPLIT distance="1300" swimtime="00:19:38.20" />
                    <SPLIT distance="1350" swimtime="00:20:22.49" />
                    <SPLIT distance="1400" swimtime="00:21:07.42" />
                    <SPLIT distance="1450" swimtime="00:21:50.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolle" lastname="Akemi Wajima" birthdate="2008-02-01" gender="F" nation="BRA" license="399346" swrid="5658056" athleteid="1866" externalid="399346">
              <RESULTS>
                <RESULT eventid="1111" points="400" swimtime="00:05:13.92" resultid="1867" heatid="2001" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:10.37" />
                    <SPLIT distance="150" swimtime="00:01:50.26" />
                    <SPLIT distance="200" swimtime="00:02:30.97" />
                    <SPLIT distance="250" swimtime="00:03:11.51" />
                    <SPLIT distance="300" swimtime="00:03:52.59" />
                    <SPLIT distance="350" swimtime="00:04:33.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" points="388" swimtime="00:20:44.86" resultid="1868" heatid="2047" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                    <SPLIT distance="100" swimtime="00:01:13.00" />
                    <SPLIT distance="150" swimtime="00:01:53.10" />
                    <SPLIT distance="200" swimtime="00:02:34.48" />
                    <SPLIT distance="250" swimtime="00:03:15.86" />
                    <SPLIT distance="300" swimtime="00:03:57.87" />
                    <SPLIT distance="350" swimtime="00:04:39.06" />
                    <SPLIT distance="400" swimtime="00:05:19.12" />
                    <SPLIT distance="450" swimtime="00:06:00.68" />
                    <SPLIT distance="500" swimtime="00:06:41.98" />
                    <SPLIT distance="550" swimtime="00:07:23.62" />
                    <SPLIT distance="600" swimtime="00:08:05.50" />
                    <SPLIT distance="650" swimtime="00:08:47.49" />
                    <SPLIT distance="700" swimtime="00:09:30.08" />
                    <SPLIT distance="750" swimtime="00:10:12.23" />
                    <SPLIT distance="800" swimtime="00:10:54.06" />
                    <SPLIT distance="850" swimtime="00:11:36.60" />
                    <SPLIT distance="900" swimtime="00:12:18.65" />
                    <SPLIT distance="950" swimtime="00:13:00.03" />
                    <SPLIT distance="1000" swimtime="00:13:42.90" />
                    <SPLIT distance="1050" swimtime="00:14:24.72" />
                    <SPLIT distance="1150" swimtime="00:15:49.60" />
                    <SPLIT distance="1200" swimtime="00:16:32.18" />
                    <SPLIT distance="1250" swimtime="00:17:14.66" />
                    <SPLIT distance="1300" swimtime="00:17:57.61" />
                    <SPLIT distance="1350" swimtime="00:18:39.70" />
                    <SPLIT distance="1400" swimtime="00:19:22.40" />
                    <SPLIT distance="1450" swimtime="00:20:05.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Alves Goncalves" birthdate="2008-10-30" gender="M" nation="BRA" license="V414514" athleteid="1872" externalid="V414514">
              <RESULTS>
                <RESULT eventid="1081" points="263" swimtime="00:01:09.98" resultid="1873" heatid="1984" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1073" points="221" swimtime="00:00:36.56" resultid="1874" heatid="1978" lane="4" />
                <RESULT eventid="1131" points="298" swimtime="00:00:30.15" resultid="1875" heatid="2013" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17319" nation="BRA" region="PR" clubid="1900" name="Colégio Estadual Eunice Borges Da Rocha, Sjpi" shortname="Sjpi-Euniceborges,Ce">
          <ATHLETES>
            <ATHLETE firstname="Monike" lastname="Lemos Carvalho" birthdate="2008-03-28" gender="F" nation="BRA" license="307796" swrid="5600199" athleteid="1901" externalid="307796">
              <RESULTS>
                <RESULT eventid="1061" points="360" swimtime="00:11:10.76" resultid="1902" heatid="1975" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="150" swimtime="00:01:53.49" />
                    <SPLIT distance="200" swimtime="00:02:34.22" />
                    <SPLIT distance="250" swimtime="00:03:15.35" />
                    <SPLIT distance="300" swimtime="00:03:58.32" />
                    <SPLIT distance="350" swimtime="00:04:41.29" />
                    <SPLIT distance="400" swimtime="00:05:24.67" />
                    <SPLIT distance="450" swimtime="00:06:07.57" />
                    <SPLIT distance="500" swimtime="00:06:50.46" />
                    <SPLIT distance="550" swimtime="00:07:33.65" />
                    <SPLIT distance="600" swimtime="00:08:17.55" />
                    <SPLIT distance="650" swimtime="00:09:02.04" />
                    <SPLIT distance="700" swimtime="00:09:44.65" />
                    <SPLIT distance="750" swimtime="00:10:27.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="423" swimtime="00:05:08.06" resultid="1903" heatid="2001" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                    <SPLIT distance="100" swimtime="00:01:12.70" />
                    <SPLIT distance="150" swimtime="00:01:51.65" />
                    <SPLIT distance="200" swimtime="00:02:31.10" />
                    <SPLIT distance="250" swimtime="00:03:10.29" />
                    <SPLIT distance="300" swimtime="00:03:50.00" />
                    <SPLIT distance="350" swimtime="00:04:29.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="363" swimtime="00:01:16.91" resultid="1904" heatid="2031" lane="8" entrytime="00:01:17.73" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3701" nation="BRA" region="PR" clubid="1512" name="Colégio Estadual Prof. Lysímaco Da Costa, Curitiba" shortname="Ctba-Lysímaco,Ce">
          <ATHLETES>
            <ATHLETE firstname="Marina" lastname="Heloisa Souza" birthdate="2007-01-15" gender="F" nation="BRA" license="336615" swrid="5600184" athleteid="1513" externalid="336615">
              <RESULTS>
                <RESULT eventid="1085" status="DNS" swimtime="00:00:00.00" resultid="1514" heatid="1990" lane="4" entrytime="00:01:00.05" entrycourse="SCM" />
                <RESULT eventid="1111" status="DNS" swimtime="00:00:00.00" resultid="1515" heatid="2002" lane="4" entrytime="00:04:32.60" entrycourse="SCM" />
                <RESULT eventid="1127" status="DNS" swimtime="00:00:00.00" resultid="1516" heatid="2009" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="8869" nation="BRA" region="PR" clubid="1700" name="Colégio Educação Dinâmica, Foz Do Iguaçu" shortname="Fozi-Dinâmica,C">
          <ATHLETES>
            <ATHLETE firstname="Vitor" lastname="Otremba Rouver" birthdate="2007-04-25" gender="M" nation="BRA" license="342152" swrid="5596919" athleteid="1701" externalid="342152">
              <RESULTS>
                <RESULT eventid="1081" points="474" swimtime="00:00:57.50" resultid="1702" heatid="1987" lane="7" entrytime="00:00:56.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="438" swimtime="00:00:26.53" resultid="1703" heatid="2017" lane="8" entrytime="00:00:25.96" entrycourse="SCM" />
                <RESULT eventid="1187" points="430" swimtime="00:00:28.81" resultid="1704" heatid="2041" lane="3" entrytime="00:00:27.44" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13383" nation="BRA" region="PR" clubid="1295" name="Colégio Bom Jesus Água Verde, Curitiba" shortname="Ctba-Bj Água Verde,C">
          <ATHLETES>
            <ATHLETE firstname="Isadora" lastname="Muller" birthdate="2009-10-10" gender="F" nation="BRA" license="376952" swrid="5600221" athleteid="1296" externalid="376952">
              <RESULTS>
                <RESULT eventid="1101" points="436" swimtime="00:00:37.40" resultid="1297" heatid="1998" lane="3" entrytime="00:00:37.42" entrycourse="SCM" />
                <RESULT eventid="1111" points="403" swimtime="00:05:12.94" resultid="1298" heatid="2002" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:12.76" />
                    <SPLIT distance="150" swimtime="00:01:51.82" />
                    <SPLIT distance="200" swimtime="00:02:31.51" />
                    <SPLIT distance="250" swimtime="00:03:11.64" />
                    <SPLIT distance="300" swimtime="00:03:52.10" />
                    <SPLIT distance="350" swimtime="00:04:32.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="453" swimtime="00:01:21.15" resultid="1299" heatid="2042" lane="3" entrytime="00:01:21.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16665" nation="BRA" region="PR" clubid="1830" name="Centro Estadual De Educação Profiss., Ponta Grossa" shortname="Pgro-Ceep,Ce">
          <ATHLETES>
            <ATHLETE firstname="Yago" lastname="Vallentin Cadene Dos Santos" birthdate="2009-10-19" gender="M" nation="BRA" license="V414499" athleteid="1831" externalid="V414499">
              <RESULTS>
                <RESULT eventid="1131" points="157" swimtime="00:00:37.33" resultid="1832" heatid="2013" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="10601" nation="BRA" region="PR" clubid="1630" name="Centro Estadual De Educação Profiss., Cascavel" shortname="Cvel-Ceep,Ce">
          <ATHLETES>
            <ATHLETE firstname="Juan" lastname="Balduíno" birthdate="2009-06-24" gender="M" nation="BRA" license="370764" swrid="5596870" athleteid="1631" externalid="370764">
              <RESULTS>
                <RESULT eventid="1073" points="365" reactiontime="+81" swimtime="00:00:30.91" resultid="1632" heatid="1979" lane="8" />
                <RESULT eventid="1139" points="378" swimtime="00:02:26.01" resultid="1633" heatid="2019" lane="4" entrytime="00:02:27.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                    <SPLIT distance="100" swimtime="00:01:10.00" />
                    <SPLIT distance="150" swimtime="00:01:48.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="392" swimtime="00:01:06.03" resultid="1634" heatid="2033" lane="7" entrytime="00:01:09.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="889" nation="BRA" region="PR" clubid="1392" name="Colégio Estadual Do Paraná, Curitiba" shortname="Ctba-Cep,Ce">
          <ATHLETES>
            <ATHLETE firstname="Pedro" lastname="De Castro Paiva Maciel" birthdate="2008-04-10" gender="M" nation="BRA" license="378333" swrid="5622275" athleteid="1393" externalid="378333">
              <RESULTS>
                <RESULT eventid="1081" points="426" swimtime="00:00:59.56" resultid="1394" heatid="1986" lane="3" entrytime="00:00:59.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="375" swimtime="00:01:06.21" resultid="1395" heatid="2021" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="424" swimtime="00:00:26.82" resultid="1396" heatid="2016" lane="7" entrytime="00:00:27.26" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wagner" lastname="Junior Cabral Gama" birthdate="2007-07-22" gender="M" nation="BRA" license="345334" swrid="5723027" athleteid="1397" externalid="345334">
              <RESULTS>
                <RESULT eventid="1073" points="339" swimtime="00:00:31.69" resultid="1398" heatid="1979" lane="2" />
                <RESULT eventid="1131" points="301" swimtime="00:00:30.08" resultid="1399" heatid="2014" lane="6" />
                <RESULT eventid="1171" points="290" swimtime="00:01:12.95" resultid="1400" heatid="2032" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mucke Buchmann" birthdate="2009-02-25" gender="F" nation="BRA" license="V414487" athleteid="1417" externalid="V414487">
              <RESULTS>
                <RESULT eventid="1077" points="113" swimtime="00:00:52.21" resultid="1418" heatid="1980" lane="5" />
                <RESULT eventid="1127" points="158" swimtime="00:00:42.34" resultid="1419" heatid="2008" lane="5" />
                <RESULT eventid="1167" points="94" swimtime="00:02:00.31" resultid="1420" heatid="2030" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Alface Cervelin" birthdate="2008-02-09" gender="M" nation="BRA" license="V414502" athleteid="1433" externalid="V414502">
              <RESULTS>
                <RESULT eventid="1073" points="172" swimtime="00:00:39.70" resultid="1434" heatid="1979" lane="7" />
                <RESULT eventid="1131" points="199" swimtime="00:00:34.53" resultid="1435" heatid="2014" lane="3" />
                <RESULT eventid="1171" status="DSQ" swimtime="00:01:33.17" resultid="1436" heatid="2032" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Bianchini De Quadros" birthdate="2009-08-04" gender="F" nation="BRA" license="V414488" athleteid="1421" externalid="V414488">
              <RESULTS>
                <RESULT eventid="1101" points="124" swimtime="00:00:56.84" resultid="1422" heatid="1997" lane="5" />
                <RESULT eventid="1127" points="190" swimtime="00:00:39.83" resultid="1423" heatid="2008" lane="3" />
                <RESULT eventid="1167" status="DSQ" swimtime="00:00:00.00" resultid="1424" heatid="2030" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Vitor Da Silva" birthdate="2008-10-23" gender="M" nation="BRA" license="V414503" athleteid="1437" externalid="V414503">
              <RESULTS>
                <RESULT eventid="1081" points="165" swimtime="00:01:21.60" resultid="1438" heatid="1984" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="121" swimtime="00:03:41.61" resultid="1439" heatid="1976" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                    <SPLIT distance="100" swimtime="00:01:35.48" />
                    <SPLIT distance="150" swimtime="00:02:48.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="170" swimtime="00:00:39.24" resultid="1440" heatid="2040" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Rodrigues Galvao" birthdate="2007-04-19" gender="M" nation="BRA" license="376586" swrid="5600247" athleteid="1401" externalid="376586">
              <RESULTS>
                <RESULT eventid="1089" status="DSQ" swimtime="00:02:32.38" resultid="1402" heatid="1991" lane="7" entrytime="00:02:31.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.23" />
                    <SPLIT distance="100" swimtime="00:01:07.27" />
                    <SPLIT distance="150" swimtime="00:01:48.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="423" swimtime="00:01:03.62" resultid="1403" heatid="2023" lane="2" entrytime="00:01:02.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="1404" heatid="2041" lane="5" entrytime="00:00:27.06" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Bilecki" birthdate="2007-05-28" gender="M" nation="BRA" license="406726" swrid="5717247" athleteid="1409" externalid="406726">
              <RESULTS>
                <RESULT eventid="1081" status="DNS" swimtime="00:00:00.00" resultid="1410" heatid="1985" lane="6" entrytime="00:01:06.54" entrycourse="SCM" />
                <RESULT eventid="1147" status="DNS" swimtime="00:00:00.00" resultid="1411" heatid="2022" lane="6" entrytime="00:01:18.82" entrycourse="SCM" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="1412" heatid="2040" lane="3" entrytime="00:00:33.15" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Torres Oliveira" birthdate="2008-04-10" gender="M" nation="BRA" license="400274" swrid="5653303" athleteid="1405" externalid="400274">
              <RESULTS>
                <RESULT eventid="1065" points="235" swimtime="00:02:57.62" resultid="1406" heatid="1976" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:21.78" />
                    <SPLIT distance="150" swimtime="00:02:13.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="210" swimtime="00:03:21.95" resultid="1407" heatid="2006" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.08" />
                    <SPLIT distance="100" swimtime="00:01:30.24" />
                    <SPLIT distance="150" swimtime="00:02:26.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="248" swimtime="00:01:27.92" resultid="1408" heatid="2044" lane="6" entrytime="00:01:27.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="Rosa Rodrigues Da Silva" birthdate="2009-03-03" gender="F" nation="BRA" license="V414489" athleteid="1425" externalid="V414489">
              <RESULTS>
                <RESULT eventid="1085" points="134" swimtime="00:01:38.15" resultid="1426" heatid="1988" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1069" status="DNS" swimtime="00:00:00.00" resultid="1427" heatid="1977" lane="3" />
                <RESULT eventid="1127" points="242" swimtime="00:00:36.76" resultid="1428" heatid="2008" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Carolina Barbosa De Oliveira" birthdate="2009-01-19" gender="F" nation="BRA" license="V414486" athleteid="1413" externalid="V414486">
              <RESULTS>
                <RESULT eventid="1085" points="153" swimtime="00:01:33.92" resultid="1414" heatid="1989" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="128" swimtime="00:00:50.07" resultid="1415" heatid="1981" lane="7" />
                <RESULT eventid="1175" points="98" swimtime="00:03:58.72" resultid="1416" heatid="2034" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.27" />
                    <SPLIT distance="100" swimtime="00:01:55.83" />
                    <SPLIT distance="150" swimtime="00:03:03.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Alixandrini" birthdate="2009-02-20" gender="F" nation="BRA" license="V414490" athleteid="1429" externalid="V414490">
              <RESULTS>
                <RESULT eventid="1085" points="96" swimtime="00:01:49.40" resultid="1430" heatid="1988" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="65" swimtime="00:01:02.56" resultid="1431" heatid="1980" lane="4" />
                <RESULT eventid="1167" status="DNS" swimtime="00:00:00.00" resultid="1432" heatid="2030" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CTBA-CEP,CE &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1161" points="424" swimtime="00:01:48.85" resultid="1443" heatid="2027" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.33" />
                    <SPLIT distance="100" swimtime="00:00:56.30" />
                    <SPLIT distance="150" swimtime="00:01:22.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1393" number="1" />
                    <RELAYPOSITION athleteid="1405" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1397" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1401" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1203" points="285" swimtime="00:02:16.18" resultid="1444" heatid="2048" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.28" />
                    <SPLIT distance="150" swimtime="00:01:49.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1397" number="1" />
                    <RELAYPOSITION athleteid="1405" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1437" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1393" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="CTBA-CEP,CE &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1159" points="192" swimtime="00:02:40.07" resultid="1441" heatid="2026" lane="5">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:02.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1421" number="1" />
                    <RELAYPOSITION athleteid="1429" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1413" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1425" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1205" status="DSQ" swimtime="00:03:13.10" resultid="1442" heatid="2049" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.28" />
                    <SPLIT distance="100" swimtime="00:01:47.10" />
                    <SPLIT distance="150" swimtime="00:02:31.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1417" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="1421" number="2" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1425" number="3" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1413" number="4" reactiontime="0" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="CTBA-CEP,CE &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1109" points="226" swimtime="00:02:36.17" resultid="1445" heatid="2000" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:28.60" />
                    <SPLIT distance="150" swimtime="00:01:56.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1397" number="1" />
                    <RELAYPOSITION athleteid="1421" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1401" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1425" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="18922" nation="BRA" region="PR" clubid="1270" name="Colégio Estadual Antônio Lacerda Braga, Colombo" shortname="Colb-Antôniobraga,Ce">
          <ATHLETES>
            <ATHLETE firstname="Kethelyn" lastname="Ribeiro Rodrigues" birthdate="2009-04-24" gender="F" nation="BRA" license="367052" swrid="5600244" athleteid="1271" externalid="367052">
              <RESULTS>
                <RESULT eventid="1085" points="379" swimtime="00:01:09.43" resultid="1272" heatid="1990" lane="6" entrytime="00:01:07.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="266" swimtime="00:00:39.26" resultid="1273" heatid="1981" lane="4" entrytime="00:00:38.51" entrycourse="SCM" />
                <RESULT eventid="1127" points="365" swimtime="00:00:32.08" resultid="1274" heatid="2010" lane="5" entrytime="00:00:30.69" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6525" nation="BRA" region="PR" clubid="1655" name="Colégio Santa Maria, Cascavel" shortname="Cvel-Santa Maria, C">
          <ATHLETES>
            <ATHLETE firstname="Milena" lastname="Gamero Prado" birthdate="2007-05-16" gender="F" nation="BRA" license="305973" swrid="5596903" athleteid="1656" externalid="305973">
              <RESULTS>
                <RESULT eventid="1061" points="448" swimtime="00:10:23.52" resultid="1657" heatid="1975" lane="3" entrytime="00:10:12.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:10.28" />
                    <SPLIT distance="150" swimtime="00:01:48.30" />
                    <SPLIT distance="200" swimtime="00:02:27.43" />
                    <SPLIT distance="250" swimtime="00:03:07.01" />
                    <SPLIT distance="300" swimtime="00:03:46.20" />
                    <SPLIT distance="350" swimtime="00:04:26.09" />
                    <SPLIT distance="400" swimtime="00:05:06.08" />
                    <SPLIT distance="450" swimtime="00:05:44.32" />
                    <SPLIT distance="500" swimtime="00:06:23.46" />
                    <SPLIT distance="550" swimtime="00:07:02.32" />
                    <SPLIT distance="600" swimtime="00:07:41.26" />
                    <SPLIT distance="650" swimtime="00:08:20.00" />
                    <SPLIT distance="700" swimtime="00:09:00.18" />
                    <SPLIT distance="750" swimtime="00:09:41.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="467" swimtime="00:04:58.05" resultid="1658" heatid="2002" lane="6" entrytime="00:04:59.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:09.52" />
                    <SPLIT distance="150" swimtime="00:01:46.92" />
                    <SPLIT distance="200" swimtime="00:02:25.69" />
                    <SPLIT distance="250" swimtime="00:03:03.65" />
                    <SPLIT distance="300" swimtime="00:03:41.79" />
                    <SPLIT distance="350" swimtime="00:04:20.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" points="404" swimtime="00:20:28.07" resultid="1659" heatid="2047" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                    <SPLIT distance="100" swimtime="00:01:12.21" />
                    <SPLIT distance="150" swimtime="00:01:50.28" />
                    <SPLIT distance="200" swimtime="00:02:29.23" />
                    <SPLIT distance="250" swimtime="00:03:09.20" />
                    <SPLIT distance="300" swimtime="00:03:50.01" />
                    <SPLIT distance="350" swimtime="00:04:31.03" />
                    <SPLIT distance="400" swimtime="00:05:11.58" />
                    <SPLIT distance="450" swimtime="00:05:52.63" />
                    <SPLIT distance="500" swimtime="00:06:33.58" />
                    <SPLIT distance="550" swimtime="00:07:14.44" />
                    <SPLIT distance="600" swimtime="00:07:55.39" />
                    <SPLIT distance="650" swimtime="00:08:36.51" />
                    <SPLIT distance="700" swimtime="00:09:17.79" />
                    <SPLIT distance="750" swimtime="00:09:57.16" />
                    <SPLIT distance="800" swimtime="00:10:36.72" />
                    <SPLIT distance="850" swimtime="00:11:17.54" />
                    <SPLIT distance="900" swimtime="00:11:59.77" />
                    <SPLIT distance="950" swimtime="00:12:41.45" />
                    <SPLIT distance="1000" swimtime="00:13:23.08" />
                    <SPLIT distance="1050" swimtime="00:14:01.23" />
                    <SPLIT distance="1100" swimtime="00:14:40.80" />
                    <SPLIT distance="1150" swimtime="00:15:20.87" />
                    <SPLIT distance="1200" swimtime="00:16:04.72" />
                    <SPLIT distance="1250" swimtime="00:16:48.27" />
                    <SPLIT distance="1300" swimtime="00:17:31.81" />
                    <SPLIT distance="1350" swimtime="00:18:15.63" />
                    <SPLIT distance="1400" swimtime="00:18:59.22" />
                    <SPLIT distance="1450" swimtime="00:19:43.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luann" lastname="Miguel Mazur" birthdate="2007-01-10" gender="M" nation="BRA" license="365682" swrid="5596915" athleteid="1664" externalid="365682">
              <RESULTS>
                <RESULT eventid="1123" points="451" swimtime="00:02:36.65" resultid="1665" heatid="2007" lane="6" entrytime="00:02:34.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.60" />
                    <SPLIT distance="100" swimtime="00:01:14.86" />
                    <SPLIT distance="150" swimtime="00:01:55.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="465" swimtime="00:05:02.95" resultid="1666" heatid="2025" lane="6" entrytime="00:04:58.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                    <SPLIT distance="100" swimtime="00:01:09.69" />
                    <SPLIT distance="150" swimtime="00:01:49.85" />
                    <SPLIT distance="200" swimtime="00:02:29.13" />
                    <SPLIT distance="250" swimtime="00:03:10.87" />
                    <SPLIT distance="300" swimtime="00:03:53.19" />
                    <SPLIT distance="350" swimtime="00:04:28.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="429" swimtime="00:01:13.29" resultid="1667" heatid="2045" lane="6" entrytime="00:01:10.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Rinaldini" birthdate="2009-04-09" gender="M" nation="BRA" license="348289" swrid="5596932" athleteid="1660" externalid="348289">
              <RESULTS>
                <RESULT eventid="1105" points="572" swimtime="00:16:59.77" resultid="1661" heatid="1999" lane="4" entrytime="00:17:16.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                    <SPLIT distance="150" swimtime="00:01:37.96" />
                    <SPLIT distance="200" swimtime="00:02:11.95" />
                    <SPLIT distance="250" swimtime="00:02:45.77" />
                    <SPLIT distance="300" swimtime="00:03:19.82" />
                    <SPLIT distance="350" swimtime="00:03:54.03" />
                    <SPLIT distance="400" swimtime="00:04:28.53" />
                    <SPLIT distance="450" swimtime="00:05:02.93" />
                    <SPLIT distance="500" swimtime="00:05:37.17" />
                    <SPLIT distance="550" swimtime="00:06:11.20" />
                    <SPLIT distance="600" swimtime="00:06:45.59" />
                    <SPLIT distance="650" swimtime="00:07:19.44" />
                    <SPLIT distance="700" swimtime="00:07:53.79" />
                    <SPLIT distance="750" swimtime="00:08:28.03" />
                    <SPLIT distance="800" swimtime="00:09:02.21" />
                    <SPLIT distance="850" swimtime="00:09:36.65" />
                    <SPLIT distance="900" swimtime="00:10:11.12" />
                    <SPLIT distance="950" swimtime="00:10:45.18" />
                    <SPLIT distance="1000" swimtime="00:11:19.45" />
                    <SPLIT distance="1050" swimtime="00:11:53.06" />
                    <SPLIT distance="1100" swimtime="00:12:27.29" />
                    <SPLIT distance="1150" swimtime="00:13:01.36" />
                    <SPLIT distance="1200" swimtime="00:13:35.36" />
                    <SPLIT distance="1250" swimtime="00:14:09.87" />
                    <SPLIT distance="1300" swimtime="00:14:43.79" />
                    <SPLIT distance="1350" swimtime="00:15:18.30" />
                    <SPLIT distance="1400" swimtime="00:15:52.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="534" swimtime="00:04:21.48" resultid="1662" heatid="2004" lane="3" entrytime="00:04:18.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.41" />
                    <SPLIT distance="100" swimtime="00:01:00.96" />
                    <SPLIT distance="150" swimtime="00:01:33.55" />
                    <SPLIT distance="200" swimtime="00:02:06.95" />
                    <SPLIT distance="250" swimtime="00:02:40.79" />
                    <SPLIT distance="300" swimtime="00:03:14.67" />
                    <SPLIT distance="350" swimtime="00:03:48.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="567" swimtime="00:08:55.44" resultid="1663" heatid="2029" lane="5" entrytime="00:09:00.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.67" />
                    <SPLIT distance="100" swimtime="00:01:03.54" />
                    <SPLIT distance="150" swimtime="00:01:36.96" />
                    <SPLIT distance="200" swimtime="00:02:10.39" />
                    <SPLIT distance="250" swimtime="00:02:44.33" />
                    <SPLIT distance="300" swimtime="00:03:18.21" />
                    <SPLIT distance="350" swimtime="00:03:52.14" />
                    <SPLIT distance="400" swimtime="00:04:25.41" />
                    <SPLIT distance="450" swimtime="00:04:59.39" />
                    <SPLIT distance="500" swimtime="00:05:32.95" />
                    <SPLIT distance="550" swimtime="00:06:07.09" />
                    <SPLIT distance="600" swimtime="00:06:41.27" />
                    <SPLIT distance="650" swimtime="00:07:15.14" />
                    <SPLIT distance="700" swimtime="00:07:49.00" />
                    <SPLIT distance="750" swimtime="00:08:22.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Do Prado Martins" birthdate="2008-10-17" gender="F" nation="BRA" license="369419" swrid="5596893" athleteid="1668" externalid="369419">
              <RESULTS>
                <RESULT eventid="1069" status="DSQ" swimtime="00:02:33.34" resultid="1669" heatid="1977" lane="5" entrytime="00:02:36.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:12.44" />
                    <SPLIT distance="150" swimtime="00:01:56.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="458" swimtime="00:02:54.47" resultid="1670" heatid="2005" lane="4" entrytime="00:02:49.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                    <SPLIT distance="100" swimtime="00:01:23.12" />
                    <SPLIT distance="150" swimtime="00:02:07.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="469" swimtime="00:05:33.16" resultid="1671" heatid="2024" lane="4" entrytime="00:05:29.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:01:16.56" />
                    <SPLIT distance="150" swimtime="00:01:59.38" />
                    <SPLIT distance="200" swimtime="00:02:41.48" />
                    <SPLIT distance="250" swimtime="00:03:28.15" />
                    <SPLIT distance="300" swimtime="00:04:15.72" />
                    <SPLIT distance="350" swimtime="00:04:54.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="CVEL-SANTA MARIA, C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1109" points="401" swimtime="00:02:09.03" resultid="1672" heatid="2000" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:05.92" />
                    <SPLIT distance="150" swimtime="00:01:39.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1660" number="1" />
                    <RELAYPOSITION athleteid="1664" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1656" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1668" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="9878" nation="BRA" region="PR" clubid="1650" name="Colégio Estadual Marilis Faria Pirotelli, Cascavel" shortname="Cvel-Marilis Piro,Ce">
          <ATHLETES>
            <ATHLETE firstname="Heloisa" lastname="Souza Garute Da Silva" birthdate="2009-01-07" gender="F" nation="BRA" license="329307" swrid="5596940" athleteid="1651" externalid="329307">
              <RESULTS>
                <RESULT eventid="1069" points="447" swimtime="00:02:39.35" resultid="1652" heatid="1977" lane="4" entrytime="00:02:32.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.46" />
                    <SPLIT distance="100" swimtime="00:01:17.74" />
                    <SPLIT distance="150" swimtime="00:02:03.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="407" swimtime="00:02:40.49" resultid="1653" heatid="2018" lane="4" entrytime="00:02:40.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                    <SPLIT distance="100" swimtime="00:01:18.45" />
                    <SPLIT distance="150" swimtime="00:01:59.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="386" swimtime="00:01:15.34" resultid="1654" heatid="2031" lane="2" entrytime="00:01:13.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2654" nation="BRA" region="PR" clubid="1803" name="Colégio Platão, Maringá" shortname="Mrga-Platão,C">
          <ATHLETES>
            <ATHLETE firstname="Beatriz" lastname="Passafaro" birthdate="2009-02-01" gender="F" nation="BRA" license="370673" swrid="5603885" athleteid="1804" externalid="370673">
              <RESULTS>
                <RESULT eventid="1085" points="330" swimtime="00:01:12.67" resultid="1805" heatid="1990" lane="7" entrytime="00:01:09.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" status="DSQ" swimtime="00:00:31.88" resultid="1806" heatid="2010" lane="3" entrytime="00:00:30.77" entrycourse="SCM" />
                <RESULT eventid="1183" status="DSQ" swimtime="00:00:34.64" resultid="1807" heatid="2038" lane="2" entrytime="00:00:34.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13438" nation="BRA" region="PR" clubid="1600" name="Colégio Santo Anjo, Curitiba" shortname="Ctba-Santo Anjo,C">
          <ATHLETES>
            <ATHLETE firstname="Camila" lastname="Duarte De Almeida" birthdate="2009-11-26" gender="F" nation="BRA" license="378819" swrid="5600152" athleteid="1601" externalid="378819">
              <RESULTS>
                <RESULT eventid="1085" points="434" swimtime="00:01:06.35" resultid="1602" heatid="1990" lane="2" entrytime="00:01:07.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="431" swimtime="00:00:30.34" resultid="1603" heatid="2011" lane="8" entrytime="00:00:30.44" entrycourse="SCM" />
                <RESULT eventid="1183" points="364" swimtime="00:00:34.13" resultid="1604" heatid="2038" lane="6" entrytime="00:00:34.28" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18920" nation="BRA" region="PR" clubid="1881" name="Instituto Federal Do Paraná, Pinhais" shortname="Pinh-Ifpr">
          <ATHLETES>
            <ATHLETE firstname="Benito" lastname="Alves Sant&apos;Ana" birthdate="2009-06-01" gender="M" nation="BRA" license="376585" swrid="5351951" athleteid="1882" externalid="376585">
              <RESULTS>
                <RESULT eventid="1065" points="430" swimtime="00:02:25.14" resultid="1883" heatid="1976" lane="5" entrytime="00:02:28.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:01:08.19" />
                    <SPLIT distance="150" swimtime="00:01:52.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="501" swimtime="00:04:27.07" resultid="1884" heatid="2004" lane="6" entrytime="00:04:32.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="100" swimtime="00:01:03.54" />
                    <SPLIT distance="150" swimtime="00:01:37.87" />
                    <SPLIT distance="200" swimtime="00:02:11.80" />
                    <SPLIT distance="250" swimtime="00:02:46.07" />
                    <SPLIT distance="300" swimtime="00:03:21.18" />
                    <SPLIT distance="350" swimtime="00:03:54.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="536" swimtime="00:09:05.63" resultid="1885" heatid="2028" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.62" />
                    <SPLIT distance="100" swimtime="00:01:03.60" />
                    <SPLIT distance="150" swimtime="00:01:37.78" />
                    <SPLIT distance="200" swimtime="00:02:12.67" />
                    <SPLIT distance="250" swimtime="00:02:46.38" />
                    <SPLIT distance="300" swimtime="00:03:19.81" />
                    <SPLIT distance="350" swimtime="00:03:54.45" />
                    <SPLIT distance="400" swimtime="00:04:29.26" />
                    <SPLIT distance="450" swimtime="00:05:04.34" />
                    <SPLIT distance="500" swimtime="00:05:39.60" />
                    <SPLIT distance="550" swimtime="00:06:15.13" />
                    <SPLIT distance="600" swimtime="00:06:50.36" />
                    <SPLIT distance="650" swimtime="00:07:25.50" />
                    <SPLIT distance="700" swimtime="00:08:00.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6506" nation="BRA" region="PR" clubid="1255" name="Colégio Adventista De Campo Mourão" shortname="Cmou-Adventista,C">
          <ATHLETES>
            <ATHLETE firstname="Arthur" lastname="Batinga Ponchielli" birthdate="2007-01-18" gender="M" nation="BRA" license="378461" swrid="5251143" athleteid="1256" externalid="378461">
              <RESULTS>
                <RESULT eventid="1073" points="249" swimtime="00:00:35.13" resultid="1257" heatid="1979" lane="3" entrytime="00:00:33.52" entrycourse="SCM" />
                <RESULT eventid="1131" points="287" swimtime="00:00:30.55" resultid="1258" heatid="2015" lane="7" entrytime="00:00:30.02" entrycourse="SCM" />
                <RESULT eventid="1171" points="218" swimtime="00:01:20.24" resultid="1259" heatid="2032" lane="4" entrytime="00:01:18.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4573" nation="BRA" region="PR" clubid="1705" name="Instituto Federal Do Paraná, Foz Do Iguaçu" shortname="Fozi-Ifpr">
          <ATHLETES>
            <ATHLETE firstname="Christopher" lastname="De Araujo" birthdate="2008-08-09" gender="M" nation="BRA" license="366376" swrid="5596884" athleteid="1706" externalid="366376" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1105" points="491" swimtime="00:17:52.91" resultid="1707" heatid="1999" lane="5" entrytime="00:17:32.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:05.11" />
                    <SPLIT distance="150" swimtime="00:01:38.63" />
                    <SPLIT distance="200" swimtime="00:02:12.91" />
                    <SPLIT distance="250" swimtime="00:02:46.77" />
                    <SPLIT distance="300" swimtime="00:03:21.94" />
                    <SPLIT distance="350" swimtime="00:03:57.43" />
                    <SPLIT distance="400" swimtime="00:04:33.26" />
                    <SPLIT distance="450" swimtime="00:05:09.25" />
                    <SPLIT distance="500" swimtime="00:05:44.95" />
                    <SPLIT distance="550" swimtime="00:06:20.77" />
                    <SPLIT distance="600" swimtime="00:06:56.94" />
                    <SPLIT distance="650" swimtime="00:07:33.11" />
                    <SPLIT distance="700" swimtime="00:08:08.96" />
                    <SPLIT distance="750" swimtime="00:08:45.22" />
                    <SPLIT distance="800" swimtime="00:09:21.55" />
                    <SPLIT distance="850" swimtime="00:09:58.34" />
                    <SPLIT distance="900" swimtime="00:10:34.82" />
                    <SPLIT distance="950" swimtime="00:11:11.43" />
                    <SPLIT distance="1000" swimtime="00:11:48.45" />
                    <SPLIT distance="1050" swimtime="00:12:25.62" />
                    <SPLIT distance="1100" swimtime="00:13:02.11" />
                    <SPLIT distance="1150" swimtime="00:13:39.25" />
                    <SPLIT distance="1200" swimtime="00:14:15.44" />
                    <SPLIT distance="1250" swimtime="00:14:52.27" />
                    <SPLIT distance="1300" swimtime="00:15:28.73" />
                    <SPLIT distance="1350" swimtime="00:16:05.58" />
                    <SPLIT distance="1400" swimtime="00:16:42.24" />
                    <SPLIT distance="1450" swimtime="00:17:18.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="455" swimtime="00:05:05.24" resultid="1708" heatid="2025" lane="3" entrytime="00:04:53.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:08.16" />
                    <SPLIT distance="150" swimtime="00:01:48.65" />
                    <SPLIT distance="200" swimtime="00:02:28.90" />
                    <SPLIT distance="250" swimtime="00:03:13.61" />
                    <SPLIT distance="300" swimtime="00:03:58.11" />
                    <SPLIT distance="350" swimtime="00:04:32.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="529" swimtime="00:02:02.81" resultid="1709" heatid="2035" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.73" />
                    <SPLIT distance="100" swimtime="00:00:58.68" />
                    <SPLIT distance="150" swimtime="00:01:30.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18918" nation="BRA" region="PR" clubid="1808" name="Colégio Pro, Maringá" shortname="Mrga-Pro,C">
          <ATHLETES>
            <ATHLETE firstname="Felipe" lastname="Berto" birthdate="2008-10-22" gender="M" nation="BRA" license="378342" swrid="5312223" athleteid="1809" externalid="378342">
              <RESULTS>
                <RESULT eventid="1081" status="DNS" swimtime="00:00:00.00" resultid="1810" heatid="1985" lane="3" entrytime="00:01:06.32" entrycourse="SCM" />
                <RESULT eventid="1123" status="DNS" swimtime="00:00:00.00" resultid="1811" heatid="2006" lane="4" entrytime="00:02:43.26" entrycourse="SCM" />
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="1812" heatid="2044" lane="5" entrytime="00:01:17.98" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11552" nation="BRA" region="PR" clubid="1635" name="Colégio Fag, Cascavel" shortname="Cvel-Fag,C">
          <ATHLETES>
            <ATHLETE firstname="Felipe" lastname="Mariotti De Castro" birthdate="2008-06-27" gender="M" nation="BRA" license="329200" swrid="5596912" athleteid="1636" externalid="329200">
              <RESULTS>
                <RESULT eventid="1089" points="540" swimtime="00:02:11.18" resultid="1637" heatid="1991" lane="4" entrytime="00:02:09.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.71" />
                    <SPLIT distance="100" swimtime="00:01:02.40" />
                    <SPLIT distance="150" swimtime="00:01:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="542" swimtime="00:04:47.90" resultid="1638" heatid="2025" lane="4" entrytime="00:04:36.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                    <SPLIT distance="100" swimtime="00:01:04.52" />
                    <SPLIT distance="150" swimtime="00:01:41.72" />
                    <SPLIT distance="200" swimtime="00:02:18.50" />
                    <SPLIT distance="250" swimtime="00:03:00.80" />
                    <SPLIT distance="300" swimtime="00:03:42.99" />
                    <SPLIT distance="350" swimtime="00:04:16.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="613" swimtime="00:08:41.72" resultid="1639" heatid="2029" lane="4" entrytime="00:08:38.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                    <SPLIT distance="100" swimtime="00:01:01.79" />
                    <SPLIT distance="150" swimtime="00:01:34.26" />
                    <SPLIT distance="200" swimtime="00:02:06.89" />
                    <SPLIT distance="250" swimtime="00:02:39.59" />
                    <SPLIT distance="300" swimtime="00:03:12.77" />
                    <SPLIT distance="350" swimtime="00:03:46.52" />
                    <SPLIT distance="400" swimtime="00:04:20.60" />
                    <SPLIT distance="450" swimtime="00:04:52.40" />
                    <SPLIT distance="500" swimtime="00:05:25.52" />
                    <SPLIT distance="550" swimtime="00:05:58.72" />
                    <SPLIT distance="600" swimtime="00:06:32.08" />
                    <SPLIT distance="650" swimtime="00:07:05.10" />
                    <SPLIT distance="700" swimtime="00:07:38.58" />
                    <SPLIT distance="750" swimtime="00:08:11.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15542" nation="BRA" region="PR" clubid="1280" name="Colégio Estadual Ângelo Gusso, Curitiba" shortname="Ctba-Ângelo Gusso,Ce">
          <ATHLETES>
            <ATHLETE firstname="Fabio" lastname="C Burak" birthdate="2009-08-29" gender="M" nation="BRA" license="343297" swrid="5600126" athleteid="1281" externalid="343297">
              <RESULTS>
                <RESULT eventid="1065" points="407" swimtime="00:02:27.92" resultid="1282" heatid="1976" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                    <SPLIT distance="100" swimtime="00:01:12.58" />
                    <SPLIT distance="150" swimtime="00:01:53.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="385" swimtime="00:00:34.27" resultid="1283" heatid="1994" lane="4" />
                <RESULT eventid="1195" points="419" swimtime="00:01:13.82" resultid="1284" heatid="2045" lane="7" entrytime="00:01:12.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2670" nation="BRA" region="PR" clubid="1517" name="Colégio Marista Paranaense, Curitiba" shortname="Ctba-Marista Pr,C">
          <ATHLETES>
            <ATHLETE firstname="Pedro" lastname="Sachser Rocha" birthdate="2008-07-09" gender="M" nation="BRA" license="330072" swrid="5600254" athleteid="1522" externalid="330072">
              <RESULTS>
                <RESULT eventid="1065" status="DNS" swimtime="00:00:00.00" resultid="1523" heatid="1976" lane="3" />
                <RESULT eventid="1147" status="DNS" swimtime="00:00:00.00" resultid="1524" heatid="2021" lane="5" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="1525" heatid="2041" lane="4" entrytime="00:00:26.95" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo" lastname="Gabriel Nascimento" birthdate="2008-11-14" gender="M" nation="BRA" license="348028" swrid="5600171" athleteid="1526" externalid="348028" level="BIG BUM">
              <RESULTS>
                <RESULT eventid="1097" points="319" swimtime="00:00:36.48" resultid="1527" heatid="1994" lane="7" />
                <RESULT eventid="1147" points="372" swimtime="00:01:06.43" resultid="1528" heatid="2023" lane="8" entrytime="00:01:04.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="426" swimtime="00:00:28.89" resultid="1529" heatid="2041" lane="2" entrytime="00:00:28.27" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Moreira Segadaes" birthdate="2008-05-15" gender="M" nation="BRA" license="331574" swrid="5600220" athleteid="1518" externalid="331574">
              <RESULTS>
                <RESULT eventid="1097" points="477" swimtime="00:00:31.92" resultid="1519" heatid="1996" lane="3" entrytime="00:00:30.80" entrycourse="SCM" />
                <RESULT eventid="1123" status="DSQ" swimtime="00:02:32.36" resultid="1520" heatid="2007" lane="2" entrytime="00:02:36.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:11.00" />
                    <SPLIT distance="150" swimtime="00:01:51.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="504" swimtime="00:01:09.44" resultid="1521" heatid="2045" lane="5" entrytime="00:01:07.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15563" nation="BRA" region="PR" clubid="1724" name="CCM Manoel Ribas, Guarapuava" shortname="Grpa-Manoelribas,CCM">
          <ATHLETES>
            <ATHLETE firstname="Nilton" lastname="Cesar Medeiros Junior" birthdate="2008-01-14" gender="M" nation="BRA" license="V371155" athleteid="1725" externalid="V371155">
              <RESULTS>
                <RESULT eventid="1115" status="DNS" swimtime="00:00:00.00" resultid="1726" heatid="2003" lane="5" />
                <RESULT eventid="1131" status="DNS" swimtime="00:00:00.00" resultid="1727" heatid="2012" lane="5" />
                <RESULT eventid="1187" status="DNS" swimtime="00:00:00.00" resultid="1728" heatid="2039" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6523" nation="BRA" region="PR" clubid="1208" name="Colégio Nossa Senhora Da Glória, Apucarana" shortname="Apuc-N.Sra.Glória,C">
          <ATHLETES>
            <ATHLETE firstname="Gustavo" lastname="Brum Nepomuceno De Souza" birthdate="2007-12-11" gender="M" nation="BRA" license="V414513" athleteid="1209" externalid="V414513">
              <RESULTS>
                <RESULT eventid="1081" status="DNS" swimtime="00:00:00.00" resultid="1210" heatid="1983" lane="5" />
                <RESULT eventid="1131" points="297" swimtime="00:00:30.20" resultid="1211" heatid="2013" lane="6" />
                <RESULT eventid="1187" points="209" swimtime="00:00:36.63" resultid="1212" heatid="2039" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="319" nation="BRA" region="PR" clubid="1213" name="Colégio São José, Apucarana" shortname="Apuc-São José,C">
          <ATHLETES>
            <ATHLETE firstname="Thiago" lastname="Henrique Ferreira" birthdate="2009-07-13" gender="M" nation="BRA" license="V383399" athleteid="1217" externalid="V383399">
              <RESULTS>
                <RESULT eventid="1073" points="142" swimtime="00:00:42.34" resultid="1218" heatid="1979" lane="1" />
                <RESULT eventid="1131" points="221" swimtime="00:00:33.31" resultid="1219" heatid="2012" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Gabriel Galhardo" birthdate="2009-10-23" gender="M" nation="BRA" license="V414506" athleteid="1220" externalid="V414506">
              <RESULTS>
                <RESULT eventid="1097" status="DSQ" swimtime="00:00:56.37" resultid="1221" heatid="1995" lane="1" />
                <RESULT eventid="1131" points="133" swimtime="00:00:39.49" resultid="1222" heatid="2013" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Henrique Ferreira" birthdate="2008-10-01" gender="M" nation="BRA" license="V383397" athleteid="1214" externalid="V383397">
              <RESULTS>
                <RESULT eventid="1097" status="DSQ" swimtime="00:00:48.95" resultid="1215" heatid="1993" lane="3" />
                <RESULT eventid="1131" points="220" swimtime="00:00:33.38" resultid="1216" heatid="2012" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Santos Miquelin" birthdate="2009-09-22" gender="M" nation="BRA" license="V414509" athleteid="1226" externalid="V414509">
              <RESULTS>
                <RESULT eventid="1097" points="112" swimtime="00:00:51.76" resultid="1227" heatid="1995" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heitor Souza Telles" lastname="Proença" birthdate="2009-06-10" gender="M" nation="BRA" license="V414558" athleteid="2061" externalid="V414558" />
            <ATHLETE firstname="Ian" lastname="Da Silva Batista" birthdate="2009-12-22" gender="M" nation="BRA" license="V414507" athleteid="1223" externalid="V414507">
              <RESULTS>
                <RESULT eventid="1097" status="DSQ" swimtime="00:00:54.00" resultid="1224" heatid="1995" lane="8" />
                <RESULT eventid="1131" points="138" swimtime="00:00:38.97" resultid="1225" heatid="2014" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="APUC-C SAO JOSE &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1161" points="196" swimtime="00:02:20.64" resultid="1228" heatid="2027" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:01:13.28" />
                    <SPLIT distance="150" swimtime="00:01:47.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1217" number="1" />
                    <RELAYPOSITION athleteid="1223" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1214" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="2061" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="2649" nation="BRA" region="PR" clubid="1905" name="Colégio Estadual Presidente Castelo Branco, Toledo" shortname="Tole-Caste.Branco,Ce">
          <ATHLETES>
            <ATHLETE firstname="Pedro" lastname="Henrique Dell Agnolo Da Silva" birthdate="2009-12-18" gender="M" nation="BRA" license="V414500" athleteid="1906" externalid="V414500">
              <RESULTS>
                <RESULT eventid="1081" points="187" swimtime="00:01:18.30" resultid="1907" heatid="1985" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" status="DSQ" swimtime="00:01:43.86" resultid="1908" heatid="2021" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alisson" lastname="Bratz Frana" birthdate="2009-10-15" gender="M" nation="BRA" license="V414501" athleteid="1909" externalid="V414501">
              <RESULTS>
                <RESULT eventid="1097" points="154" swimtime="00:00:46.49" resultid="1910" heatid="1993" lane="5" />
                <RESULT eventid="1131" points="248" swimtime="00:00:32.06" resultid="1911" heatid="2013" lane="3" />
                <RESULT eventid="1187" status="DSQ" swimtime="00:00:39.58" resultid="1912" heatid="2040" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15583" nation="BRA" region="PR" clubid="1581" name="Colégio Positivo Boa Vista, Curitiba" shortname="Ctba-Posi. B.Vista,C">
          <ATHLETES>
            <ATHLETE firstname="Pedro" lastname="Giuseppe Bulla Lanaro" birthdate="2007-05-22" gender="M" nation="BRA" license="331630" swrid="5600174" athleteid="1582" externalid="331630">
              <RESULTS>
                <RESULT eventid="1081" points="552" swimtime="00:00:54.64" resultid="1583" heatid="1987" lane="4" entrytime="00:00:53.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="596" swimtime="00:04:12.17" resultid="1584" heatid="2004" lane="4" entrytime="00:04:11.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.11" />
                    <SPLIT distance="100" swimtime="00:00:59.44" />
                    <SPLIT distance="150" swimtime="00:01:31.29" />
                    <SPLIT distance="200" swimtime="00:02:03.67" />
                    <SPLIT distance="250" swimtime="00:02:36.08" />
                    <SPLIT distance="300" swimtime="00:03:08.75" />
                    <SPLIT distance="350" swimtime="00:03:41.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="616" swimtime="00:01:56.78" resultid="1585" heatid="2036" lane="4" entrytime="00:01:55.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.73" />
                    <SPLIT distance="100" swimtime="00:00:55.60" />
                    <SPLIT distance="150" swimtime="00:01:25.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17317" nation="BRA" region="PR" clubid="1502" name="Colégio Estadual Ernani Vidal, Curitiba" shortname="Ctba-Ernani Vidal,Ce">
          <ATHLETES>
            <ATHLETE firstname="Giovana" lastname="Reis" birthdate="2008-04-07" gender="F" nation="BRA" license="378820" swrid="5600243" athleteid="1503" externalid="378820" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1085" points="216" swimtime="00:01:23.68" resultid="1504" heatid="1989" lane="3" entrytime="00:01:22.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="240" swimtime="00:00:36.88" resultid="1505" heatid="2010" lane="7" entrytime="00:00:38.25" entrycourse="SCM" />
                <RESULT eventid="1183" points="167" swimtime="00:00:44.27" resultid="1506" heatid="2038" lane="1" entrytime="00:00:44.10" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18911" nation="BRA" region="PR" clubid="1729" name="Colégio Premier, Londrina" shortname="Ldna-Premier,C">
          <ATHLETES>
            <ATHLETE firstname="Guilherme" lastname="Kikuchi Fujii" birthdate="2007-01-04" gender="M" nation="BRA" license="297805" swrid="5603863" athleteid="1730" externalid="297805" level="G-OLIMPICA">
              <RESULTS>
                <RESULT eventid="1097" points="543" swimtime="00:00:30.57" resultid="1731" heatid="1996" lane="4" entrytime="00:00:30.35" entrycourse="SCM" />
                <RESULT eventid="1123" points="642" swimtime="00:02:19.23" resultid="1732" heatid="2007" lane="4" entrytime="00:02:24.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                    <SPLIT distance="100" swimtime="00:01:07.32" />
                    <SPLIT distance="150" swimtime="00:01:43.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="614" swimtime="00:01:05.02" resultid="1733" heatid="2045" lane="4" entrytime="00:01:05.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Betina" lastname="Tramontini Queiroz" birthdate="2007-09-11" gender="F" nation="BRA" license="357155" swrid="5658063" athleteid="1734" externalid="357155" level="VIBE">
              <RESULTS>
                <RESULT eventid="1085" status="WDR" swimtime="00:00:00.00" resultid="1735" entrytime="00:01:02.50" entrycourse="SCM" />
                <RESULT eventid="1111" status="WDR" swimtime="00:00:00.00" resultid="1736" entrytime="00:04:47.51" entrycourse="SCM" />
                <RESULT eventid="1175" status="WDR" swimtime="00:00:00.00" resultid="1737" entrytime="00:02:12.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4222" nation="BRA" region="PR" clubid="1682" name="Colégio Bertoni Internacional, Foz Do Iguaçu" shortname="Fozi-Bertoni Int.,C">
          <ATHLETES>
            <ATHLETE firstname="Lucas" lastname="Marques Petry" birthdate="2008-01-08" gender="M" nation="BRA" license="392351" swrid="4711489" athleteid="1683" externalid="392351" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1105" points="385" swimtime="00:19:23.33" resultid="1684" heatid="1999" lane="2" entrytime="00:19:05.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                    <SPLIT distance="100" swimtime="00:01:10.29" />
                    <SPLIT distance="150" swimtime="00:01:48.49" />
                    <SPLIT distance="200" swimtime="00:02:27.27" />
                    <SPLIT distance="250" swimtime="00:03:06.46" />
                    <SPLIT distance="300" swimtime="00:03:45.33" />
                    <SPLIT distance="350" swimtime="00:04:23.47" />
                    <SPLIT distance="400" swimtime="00:05:02.31" />
                    <SPLIT distance="450" swimtime="00:05:42.24" />
                    <SPLIT distance="500" swimtime="00:06:21.68" />
                    <SPLIT distance="550" swimtime="00:07:00.64" />
                    <SPLIT distance="600" swimtime="00:07:40.01" />
                    <SPLIT distance="650" swimtime="00:08:19.76" />
                    <SPLIT distance="700" swimtime="00:08:59.94" />
                    <SPLIT distance="750" swimtime="00:09:41.55" />
                    <SPLIT distance="800" swimtime="00:10:20.77" />
                    <SPLIT distance="850" swimtime="00:10:59.78" />
                    <SPLIT distance="900" swimtime="00:11:38.52" />
                    <SPLIT distance="950" swimtime="00:12:16.64" />
                    <SPLIT distance="1000" swimtime="00:12:54.60" />
                    <SPLIT distance="1050" swimtime="00:13:33.22" />
                    <SPLIT distance="1100" swimtime="00:14:11.12" />
                    <SPLIT distance="1150" swimtime="00:14:49.87" />
                    <SPLIT distance="1200" swimtime="00:15:29.27" />
                    <SPLIT distance="1250" swimtime="00:16:08.73" />
                    <SPLIT distance="1300" swimtime="00:16:48.73" />
                    <SPLIT distance="1350" swimtime="00:17:27.73" />
                    <SPLIT distance="1400" swimtime="00:18:06.39" />
                    <SPLIT distance="1450" swimtime="00:18:45.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="365" swimtime="00:04:56.75" resultid="1685" heatid="2004" lane="2" entrytime="00:04:42.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:07.62" />
                    <SPLIT distance="150" swimtime="00:01:45.59" />
                    <SPLIT distance="200" swimtime="00:02:25.19" />
                    <SPLIT distance="250" swimtime="00:03:03.29" />
                    <SPLIT distance="300" swimtime="00:03:41.80" />
                    <SPLIT distance="350" swimtime="00:04:20.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="356" swimtime="00:10:25.23" resultid="1686" heatid="2029" lane="3" entrytime="00:10:13.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="100" swimtime="00:01:13.58" />
                    <SPLIT distance="150" swimtime="00:01:53.16" />
                    <SPLIT distance="200" swimtime="00:02:33.29" />
                    <SPLIT distance="250" swimtime="00:03:13.20" />
                    <SPLIT distance="300" swimtime="00:03:53.41" />
                    <SPLIT distance="350" swimtime="00:04:33.26" />
                    <SPLIT distance="400" swimtime="00:05:13.09" />
                    <SPLIT distance="450" swimtime="00:05:53.30" />
                    <SPLIT distance="500" swimtime="00:06:32.36" />
                    <SPLIT distance="550" swimtime="00:07:11.47" />
                    <SPLIT distance="600" swimtime="00:07:51.47" />
                    <SPLIT distance="650" swimtime="00:08:30.99" />
                    <SPLIT distance="700" swimtime="00:09:11.03" />
                    <SPLIT distance="750" swimtime="00:09:48.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Marques Petry" birthdate="2008-01-08" gender="M" nation="BRA" license="392352" swrid="4795316" athleteid="1687" externalid="392352" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1081" points="383" swimtime="00:01:01.72" resultid="1688" heatid="1986" lane="1" entrytime="00:01:01.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="342" swimtime="00:05:03.48" resultid="1689" heatid="2004" lane="1" entrytime="00:05:03.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="100" swimtime="00:01:09.72" />
                    <SPLIT distance="150" swimtime="00:01:47.43" />
                    <SPLIT distance="200" swimtime="00:02:26.07" />
                    <SPLIT distance="250" swimtime="00:03:05.01" />
                    <SPLIT distance="300" swimtime="00:03:44.70" />
                    <SPLIT distance="350" swimtime="00:04:25.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="374" swimtime="00:02:17.86" resultid="1690" heatid="2036" lane="7" entrytime="00:02:16.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="100" swimtime="00:01:06.01" />
                    <SPLIT distance="150" swimtime="00:01:41.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Victoria Portela" birthdate="2009-12-04" gender="F" nation="BRA" license="383047" swrid="5596945" athleteid="1691" externalid="383047">
              <RESULTS>
                <RESULT eventid="1077" points="315" swimtime="00:00:37.10" resultid="1692" heatid="1982" lane="8" entrytime="00:00:37.77" entrycourse="SCM" />
                <RESULT eventid="1127" points="452" swimtime="00:00:29.87" resultid="1693" heatid="2011" lane="6" entrytime="00:00:29.33" entrycourse="SCM" />
                <RESULT eventid="1175" points="433" swimtime="00:02:25.75" resultid="1694" heatid="2034" lane="5" entrytime="00:02:29.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                    <SPLIT distance="100" swimtime="00:01:09.16" />
                    <SPLIT distance="150" swimtime="00:01:46.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18926" nation="BRA" region="PR" clubid="1913" name="Colégio Estadual Dario Vellozo, Londrina" shortname="Ldna-Dario Vello.,Ce">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Eduarda Larsen De Godoi Pinton" birthdate="2009-02-20" gender="F" nation="BRA" license="V414485" athleteid="1914" externalid="V414485">
              <RESULTS>
                <RESULT eventid="1199" status="DSQ" swimtime="00:00:00.00" resultid="1915" heatid="2047" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.38" />
                    <SPLIT distance="100" swimtime="00:01:53.15" />
                    <SPLIT distance="150" swimtime="00:02:54.47" />
                    <SPLIT distance="200" swimtime="00:03:58.13" />
                    <SPLIT distance="250" swimtime="00:05:03.24" />
                    <SPLIT distance="300" swimtime="00:06:08.46" />
                    <SPLIT distance="350" swimtime="00:07:14.18" />
                    <SPLIT distance="400" swimtime="00:08:20.41" />
                    <SPLIT distance="450" swimtime="00:09:26.99" />
                    <SPLIT distance="500" swimtime="00:10:34.46" />
                    <SPLIT distance="550" swimtime="00:11:42.86" />
                    <SPLIT distance="600" swimtime="00:12:51.06" />
                    <SPLIT distance="650" swimtime="00:14:00.33" />
                    <SPLIT distance="700" swimtime="00:15:10.44" />
                    <SPLIT distance="750" swimtime="00:16:21.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="135" swimtime="00:03:34.71" resultid="1916" heatid="2034" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.01" />
                    <SPLIT distance="100" swimtime="00:01:39.39" />
                    <SPLIT distance="150" swimtime="00:02:37.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18909" nation="BRA" region="PR" clubid="1229" name="Colégio Ecel Bandeirantes" shortname="Btes-Ecel,C">
          <ATHLETES>
            <ATHLETE firstname="Luis" lastname="Otavio Pedrozo De Lazzari" birthdate="2008-05-22" gender="M" nation="BRA" license="V414516" athleteid="1233" externalid="V414516">
              <RESULTS>
                <RESULT eventid="1081" points="194" swimtime="00:01:17.39" resultid="1234" heatid="1983" lane="3" />
                <RESULT eventid="1131" points="219" swimtime="00:00:33.41" resultid="1235" heatid="2012" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Guidi Amaro Costa" birthdate="2008-11-08" gender="M" nation="BRA" license="V414515" athleteid="1230" externalid="V414515">
              <RESULTS>
                <RESULT eventid="1081" points="254" swimtime="00:01:10.80" resultid="1231" heatid="1984" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="295" swimtime="00:00:30.27" resultid="1232" heatid="2014" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17332" nation="BRA" region="PR" clubid="1285" name="Colégio Estadual Ângelo Trevisan, Curitiba" shortname="Ctba-Ângelo Trev.,Ce">
          <ATHLETES>
            <ATHLETE firstname="Mayara" lastname="Fieber" birthdate="2008-08-20" gender="F" nation="BRA" license="391147" swrid="5600161" athleteid="1286" externalid="391147">
              <RESULTS>
                <RESULT eventid="1085" points="322" swimtime="00:01:13.26" resultid="1287" heatid="1989" lane="4" entrytime="00:01:13.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" status="DSQ" swimtime="00:00:00.00" resultid="1288" heatid="2024" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                    <SPLIT distance="100" swimtime="00:01:27.83" />
                    <SPLIT distance="150" swimtime="00:02:18.37" />
                    <SPLIT distance="200" swimtime="00:03:13.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="316" swimtime="00:00:35.77" resultid="1289" heatid="2037" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="8871" nation="BRA" region="PR" clubid="1530" name="Colégio Marista Santa Maria, Curitiba" shortname="Ctba-Marista St.Mª,C">
          <ATHLETES>
            <ATHLETE firstname="Laura" lastname="Da Costa Riekes" birthdate="2008-06-19" gender="F" nation="BRA" license="331686" swrid="5600143" athleteid="1531" externalid="331686" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1077" points="391" swimtime="00:00:34.53" resultid="1532" heatid="1980" lane="2" />
                <RESULT eventid="1127" points="453" swimtime="00:00:29.84" resultid="1533" heatid="2011" lane="2" entrytime="00:00:29.55" entrycourse="SCM" />
                <RESULT eventid="1183" points="449" swimtime="00:00:31.82" resultid="1534" heatid="2038" lane="5" entrytime="00:00:31.98" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17646" nation="BRA" region="PR" clubid="1620" name="Colégio Adventista De Cascavel" shortname="Cvel-Adventista,C">
          <ATHLETES>
            <ATHLETE firstname="Alice" lastname="Sehn Uren" birthdate="2009-10-15" gender="F" nation="BRA" license="357159" swrid="5596937" athleteid="1621" externalid="357159">
              <RESULTS>
                <RESULT eventid="1101" points="390" swimtime="00:00:38.81" resultid="1622" heatid="1997" lane="4" />
                <RESULT eventid="1135" points="374" swimtime="00:02:44.94" resultid="1623" heatid="2018" lane="6" entrytime="00:02:52.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                    <SPLIT distance="100" swimtime="00:01:20.56" />
                    <SPLIT distance="150" swimtime="00:02:03.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="374" swimtime="00:01:26.51" resultid="1624" heatid="2042" lane="6" entrytime="00:01:26.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13980" nation="BRA" region="PR" clubid="1695" name="CCM Presidente Costa E Silva, Foz Do Iguaçu" shortname="Fozi-Costa Silva,CCM">
          <ATHLETES>
            <ATHLETE firstname="Ana" lastname="Carolina Ghellere" birthdate="2007-06-05" gender="F" nation="BRA" license="312662" swrid="5596874" athleteid="1696" externalid="312662" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1093" points="540" swimtime="00:02:26.88" resultid="1697" heatid="1992" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                    <SPLIT distance="100" swimtime="00:01:09.63" />
                    <SPLIT distance="150" swimtime="00:01:47.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="502" swimtime="00:05:25.63" resultid="1698" heatid="2024" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:10.89" />
                    <SPLIT distance="150" swimtime="00:01:55.04" />
                    <SPLIT distance="200" swimtime="00:02:38.19" />
                    <SPLIT distance="250" swimtime="00:03:24.54" />
                    <SPLIT distance="300" swimtime="00:04:11.80" />
                    <SPLIT distance="350" swimtime="00:04:49.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="590" swimtime="00:02:11.48" resultid="1699" heatid="2034" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.19" />
                    <SPLIT distance="100" swimtime="00:01:03.70" />
                    <SPLIT distance="150" swimtime="00:01:37.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2633" nation="BRA" region="PR" clubid="1640" name="Colégio Ideal, Cascavel" shortname="Cvel-Ideal,C">
          <ATHLETES>
            <ATHLETE firstname="Henrique" lastname="Tolentino Smarczewski" birthdate="2008-09-01" gender="M" nation="BRA" license="378818" swrid="5596941" athleteid="1641" externalid="378818">
              <RESULTS>
                <RESULT eventid="1105" points="454" swimtime="00:18:21.67" resultid="1642" heatid="1999" lane="3" entrytime="00:18:32.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                    <SPLIT distance="100" swimtime="00:01:06.94" />
                    <SPLIT distance="150" swimtime="00:01:42.51" />
                    <SPLIT distance="200" swimtime="00:02:18.70" />
                    <SPLIT distance="250" swimtime="00:02:55.03" />
                    <SPLIT distance="350" swimtime="00:04:07.22" />
                    <SPLIT distance="400" swimtime="00:04:44.43" />
                    <SPLIT distance="450" swimtime="00:05:20.93" />
                    <SPLIT distance="500" swimtime="00:05:58.14" />
                    <SPLIT distance="550" swimtime="00:06:35.58" />
                    <SPLIT distance="600" swimtime="00:07:12.71" />
                    <SPLIT distance="650" swimtime="00:07:49.89" />
                    <SPLIT distance="700" swimtime="00:08:26.77" />
                    <SPLIT distance="750" swimtime="00:09:04.70" />
                    <SPLIT distance="800" swimtime="00:09:41.97" />
                    <SPLIT distance="850" swimtime="00:10:19.35" />
                    <SPLIT distance="900" swimtime="00:10:56.80" />
                    <SPLIT distance="950" swimtime="00:11:34.53" />
                    <SPLIT distance="1000" swimtime="00:12:12.24" />
                    <SPLIT distance="1050" swimtime="00:12:49.23" />
                    <SPLIT distance="1100" swimtime="00:13:27.13" />
                    <SPLIT distance="1150" swimtime="00:14:04.44" />
                    <SPLIT distance="1200" swimtime="00:14:43.19" />
                    <SPLIT distance="1250" swimtime="00:15:19.03" />
                    <SPLIT distance="1300" swimtime="00:15:56.49" />
                    <SPLIT distance="1350" swimtime="00:16:33.84" />
                    <SPLIT distance="1400" swimtime="00:17:11.54" />
                    <SPLIT distance="1450" swimtime="00:17:47.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" status="DSQ" swimtime="00:02:50.56" resultid="1643" heatid="2007" lane="8" entrytime="00:02:41.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:01:20.98" />
                    <SPLIT distance="150" swimtime="00:02:05.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="446" swimtime="00:02:10.05" resultid="1644" heatid="2036" lane="6" entrytime="00:02:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="100" swimtime="00:01:02.03" />
                    <SPLIT distance="150" swimtime="00:01:35.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15598" nation="BRA" region="PR" clubid="1748" name="Colégio De Aplicação Pedagógica Uem, Maringá" shortname="Mrga-Aplicação Uem,C">
          <ATHLETES>
            <ATHLETE firstname="Gabriel" lastname="Casavechia Carraro" birthdate="2009-07-28" gender="M" nation="BRA" license="368150" swrid="5384752" athleteid="1749" externalid="368150">
              <RESULTS>
                <RESULT eventid="1081" points="566" swimtime="00:00:54.20" resultid="1750" heatid="1987" lane="3" entrytime="00:00:54.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="519" swimtime="00:00:59.42" resultid="1751" heatid="2023" lane="4" entrytime="00:01:00.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="561" swimtime="00:02:00.43" resultid="1752" heatid="2036" lane="5" entrytime="00:01:58.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.29" />
                    <SPLIT distance="100" swimtime="00:00:57.02" />
                    <SPLIT distance="150" swimtime="00:01:27.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2603" nation="BRA" region="PR" clubid="1851" name="Colégio Sagrada Família, Ponta Grossa" shortname="Pgro-Sagrada Fami.,C">
          <ATHLETES>
            <ATHLETE firstname="Victor" lastname="Carraro Borges" birthdate="2009-05-11" gender="M" nation="BRA" license="345590" swrid="5622267" athleteid="1852" externalid="345590" level="SAGRADA FA">
              <RESULTS>
                <RESULT eventid="1105" points="402" swimtime="00:19:07.28" resultid="1853" heatid="1999" lane="6" entrytime="00:18:48.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:09.96" />
                    <SPLIT distance="150" swimtime="00:01:47.30" />
                    <SPLIT distance="200" swimtime="00:02:25.00" />
                    <SPLIT distance="250" swimtime="00:03:02.54" />
                    <SPLIT distance="300" swimtime="00:03:41.59" />
                    <SPLIT distance="350" swimtime="00:04:20.09" />
                    <SPLIT distance="400" swimtime="00:04:59.13" />
                    <SPLIT distance="450" swimtime="00:05:38.41" />
                    <SPLIT distance="500" swimtime="00:06:18.19" />
                    <SPLIT distance="550" swimtime="00:06:56.83" />
                    <SPLIT distance="600" swimtime="00:07:36.07" />
                    <SPLIT distance="650" swimtime="00:08:15.19" />
                    <SPLIT distance="700" swimtime="00:08:54.14" />
                    <SPLIT distance="750" swimtime="00:09:33.32" />
                    <SPLIT distance="800" swimtime="00:10:12.74" />
                    <SPLIT distance="850" swimtime="00:10:51.54" />
                    <SPLIT distance="900" swimtime="00:11:30.16" />
                    <SPLIT distance="950" swimtime="00:12:09.63" />
                    <SPLIT distance="1000" swimtime="00:12:48.20" />
                    <SPLIT distance="1050" swimtime="00:13:26.47" />
                    <SPLIT distance="1100" swimtime="00:14:04.70" />
                    <SPLIT distance="1150" swimtime="00:14:41.92" />
                    <SPLIT distance="1200" swimtime="00:15:19.71" />
                    <SPLIT distance="1250" swimtime="00:15:57.90" />
                    <SPLIT distance="1300" swimtime="00:16:35.88" />
                    <SPLIT distance="1350" swimtime="00:17:13.86" />
                    <SPLIT distance="1400" swimtime="00:17:52.21" />
                    <SPLIT distance="1450" swimtime="00:18:25.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="416" swimtime="00:04:44.21" resultid="1854" heatid="2004" lane="7" entrytime="00:04:45.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:40.96" />
                    <SPLIT distance="200" swimtime="00:02:17.79" />
                    <SPLIT distance="250" swimtime="00:02:54.46" />
                    <SPLIT distance="300" swimtime="00:03:31.57" />
                    <SPLIT distance="350" swimtime="00:04:08.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="393" swimtime="00:10:05.32" resultid="1855" heatid="2029" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                    <SPLIT distance="100" swimtime="00:01:11.38" />
                    <SPLIT distance="150" swimtime="00:01:49.47" />
                    <SPLIT distance="200" swimtime="00:02:26.98" />
                    <SPLIT distance="250" swimtime="00:03:05.88" />
                    <SPLIT distance="300" swimtime="00:03:44.09" />
                    <SPLIT distance="350" swimtime="00:04:23.32" />
                    <SPLIT distance="400" swimtime="00:05:01.90" />
                    <SPLIT distance="450" swimtime="00:05:41.31" />
                    <SPLIT distance="500" swimtime="00:06:20.35" />
                    <SPLIT distance="550" swimtime="00:06:58.39" />
                    <SPLIT distance="600" swimtime="00:07:37.11" />
                    <SPLIT distance="650" swimtime="00:08:14.86" />
                    <SPLIT distance="700" swimtime="00:08:52.41" />
                    <SPLIT distance="750" swimtime="00:09:29.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13349" nation="BRA" region="PR" clubid="1300" name="Colégio Bom Jesus Centro, Curitiba" shortname="Ctba-Bj Centro,C">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Carolina Biella Misocami" birthdate="2009-02-19" gender="F" nation="BRA" license="V339455" athleteid="1313" externalid="V339455">
              <RESULTS>
                <RESULT eventid="1085" points="188" swimtime="00:01:27.59" resultid="1314" heatid="1989" lane="6" entrytime="00:01:33.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="182" swimtime="00:00:49.99" resultid="1315" heatid="1998" lane="7" entrytime="00:00:56.42" entrycourse="SCM" />
                <RESULT eventid="1127" points="191" swimtime="00:00:39.80" resultid="1316" heatid="2009" lane="4" entrytime="00:00:41.69" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Garcia De Fraga" birthdate="2009-03-24" gender="M" nation="BRA" license="342147" swrid="5600172" athleteid="1301" externalid="342147" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1065" points="537" swimtime="00:02:14.86" resultid="1302" heatid="1976" lane="4" entrytime="00:02:11.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.54" />
                    <SPLIT distance="100" swimtime="00:01:01.72" />
                    <SPLIT distance="150" swimtime="00:01:41.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="521" swimtime="00:02:11.19" resultid="1303" heatid="2019" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.54" />
                    <SPLIT distance="100" swimtime="00:01:02.68" />
                    <SPLIT distance="150" swimtime="00:01:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="534" swimtime="00:00:59.57" resultid="1304" heatid="2033" lane="4" entrytime="00:00:59.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Zanini Duarte" birthdate="2009-03-27" gender="M" nation="BRA" license="V383394" athleteid="1317" externalid="V383394">
              <RESULTS>
                <RESULT eventid="1097" points="232" swimtime="00:00:40.58" resultid="1318" heatid="1995" lane="6" entrytime="00:00:43.91" entrycourse="SCM" />
                <RESULT eventid="1131" points="251" swimtime="00:00:31.93" resultid="1319" heatid="2012" lane="3" />
                <RESULT eventid="1163" status="DSQ" swimtime="00:00:00.00" resultid="1320" heatid="2028" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                    <SPLIT distance="100" swimtime="00:01:17.99" />
                    <SPLIT distance="150" swimtime="00:02:03.59" />
                    <SPLIT distance="200" swimtime="00:02:51.53" />
                    <SPLIT distance="250" swimtime="00:03:40.51" />
                    <SPLIT distance="300" swimtime="00:04:29.98" />
                    <SPLIT distance="350" swimtime="00:05:20.54" />
                    <SPLIT distance="400" swimtime="00:06:11.88" />
                    <SPLIT distance="450" swimtime="00:07:03.67" />
                    <SPLIT distance="500" swimtime="00:07:59.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo" lastname="De Lima Cavalcanti" birthdate="2009-12-17" gender="M" nation="BRA" license="380965" swrid="5634589" athleteid="1305" externalid="380965">
              <RESULTS>
                <RESULT eventid="1089" points="382" swimtime="00:02:27.17" resultid="1306" heatid="1991" lane="3" entrytime="00:02:22.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:10.91" />
                    <SPLIT distance="150" swimtime="00:01:49.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="426" swimtime="00:01:03.48" resultid="1307" heatid="2023" lane="6" entrytime="00:01:01.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="438" swimtime="00:00:26.54" resultid="1308" heatid="2017" lane="1" entrytime="00:00:25.95" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Neves Vianna" birthdate="2007-12-30" gender="F" nation="BRA" license="391106" swrid="5600223" athleteid="1309" externalid="391106">
              <RESULTS>
                <RESULT eventid="1085" points="271" swimtime="00:01:17.61" resultid="1310" heatid="1989" lane="5" entrytime="00:01:22.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="223" swimtime="00:01:30.49" resultid="1311" heatid="2030" lane="5" entrytime="00:01:31.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="226" swimtime="00:03:00.97" resultid="1312" heatid="2034" lane="6" entrytime="00:03:00.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                    <SPLIT distance="100" swimtime="00:01:26.01" />
                    <SPLIT distance="150" swimtime="00:02:13.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2653" nation="BRA" region="PR" clubid="1605" name="Escola Seb Dom Bosco Batel, Curitiba" shortname="Ctba-Seb Batel,E">
          <ATHLETES>
            <ATHLETE firstname="Rafaela" lastname="Yolanda Ferreira" birthdate="2008-03-17" gender="F" nation="BRA" license="358335" swrid="5600276" athleteid="1606" externalid="358335">
              <RESULTS>
                <RESULT eventid="1101" points="414" swimtime="00:00:38.06" resultid="1607" heatid="1998" lane="5" entrytime="00:00:36.77" entrycourse="SCM" />
                <RESULT eventid="1119" points="447" swimtime="00:02:55.87" resultid="1608" heatid="2005" lane="5" entrytime="00:02:52.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                    <SPLIT distance="100" swimtime="00:01:23.68" />
                    <SPLIT distance="150" swimtime="00:02:09.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="436" swimtime="00:01:22.19" resultid="1609" heatid="2042" lane="5" entrytime="00:01:19.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17330" nation="BRA" region="PR" clubid="1245" name="Instituto Federal Do Paraná, Colombo" shortname="Clbo-Ifpr">
          <ATHLETES>
            <ATHLETE firstname="Arthur" lastname="Arceli Silva" birthdate="2008-03-04" gender="M" nation="BRA" license="331565" swrid="5385686" athleteid="1246" externalid="331565" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1081" points="322" swimtime="00:01:05.37" resultid="1247" heatid="1984" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="292" swimtime="00:01:11.98" resultid="1248" heatid="2022" lane="4" entrytime="00:01:08.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="316" swimtime="00:01:10.90" resultid="1249" heatid="2033" lane="1" entrytime="00:01:09.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="9861" nation="BRA" region="PR" clubid="1558" name="Colégio Positivo Ângelo Sampaio, Curitiba" shortname="Ctba-Posi. Ângelo,C">
          <ATHLETES>
            <ATHLETE firstname="Fabiana" lastname="Zaleski Dallazem" birthdate="2009-05-16" gender="F" nation="BRA" license="344287" swrid="5600279" athleteid="1559" externalid="344287" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1077" points="501" swimtime="00:00:31.79" resultid="1560" heatid="1982" lane="5" entrytime="00:00:32.02" entrycourse="SCM" />
                <RESULT eventid="1135" points="461" swimtime="00:02:33.90" resultid="1561" heatid="2018" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                    <SPLIT distance="100" swimtime="00:01:14.31" />
                    <SPLIT distance="150" swimtime="00:01:54.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="488" swimtime="00:01:09.68" resultid="1562" heatid="2031" lane="5" entrytime="00:01:09.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Araujo Do Rego Barros" birthdate="2009-04-30" gender="M" nation="BRA" license="376325" swrid="5377739" athleteid="1575" externalid="376325">
              <RESULTS>
                <RESULT eventid="1081" points="344" swimtime="00:01:03.97" resultid="1576" heatid="1985" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1089" status="DSQ" swimtime="00:03:36.00" resultid="1577" heatid="1991" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="279" swimtime="00:01:13.09" resultid="1578" heatid="2022" lane="3" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Araujo Barros" birthdate="2008-12-26" gender="M" nation="BRA" license="331713" swrid="5367497" athleteid="1563" externalid="331713">
              <RESULTS>
                <RESULT eventid="1115" points="572" swimtime="00:04:15.66" resultid="1564" heatid="2004" lane="5" entrytime="00:04:11.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.07" />
                    <SPLIT distance="100" swimtime="00:00:59.51" />
                    <SPLIT distance="150" swimtime="00:01:31.26" />
                    <SPLIT distance="200" swimtime="00:02:03.39" />
                    <SPLIT distance="250" swimtime="00:02:36.30" />
                    <SPLIT distance="300" swimtime="00:03:09.68" />
                    <SPLIT distance="350" swimtime="00:03:43.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="542" swimtime="00:02:01.83" resultid="1565" heatid="2035" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.27" />
                    <SPLIT distance="100" swimtime="00:00:57.90" />
                    <SPLIT distance="150" swimtime="00:01:30.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="566" swimtime="00:08:56.02" resultid="1566" heatid="2028" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                    <SPLIT distance="100" swimtime="00:01:02.49" />
                    <SPLIT distance="150" swimtime="00:01:35.40" />
                    <SPLIT distance="200" swimtime="00:02:08.80" />
                    <SPLIT distance="250" swimtime="00:02:41.81" />
                    <SPLIT distance="300" swimtime="00:03:15.24" />
                    <SPLIT distance="350" swimtime="00:03:48.99" />
                    <SPLIT distance="400" swimtime="00:04:22.84" />
                    <SPLIT distance="450" swimtime="00:04:56.97" />
                    <SPLIT distance="500" swimtime="00:05:30.89" />
                    <SPLIT distance="550" swimtime="00:06:05.37" />
                    <SPLIT distance="600" swimtime="00:06:39.58" />
                    <SPLIT distance="650" swimtime="00:07:14.00" />
                    <SPLIT distance="700" swimtime="00:07:48.40" />
                    <SPLIT distance="750" swimtime="00:08:22.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Guimaraes E Souza" birthdate="2008-12-21" gender="M" nation="BRA" license="376972" swrid="5600182" athleteid="1567" externalid="376972">
              <RESULTS>
                <RESULT eventid="1065" status="WDR" swimtime="00:00:00.00" resultid="1568" entrytime="00:02:31.56" entrycourse="SCM" />
                <RESULT eventid="1123" status="WDR" swimtime="00:00:00.00" resultid="1569" />
                <RESULT eventid="1195" status="WDR" swimtime="00:00:00.00" resultid="1570" entrytime="00:01:12.63" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Zaleski Dallazem" birthdate="2009-05-16" gender="M" nation="BRA" license="344286" swrid="5600280" athleteid="1571" externalid="344286" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1081" points="405" swimtime="00:01:00.60" resultid="1572" heatid="1986" lane="7" entrytime="00:01:00.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" status="DSQ" swimtime="00:01:07.66" resultid="1573" heatid="2022" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="392" swimtime="00:01:15.53" resultid="1574" heatid="2045" lane="8" entrytime="00:01:15.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="COL POSI ANG SAMPAIO &apos;&apos;A&apos;&apos;" number="1">
              <RESULTS>
                <RESULT eventid="1161" status="WDR" swimtime="00:00:00.00" resultid="1579" heatid="2027" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="2" reactiontime="0" />
                    <RELAYPOSITION number="3" reactiontime="0" />
                    <RELAYPOSITION number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1203" status="WDR" swimtime="00:00:00.00" resultid="1580" heatid="2048" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="2" reactiontime="0" />
                    <RELAYPOSITION number="3" reactiontime="0" />
                    <RELAYPOSITION number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="11380" nation="BRA" region="PR" clubid="1625" name="Colégio Nossa Srª. Auxiliadora, Cascavel" shortname="Cvel-Auxiliadora,C">
          <ATHLETES>
            <ATHLETE firstname="Gabriel" lastname="Alves Serafini" birthdate="2008-04-15" gender="M" nation="BRA" license="351644" swrid="5596867" athleteid="1626" externalid="351644">
              <RESULTS>
                <RESULT eventid="1089" points="434" swimtime="00:02:21.05" resultid="1627" heatid="1991" lane="6" entrytime="00:02:23.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.52" />
                    <SPLIT distance="100" swimtime="00:01:04.49" />
                    <SPLIT distance="150" swimtime="00:01:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="392" swimtime="00:01:05.26" resultid="1628" heatid="2023" lane="3" entrytime="00:01:01.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1179" points="450" swimtime="00:02:09.61" resultid="1629" heatid="2036" lane="3" entrytime="00:02:07.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.91" />
                    <SPLIT distance="100" swimtime="00:01:01.15" />
                    <SPLIT distance="150" swimtime="00:01:35.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15584" nation="BRA" region="PR" clubid="1753" name="Colégio Axia, Maringá" shortname="Mrga-Axia,C">
          <ATHLETES>
            <ATHLETE firstname="Wellington" lastname="De Lima" birthdate="2008-03-01" gender="M" nation="BRA" license="370024" swrid="5470912" athleteid="1754" externalid="370024">
              <RESULTS>
                <RESULT eventid="1081" points="472" swimtime="00:00:57.57" resultid="1755" heatid="1987" lane="1" entrytime="00:00:56.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="466" swimtime="00:00:25.99" resultid="1756" heatid="2016" lane="4" entrytime="00:00:26.13" entrycourse="SCM" />
                <RESULT eventid="1179" status="DSQ" swimtime="00:02:08.28" resultid="1757" heatid="2036" lane="2" entrytime="00:02:10.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.34" />
                    <SPLIT distance="100" swimtime="00:01:00.39" />
                    <SPLIT distance="150" swimtime="00:01:34.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Antonio Mendes" birthdate="2008-12-04" gender="M" nation="BRA" license="366962" swrid="5196287" athleteid="1758" externalid="366962">
              <RESULTS>
                <RESULT eventid="1097" points="501" swimtime="00:00:31.40" resultid="1759" heatid="1996" lane="6" entrytime="00:00:31.69" entrycourse="SCM" />
                <RESULT eventid="1123" points="527" swimtime="00:02:28.73" resultid="1760" heatid="2007" lane="3" entrytime="00:02:34.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                    <SPLIT distance="100" swimtime="00:01:10.36" />
                    <SPLIT distance="150" swimtime="00:01:48.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="536" swimtime="00:01:08.02" resultid="1761" heatid="2045" lane="3" entrytime="00:01:08.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="739" nation="BRA" region="PR" clubid="1265" name="CCM Marechal Rondon, Campo Mourão" shortname="Cmou-Mar. Rondon,CCM">
          <ATHLETES>
            <ATHLETE firstname="Pedro" lastname="Henrique De Oliveira" birthdate="2009-07-28" gender="M" nation="BRA" license="V414505" athleteid="1266" externalid="V414505">
              <RESULTS>
                <RESULT eventid="1081" points="296" swimtime="00:01:07.28" resultid="1267" heatid="1983" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="327" swimtime="00:00:29.25" resultid="1268" heatid="2013" lane="4" />
                <RESULT eventid="1187" points="296" swimtime="00:00:32.62" resultid="1269" heatid="2040" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6582" nation="BRA" region="PR" clubid="1290" name="Colégio Padre João Bagozzi, Curitiba" shortname="Ctba-Bagozzi,C">
          <ATHLETES>
            <ATHLETE firstname="Bianca" lastname="Liz Skowronski" birthdate="2008-01-24" gender="F" nation="BRA" license="358245" swrid="5600202" athleteid="1291" externalid="358245">
              <RESULTS>
                <RESULT eventid="1077" points="324" swimtime="00:00:36.76" resultid="1292" heatid="1982" lane="1" entrytime="00:00:37.30" entrycourse="SCM" />
                <RESULT eventid="1135" points="359" swimtime="00:02:47.35" resultid="1293" heatid="2018" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.22" />
                    <SPLIT distance="100" swimtime="00:01:21.08" />
                    <SPLIT distance="150" swimtime="00:02:03.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="328" swimtime="00:01:19.54" resultid="1294" heatid="2031" lane="1" entrytime="00:01:17.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18905" nation="BRA" region="PR" clubid="1275" name="3º Colégio Da Polícia Militar, Cornélio Procópio" shortname="Cpro-3ºcpm,C">
          <ATHLETES>
            <ATHLETE firstname="Gustavo" lastname="Taborda Medeiros" birthdate="2007-09-21" gender="M" nation="BRA" license="V414517" athleteid="1276" externalid="V414517">
              <RESULTS>
                <RESULT eventid="1081" points="222" swimtime="00:01:13.95" resultid="1277" heatid="1984" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="289" swimtime="00:00:30.47" resultid="1278" heatid="2013" lane="8" />
                <RESULT eventid="1187" points="159" swimtime="00:00:40.11" resultid="1279" heatid="2040" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13350" nation="BRA" region="PR" clubid="1321" name="Colégio Bom Jesus Nossa Srª. De Lourdes, Curitiba" shortname="Ctba-Bj Lourdes,C">
          <ATHLETES>
            <ATHLETE firstname="Enzo" lastname="Inoue Kuroda" birthdate="2009-04-18" gender="M" nation="BRA" license="324700" swrid="5600190" athleteid="1334" externalid="324700">
              <RESULTS>
                <RESULT eventid="1105" points="463" swimtime="00:18:14.22" resultid="1335" heatid="1999" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="100" swimtime="00:01:07.40" />
                    <SPLIT distance="150" swimtime="00:01:44.00" />
                    <SPLIT distance="200" swimtime="00:02:20.47" />
                    <SPLIT distance="250" swimtime="00:02:57.35" />
                    <SPLIT distance="300" swimtime="00:03:34.91" />
                    <SPLIT distance="350" swimtime="00:04:12.07" />
                    <SPLIT distance="400" swimtime="00:04:49.55" />
                    <SPLIT distance="450" swimtime="00:05:26.70" />
                    <SPLIT distance="500" swimtime="00:06:03.45" />
                    <SPLIT distance="550" swimtime="00:06:41.17" />
                    <SPLIT distance="600" swimtime="00:07:18.20" />
                    <SPLIT distance="650" swimtime="00:07:56.60" />
                    <SPLIT distance="700" swimtime="00:08:32.86" />
                    <SPLIT distance="750" swimtime="00:09:10.33" />
                    <SPLIT distance="800" swimtime="00:09:47.05" />
                    <SPLIT distance="850" swimtime="00:10:23.57" />
                    <SPLIT distance="900" swimtime="00:10:59.98" />
                    <SPLIT distance="950" swimtime="00:11:36.61" />
                    <SPLIT distance="1000" swimtime="00:12:13.74" />
                    <SPLIT distance="1050" swimtime="00:12:50.93" />
                    <SPLIT distance="1100" swimtime="00:13:27.54" />
                    <SPLIT distance="1150" swimtime="00:14:04.04" />
                    <SPLIT distance="1200" swimtime="00:14:41.42" />
                    <SPLIT distance="1250" swimtime="00:15:17.49" />
                    <SPLIT distance="1300" swimtime="00:15:54.02" />
                    <SPLIT distance="1350" swimtime="00:16:30.88" />
                    <SPLIT distance="1400" swimtime="00:17:07.80" />
                    <SPLIT distance="1450" swimtime="00:17:49.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="419" swimtime="00:00:26.94" resultid="1336" heatid="2016" lane="3" entrytime="00:00:26.61" entrycourse="SCM" />
                <RESULT eventid="1163" points="543" swimtime="00:09:03.45" resultid="1337" heatid="2029" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.44" />
                    <SPLIT distance="150" swimtime="00:01:36.38" />
                    <SPLIT distance="200" swimtime="00:02:10.61" />
                    <SPLIT distance="250" swimtime="00:02:44.58" />
                    <SPLIT distance="300" swimtime="00:03:18.84" />
                    <SPLIT distance="350" swimtime="00:03:52.74" />
                    <SPLIT distance="400" swimtime="00:04:27.14" />
                    <SPLIT distance="450" swimtime="00:05:01.75" />
                    <SPLIT distance="500" swimtime="00:05:36.42" />
                    <SPLIT distance="550" swimtime="00:06:10.91" />
                    <SPLIT distance="600" swimtime="00:06:46.04" />
                    <SPLIT distance="650" swimtime="00:07:20.67" />
                    <SPLIT distance="700" swimtime="00:07:55.30" />
                    <SPLIT distance="750" swimtime="00:08:29.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thiago" lastname="Kozera Chiarato" birthdate="2008-01-22" gender="M" nation="BRA" license="406728" swrid="5717276" athleteid="1354" externalid="406728">
              <RESULTS>
                <RESULT eventid="1081" points="393" swimtime="00:01:01.21" resultid="1355" heatid="1985" lane="2" entrytime="00:01:06.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="339" swimtime="00:00:28.90" resultid="1356" heatid="2015" lane="6" entrytime="00:00:29.27" entrycourse="SCM" />
                <RESULT eventid="1187" status="DSQ" swimtime="00:00:30.90" resultid="1357" heatid="2040" lane="5" entrytime="00:00:32.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Oenning Ihlenffeldt" birthdate="2009-05-29" gender="F" nation="BRA" license="V414478" athleteid="1370" externalid="V414478">
              <RESULTS>
                <RESULT eventid="1085" points="221" swimtime="00:01:23.03" resultid="1371" heatid="1988" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="200" swimtime="00:00:43.14" resultid="1372" heatid="1980" lane="6" />
                <RESULT eventid="1101" points="191" swimtime="00:00:49.26" resultid="1373" heatid="1997" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="De Curcio" birthdate="2009-07-24" gender="F" nation="BRA" license="V383045" athleteid="1358" externalid="V383045">
              <RESULTS>
                <RESULT eventid="1077" status="WDR" swimtime="00:00:00.00" resultid="1359" />
                <RESULT eventid="1101" status="WDR" swimtime="00:00:00.00" resultid="1360" entrytime="00:00:50.58" entrycourse="SCM" />
                <RESULT eventid="1191" status="WDR" swimtime="00:00:00.00" resultid="1361" entrytime="00:01:59.11" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="F" nation="BRA" license="344301" swrid="5569976" athleteid="1322" externalid="344301">
              <RESULTS>
                <RESULT eventid="1093" points="483" swimtime="00:02:32.39" resultid="1323" heatid="1992" lane="4" entrytime="00:02:30.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:11.73" />
                    <SPLIT distance="150" swimtime="00:01:51.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="494" swimtime="00:01:08.37" resultid="1324" heatid="2020" lane="4" entrytime="00:01:06.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1183" points="476" swimtime="00:00:31.21" resultid="1325" heatid="2038" lane="4" entrytime="00:00:30.68" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Ieger" birthdate="2009-02-20" gender="M" nation="BRA" license="356888" swrid="5600180" athleteid="1338" externalid="356888">
              <RESULTS>
                <RESULT eventid="1097" points="352" swimtime="00:00:35.32" resultid="1339" heatid="1994" lane="6" />
                <RESULT eventid="1131" points="385" swimtime="00:00:27.71" resultid="1340" heatid="2016" lane="6" entrytime="00:00:26.62" entrycourse="SCM" />
                <RESULT eventid="1195" points="325" swimtime="00:01:20.34" resultid="1341" heatid="2045" lane="1" entrytime="00:01:15.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathalia" lastname="Lourenco Osorio" birthdate="2007-04-14" gender="F" nation="BRA" license="307465" swrid="5600203" athleteid="1326" externalid="307465">
              <RESULTS>
                <RESULT eventid="1077" status="WDR" swimtime="00:00:00.00" resultid="1327" entrytime="00:00:31.77" entrycourse="SCM" />
                <RESULT eventid="1127" status="WDR" swimtime="00:00:00.00" resultid="1328" entrytime="00:00:28.10" entrycourse="SCM" />
                <RESULT eventid="1167" status="WDR" swimtime="00:00:00.00" resultid="1329" entrytime="00:01:08.06" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anita" lastname="Gomes Saldanha" birthdate="2009-02-26" gender="F" nation="BRA" license="V399518" athleteid="1346" externalid="V399518">
              <RESULTS>
                <RESULT eventid="1085" points="194" swimtime="00:01:26.73" resultid="1347" heatid="1989" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="244" swimtime="00:00:36.66" resultid="1348" heatid="2010" lane="8" entrytime="00:00:38.77" entrycourse="SCM" />
                <RESULT eventid="1183" points="218" swimtime="00:00:40.48" resultid="1349" heatid="2038" lane="7" entrytime="00:00:43.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Zanardi" birthdate="2008-10-02" gender="F" nation="BRA" license="V398572" athleteid="1342" externalid="V398572">
              <RESULTS>
                <RESULT eventid="1069" points="241" swimtime="00:03:15.78" resultid="1343" heatid="1977" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.97" />
                    <SPLIT distance="100" swimtime="00:01:33.01" />
                    <SPLIT distance="150" swimtime="00:02:29.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="225" swimtime="00:00:46.61" resultid="1344" heatid="1998" lane="1" />
                <RESULT eventid="1127" points="284" swimtime="00:00:34.86" resultid="1345" heatid="2009" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Pacheco E Silva" birthdate="2008-04-28" gender="M" nation="BRA" license="V383390" athleteid="1362" externalid="V383390">
              <RESULTS>
                <RESULT eventid="1081" points="214" swimtime="00:01:14.96" resultid="1363" heatid="1984" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" status="DNS" swimtime="00:00:00.00" resultid="1364" heatid="1994" lane="2" />
                <RESULT eventid="1195" points="215" swimtime="00:01:32.24" resultid="1365" heatid="2043" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Bastos Costa" birthdate="2009-09-26" gender="F" nation="BRA" license="V399683" athleteid="1350" externalid="V399683">
              <RESULTS>
                <RESULT eventid="1085" points="260" swimtime="00:01:18.71" resultid="1351" heatid="1989" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="225" swimtime="00:00:41.48" resultid="1352" heatid="1981" lane="3" entrytime="00:00:45.16" entrycourse="SCM" />
                <RESULT eventid="1127" points="330" swimtime="00:00:33.18" resultid="1353" heatid="2010" lane="2" entrytime="00:00:35.46" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Henrique Ercoli" birthdate="2009-02-12" gender="M" nation="BRA" license="V383392" athleteid="1366" externalid="V383392">
              <RESULTS>
                <RESULT eventid="1081" points="223" swimtime="00:01:13.85" resultid="1367" heatid="1985" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1115" points="222" swimtime="00:05:50.46" resultid="1368" heatid="2003" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.27" />
                    <SPLIT distance="100" swimtime="00:01:18.14" />
                    <SPLIT distance="150" swimtime="00:02:01.74" />
                    <SPLIT distance="200" swimtime="00:02:46.16" />
                    <SPLIT distance="250" swimtime="00:03:31.53" />
                    <SPLIT distance="300" swimtime="00:04:18.00" />
                    <SPLIT distance="350" swimtime="00:05:04.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" status="DSQ" swimtime="00:00:00.00" resultid="1369" heatid="2029" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabrizio" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="M" nation="BRA" license="344303" swrid="5559846" athleteid="1330" externalid="344303">
              <RESULTS>
                <RESULT eventid="1089" status="DSQ" swimtime="00:02:32.69" resultid="1331" heatid="1991" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.47" />
                    <SPLIT distance="100" swimtime="00:01:10.04" />
                    <SPLIT distance="150" swimtime="00:01:50.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="389" swimtime="00:01:05.41" resultid="1332" heatid="2023" lane="7" entrytime="00:01:03.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="454" swimtime="00:00:28.28" resultid="1333" heatid="2041" lane="7" entrytime="00:00:28.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CTBA-BJ LOURDES,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1161" points="423" swimtime="00:01:48.91" resultid="1376" heatid="2027" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.54" />
                    <SPLIT distance="100" swimtime="00:00:55.46" />
                    <SPLIT distance="150" swimtime="00:01:22.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1338" number="1" />
                    <RELAYPOSITION athleteid="1354" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1330" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1334" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1203" points="398" swimtime="00:02:01.94" resultid="1377" heatid="2048" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                    <SPLIT distance="100" swimtime="00:01:06.01" />
                    <SPLIT distance="150" swimtime="00:01:34.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1334" number="1" />
                    <RELAYPOSITION athleteid="1338" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1330" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1354" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="CTBA-BJ LOURDES,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1159" points="340" swimtime="00:02:12.52" resultid="1374" heatid="2026" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.49" />
                    <SPLIT distance="150" swimtime="00:01:39.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1322" number="1" />
                    <RELAYPOSITION athleteid="1346" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1342" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1350" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1205" points="277" swimtime="00:02:36.96" resultid="1375" heatid="2049" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                    <SPLIT distance="100" swimtime="00:01:28.83" />
                    <SPLIT distance="150" swimtime="00:02:00.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1350" number="1" />
                    <RELAYPOSITION athleteid="1342" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1322" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1346" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="CTBA-BJ LOURDES,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1109" points="360" swimtime="00:02:13.65" resultid="1378" heatid="2000" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:07.70" />
                    <SPLIT distance="150" swimtime="00:01:38.74" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1334" number="1" />
                    <RELAYPOSITION athleteid="1338" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1322" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1342" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="17679" nation="BRA" region="PR" clubid="1487" name="Colégio Estadual D. Branca Do Nasci. Miranda, Ctba" shortname="Ctba-Dona Branca,Ce">
          <ATHLETES>
            <ATHLETE firstname="Stella" lastname="Magalhaes Birnbaum" birthdate="2009-05-14" gender="F" nation="BRA" license="399684" swrid="5653298" athleteid="1488" externalid="399684">
              <RESULTS>
                <RESULT eventid="1085" points="352" swimtime="00:01:11.14" resultid="1489" heatid="1990" lane="8" entrytime="00:01:12.10" entrycourse="SCM" />
                <RESULT eventid="1077" points="310" swimtime="00:00:37.28" resultid="1490" heatid="1981" lane="5" entrytime="00:00:43.20" entrycourse="SCM" />
                <RESULT eventid="1127" points="361" swimtime="00:00:32.18" resultid="1491" heatid="2010" lane="6" entrytime="00:00:32.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17325" nation="BRA" region="PR" clubid="1236" name="Colégio Estadual Sagrada Família, Campo Largo" shortname="Clar-Sagrada Fami,Ce">
          <ATHLETES>
            <ATHLETE firstname="Vitor" lastname="Ferreira Rais" birthdate="2007-04-07" gender="M" nation="BRA" license="V387152" swrid="5697227" athleteid="1237" externalid="V387152">
              <RESULTS>
                <RESULT eventid="1081" points="360" swimtime="00:01:03.01" resultid="1238" heatid="1984" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="386" swimtime="00:00:27.67" resultid="1239" heatid="2012" lane="2" />
                <RESULT eventid="1187" points="304" swimtime="00:00:32.34" resultid="1240" heatid="2039" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Guilherme Ballatka" birthdate="2007-06-24" gender="M" nation="BRA" license="398616" swrid="5697228" athleteid="1241" externalid="398616">
              <RESULTS>
                <RESULT eventid="1073" points="390" swimtime="00:00:30.26" resultid="1242" heatid="1979" lane="5" entrytime="00:00:30.87" entrycourse="SCM" />
                <RESULT eventid="1131" points="431" swimtime="00:00:26.67" resultid="1243" heatid="2016" lane="2" entrytime="00:00:27.17" entrycourse="SCM" />
                <RESULT eventid="1171" points="377" swimtime="00:01:06.85" resultid="1244" heatid="2033" lane="8" entrytime="00:01:10.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2647" nation="BRA" region="PR" clubid="1856" name="Colégio Sepam, Ponta Grossa" shortname="Pgro-Sepam,C">
          <ATHLETES>
            <ATHLETE firstname="Felipe" lastname="Chi Kravchychyn" birthdate="2009-09-27" gender="M" nation="BRA" license="344268" swrid="5600134" athleteid="1857" externalid="344268">
              <RESULTS>
                <RESULT eventid="1097" points="463" swimtime="00:00:32.23" resultid="1858" heatid="1996" lane="2" entrytime="00:00:32.19" entrycourse="SCM" />
                <RESULT eventid="1123" points="519" swimtime="00:02:29.50" resultid="1859" heatid="2007" lane="5" entrytime="00:02:27.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:11.94" />
                    <SPLIT distance="150" swimtime="00:01:50.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="482" swimtime="00:04:59.45" resultid="1860" heatid="2025" lane="5" entrytime="00:04:53.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:08.17" />
                    <SPLIT distance="150" swimtime="00:01:48.54" />
                    <SPLIT distance="200" swimtime="00:02:28.42" />
                    <SPLIT distance="250" swimtime="00:03:09.64" />
                    <SPLIT distance="300" swimtime="00:03:51.26" />
                    <SPLIT distance="350" swimtime="00:04:25.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Campagnoli" birthdate="2009-04-13" gender="F" nation="BRA" license="366915" swrid="5600128" athleteid="1861" externalid="366915">
              <RESULTS>
                <RESULT eventid="1077" points="416" swimtime="00:00:33.81" resultid="1862" heatid="1982" lane="6" entrytime="00:00:32.73" entrycourse="SCM" />
                <RESULT eventid="1127" points="453" swimtime="00:00:29.85" resultid="1863" heatid="2011" lane="3" entrytime="00:00:29.31" entrycourse="SCM" />
                <RESULT eventid="1167" points="418" swimtime="00:01:13.36" resultid="1864" heatid="2031" lane="6" entrytime="00:01:13.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2273" nation="BRA" region="PR" clubid="1772" name="Colégio Marista, Maringá" shortname="Mrga-Marista,C">
          <ATHLETES>
            <ATHLETE firstname="Carina" lastname="Costa Profeta" birthdate="2008-03-20" gender="F" nation="BRA" license="366964" swrid="5591584" athleteid="1773" externalid="366964">
              <RESULTS>
                <RESULT eventid="1101" points="502" swimtime="00:00:35.68" resultid="1774" heatid="1998" lane="4" entrytime="00:00:35.51" entrycourse="SCM" />
                <RESULT eventid="1119" points="413" swimtime="00:03:00.64" resultid="1775" heatid="2005" lane="3" entrytime="00:02:52.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                    <SPLIT distance="100" swimtime="00:01:24.77" />
                    <SPLIT distance="150" swimtime="00:02:11.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="461" swimtime="00:01:20.71" resultid="1776" heatid="2042" lane="4" entrytime="00:01:17.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16003" nation="BRA" region="PR" clubid="1591" name="Colégio Saber, Curitiba" shortname="Ctba-Saber,C">
          <ATHLETES>
            <ATHLETE firstname="Bruna" lastname="Bussmann" birthdate="2007-01-16" gender="F" nation="BRA" license="313781" swrid="5579983" athleteid="1592" externalid="313781">
              <RESULTS>
                <RESULT eventid="1069" status="WDR" swimtime="00:00:00.00" resultid="1593" entrytime="00:02:33.56" entrycourse="SCM" />
                <RESULT eventid="1119" status="WDR" swimtime="00:00:00.00" resultid="1594" />
                <RESULT eventid="1183" status="WDR" swimtime="00:00:00.00" resultid="1595" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Francisco Saldo" birthdate="2007-01-23" gender="M" nation="BRA" license="313537" swrid="5600169" athleteid="1596" externalid="313537">
              <RESULTS>
                <RESULT eventid="1089" status="WDR" swimtime="00:00:00.00" resultid="1597" />
                <RESULT eventid="1147" status="WDR" swimtime="00:00:00.00" resultid="1598" />
                <RESULT eventid="1155" status="WDR" swimtime="00:00:00.00" resultid="1599" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13983" nation="BRA" region="PR" clubid="1586" name="Colégio Positivo Vicente Machado, Curitiba" shortname="Ctba-Posi. Vicente,C">
          <ATHLETES>
            <ATHLETE firstname="Caio" lastname="Rocha Silva" birthdate="2007-10-10" gender="M" nation="BRA" license="372280" swrid="5717294" athleteid="1587" externalid="372280">
              <RESULTS>
                <RESULT eventid="1081" status="WDR" swimtime="00:00:00.00" resultid="1588" entrytime="00:00:50.69" entrycourse="SCM" />
                <RESULT eventid="1131" status="WDR" swimtime="00:00:00.00" resultid="1589" entrytime="00:00:23.61" entrycourse="SCM" />
                <RESULT eventid="1179" status="WDR" swimtime="00:00:00.00" resultid="1590" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18915" nation="BRA" region="PR" clubid="1719" name="CCM Tarquino Santos, Foz Do Iguaçu" shortname="Fozi-Tarq.Santos,CCM">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Eduarda Targat Pinheiro" birthdate="2008-09-04" gender="F" nation="BRA" license="331610" swrid="5596894" athleteid="1720" externalid="331610" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1061" points="483" swimtime="00:10:08.14" resultid="1721" heatid="1975" lane="5" entrytime="00:10:09.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                    <SPLIT distance="100" swimtime="00:01:09.71" />
                    <SPLIT distance="150" swimtime="00:01:47.47" />
                    <SPLIT distance="200" swimtime="00:02:24.76" />
                    <SPLIT distance="250" swimtime="00:03:02.54" />
                    <SPLIT distance="300" swimtime="00:03:40.40" />
                    <SPLIT distance="350" swimtime="00:04:19.13" />
                    <SPLIT distance="400" swimtime="00:04:57.50" />
                    <SPLIT distance="450" swimtime="00:05:36.61" />
                    <SPLIT distance="500" swimtime="00:06:16.29" />
                    <SPLIT distance="550" swimtime="00:06:56.51" />
                    <SPLIT distance="600" swimtime="00:07:35.73" />
                    <SPLIT distance="650" swimtime="00:08:14.39" />
                    <SPLIT distance="700" swimtime="00:08:54.24" />
                    <SPLIT distance="750" swimtime="00:09:33.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="421" swimtime="00:05:45.28" resultid="1722" heatid="2024" lane="5" entrytime="00:05:41.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                    <SPLIT distance="100" swimtime="00:01:14.91" />
                    <SPLIT distance="150" swimtime="00:02:00.61" />
                    <SPLIT distance="200" swimtime="00:02:43.01" />
                    <SPLIT distance="250" swimtime="00:03:34.30" />
                    <SPLIT distance="300" swimtime="00:04:27.09" />
                    <SPLIT distance="350" swimtime="00:05:06.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" points="450" swimtime="00:19:44.51" resultid="1723" heatid="2047" lane="5" entrytime="00:20:01.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                    <SPLIT distance="100" swimtime="00:01:12.13" />
                    <SPLIT distance="150" swimtime="00:01:49.70" />
                    <SPLIT distance="200" swimtime="00:02:26.84" />
                    <SPLIT distance="250" swimtime="00:03:04.46" />
                    <SPLIT distance="300" swimtime="00:03:42.05" />
                    <SPLIT distance="350" swimtime="00:04:21.23" />
                    <SPLIT distance="400" swimtime="00:05:01.18" />
                    <SPLIT distance="450" swimtime="00:05:40.15" />
                    <SPLIT distance="500" swimtime="00:06:20.15" />
                    <SPLIT distance="550" swimtime="00:07:00.45" />
                    <SPLIT distance="600" swimtime="00:07:39.59" />
                    <SPLIT distance="650" swimtime="00:08:20.46" />
                    <SPLIT distance="700" swimtime="00:08:59.95" />
                    <SPLIT distance="750" swimtime="00:09:40.65" />
                    <SPLIT distance="800" swimtime="00:10:21.77" />
                    <SPLIT distance="850" swimtime="00:11:01.49" />
                    <SPLIT distance="900" swimtime="00:11:42.62" />
                    <SPLIT distance="950" swimtime="00:12:22.97" />
                    <SPLIT distance="1000" swimtime="00:13:02.87" />
                    <SPLIT distance="1050" swimtime="00:13:43.17" />
                    <SPLIT distance="1100" swimtime="00:14:24.11" />
                    <SPLIT distance="1150" swimtime="00:15:04.90" />
                    <SPLIT distance="1200" swimtime="00:15:45.87" />
                    <SPLIT distance="1250" swimtime="00:16:26.31" />
                    <SPLIT distance="1300" swimtime="00:17:08.09" />
                    <SPLIT distance="1350" swimtime="00:17:47.12" />
                    <SPLIT distance="1400" swimtime="00:18:26.71" />
                    <SPLIT distance="1450" swimtime="00:19:07.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18913" nation="BRA" region="PR" clubid="1886" name="CCM Sebastião Paraná, Palmas" shortname="Pmas-Sebastiã.Pr,CCM">
          <ATHLETES>
            <ATHLETE firstname="Lohan" lastname="Henrique Oliveira" birthdate="2009-03-13" gender="M" nation="BRA" license="410110" athleteid="1887" externalid="410110">
              <RESULTS>
                <RESULT eventid="1081" points="231" swimtime="00:01:12.98" resultid="1888" heatid="1984" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="237" swimtime="00:00:32.55" resultid="1889" heatid="2015" lane="8" entrytime="00:00:32.39" entrycourse="SCM" />
                <RESULT eventid="1179" points="215" swimtime="00:02:45.74" resultid="1890" heatid="2035" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="100" swimtime="00:01:18.13" />
                    <SPLIT distance="150" swimtime="00:02:02.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18903" nation="BRA" region="PR" clubid="1895" name="Colégio Adventista Centro, São José Dos Pinhais" shortname="Sjpi-Adven.Centro,C">
          <ATHLETES>
            <ATHLETE firstname="Ana" lastname="Luiza Rimbano De Jesus" birthdate="2008-09-02" gender="F" nation="BRA" license="366819" swrid="5653297" athleteid="1896" externalid="366819">
              <RESULTS>
                <RESULT eventid="1085" points="539" swimtime="00:01:01.71" resultid="1897" heatid="1990" lane="5" entrytime="00:01:04.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="526" swimtime="00:00:28.40" resultid="1898" heatid="2011" lane="5" entrytime="00:00:29.16" entrycourse="SCM" />
                <RESULT eventid="1175" points="473" swimtime="00:02:21.54" resultid="1899" heatid="2034" lane="4" entrytime="00:02:25.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:07.84" />
                    <SPLIT distance="150" swimtime="00:01:44.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3727" nation="BRA" region="PR" clubid="1917" name="Colégio Estadual Dario Vellozo, Toledo" shortname="Tole-Dario Vello.,Ce">
          <ATHLETES>
            <ATHLETE firstname="Pedro" lastname="Feder" birthdate="2008-11-13" gender="M" nation="BRA" license="347224" swrid="5622278" athleteid="1918" externalid="347224">
              <RESULTS>
                <RESULT eventid="1073" points="380" swimtime="00:00:30.51" resultid="1919" heatid="1979" lane="4" entrytime="00:00:29.80" entrycourse="SCM" />
                <RESULT eventid="1171" points="385" swimtime="00:01:06.41" resultid="1920" heatid="2033" lane="3" entrytime="00:01:05.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="391" swimtime="00:00:29.74" resultid="1921" heatid="2041" lane="1" entrytime="00:00:28.87" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1921" nation="BRA" region="PR" clubid="1794" name="Colégio Objetivo, Maringá" shortname="Mrga-Objetivo,C">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Paiva Boeing" birthdate="2008-01-22" gender="F" nation="BRA" license="318185" swrid="5603884" athleteid="1795" externalid="318185">
              <RESULTS>
                <RESULT eventid="1101" points="342" swimtime="00:00:40.54" resultid="1796" heatid="1998" lane="6" entrytime="00:00:39.57" entrycourse="SCM" />
                <RESULT eventid="1127" points="386" swimtime="00:00:31.49" resultid="1797" heatid="2011" lane="1" entrytime="00:00:29.72" entrycourse="SCM" />
                <RESULT eventid="1183" points="330" swimtime="00:00:35.28" resultid="1798" heatid="2038" lane="3" entrytime="00:00:33.73" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Biason Santana" birthdate="2009-01-21" gender="M" nation="BRA" license="366969" swrid="5317765" athleteid="1799" externalid="366969">
              <RESULTS>
                <RESULT eventid="1089" points="368" swimtime="00:02:28.99" resultid="1800" heatid="1991" lane="2" entrytime="00:02:30.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:11.27" />
                    <SPLIT distance="150" swimtime="00:01:50.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1147" points="407" swimtime="00:01:04.43" resultid="1801" heatid="2023" lane="1" entrytime="00:01:03.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1187" points="461" swimtime="00:00:28.15" resultid="1802" heatid="2041" lane="8" entrytime="00:00:29.07" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17693" nation="BRA" region="PR" clubid="1922" name="7º Colégio Da Polícia Militar, União Da Vitória" shortname="Unvt-7ºcpm,C">
          <ATHLETES>
            <ATHLETE firstname="Pietra" lastname="Cotosky Roveda" birthdate="2009-07-11" gender="F" nation="BRA" license="V399609" athleteid="1923" externalid="V399609">
              <RESULTS>
                <RESULT eventid="1061" points="330" swimtime="00:11:30.66" resultid="1924" heatid="1975" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:17.31" />
                    <SPLIT distance="150" swimtime="00:01:59.50" />
                    <SPLIT distance="200" swimtime="00:02:42.74" />
                    <SPLIT distance="250" swimtime="00:03:26.80" />
                    <SPLIT distance="300" swimtime="00:04:11.00" />
                    <SPLIT distance="350" swimtime="00:04:55.28" />
                    <SPLIT distance="400" swimtime="00:05:39.93" />
                    <SPLIT distance="450" swimtime="00:06:23.34" />
                    <SPLIT distance="500" swimtime="00:07:07.50" />
                    <SPLIT distance="550" swimtime="00:07:52.02" />
                    <SPLIT distance="600" swimtime="00:08:36.22" />
                    <SPLIT distance="650" swimtime="00:09:21.34" />
                    <SPLIT distance="700" swimtime="00:10:07.15" />
                    <SPLIT distance="750" swimtime="00:10:52.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" status="DSQ" swimtime="00:03:02.25" resultid="1925" heatid="2018" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.30" />
                    <SPLIT distance="100" swimtime="00:01:27.70" />
                    <SPLIT distance="150" swimtime="00:02:15.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" points="330" swimtime="00:21:54.00" resultid="1926" heatid="2047" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                    <SPLIT distance="100" swimtime="00:01:15.89" />
                    <SPLIT distance="150" swimtime="00:01:57.97" />
                    <SPLIT distance="200" swimtime="00:02:40.88" />
                    <SPLIT distance="250" swimtime="00:03:23.39" />
                    <SPLIT distance="300" swimtime="00:04:06.64" />
                    <SPLIT distance="350" swimtime="00:04:50.56" />
                    <SPLIT distance="400" swimtime="00:05:21.63" />
                    <SPLIT distance="450" swimtime="00:06:18.97" />
                    <SPLIT distance="500" swimtime="00:07:03.34" />
                    <SPLIT distance="550" swimtime="00:07:47.74" />
                    <SPLIT distance="600" swimtime="00:08:32.50" />
                    <SPLIT distance="650" swimtime="00:09:17.19" />
                    <SPLIT distance="700" swimtime="00:10:01.33" />
                    <SPLIT distance="750" swimtime="00:10:45.56" />
                    <SPLIT distance="800" swimtime="00:11:30.72" />
                    <SPLIT distance="850" swimtime="00:12:15.95" />
                    <SPLIT distance="900" swimtime="00:13:00.27" />
                    <SPLIT distance="950" swimtime="00:13:45.77" />
                    <SPLIT distance="1000" swimtime="00:14:30.43" />
                    <SPLIT distance="1050" swimtime="00:15:16.36" />
                    <SPLIT distance="1100" swimtime="00:16:01.46" />
                    <SPLIT distance="1150" swimtime="00:16:45.40" />
                    <SPLIT distance="1200" swimtime="00:17:31.23" />
                    <SPLIT distance="1250" swimtime="00:18:16.44" />
                    <SPLIT distance="1300" swimtime="00:19:01.35" />
                    <SPLIT distance="1350" swimtime="00:19:45.86" />
                    <SPLIT distance="1400" swimtime="00:20:31.50" />
                    <SPLIT distance="1450" swimtime="00:21:15.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4575" nation="BRA" region="PR" clubid="1710" name="Colégio Monjolo, Foz Do Iguaçu" shortname="Fozi-Monjolo,C">
          <ATHLETES>
            <ATHLETE firstname="Geórgia" lastname="Adeli Jesus" birthdate="2008-03-27" gender="F" nation="BRA" license="312649" swrid="5596864" athleteid="1711" externalid="312649">
              <RESULTS>
                <RESULT eventid="1061" points="357" swimtime="00:11:12.65" resultid="1712" heatid="1975" lane="6" entrytime="00:10:56.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:16.04" />
                    <SPLIT distance="150" swimtime="00:01:55.03" />
                    <SPLIT distance="200" swimtime="00:02:35.89" />
                    <SPLIT distance="250" swimtime="00:03:18.07" />
                    <SPLIT distance="300" swimtime="00:04:00.79" />
                    <SPLIT distance="350" swimtime="00:04:43.55" />
                    <SPLIT distance="400" swimtime="00:05:26.67" />
                    <SPLIT distance="450" swimtime="00:06:09.41" />
                    <SPLIT distance="500" swimtime="00:06:52.21" />
                    <SPLIT distance="550" swimtime="00:07:35.30" />
                    <SPLIT distance="600" swimtime="00:08:19.16" />
                    <SPLIT distance="650" swimtime="00:09:03.60" />
                    <SPLIT distance="700" swimtime="00:09:46.71" />
                    <SPLIT distance="750" swimtime="00:10:30.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="366" swimtime="00:05:23.35" resultid="1713" heatid="2002" lane="2" entrytime="00:05:11.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:13.55" />
                    <SPLIT distance="150" swimtime="00:01:53.24" />
                    <SPLIT distance="200" swimtime="00:02:34.35" />
                    <SPLIT distance="250" swimtime="00:03:16.85" />
                    <SPLIT distance="300" swimtime="00:03:59.07" />
                    <SPLIT distance="350" swimtime="00:04:41.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" status="WDR" swimtime="00:00:00.00" resultid="1714" heatid="2046" lane="4" entrytime="00:21:19.63" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yago" lastname="Simon Pires" birthdate="2008-10-29" gender="M" nation="BRA" license="328942" swrid="5596939" athleteid="1715" externalid="328942">
              <RESULTS>
                <RESULT eventid="1081" points="431" swimtime="00:00:59.33" resultid="1716" heatid="1986" lane="5" entrytime="00:00:58.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="402" swimtime="00:00:27.31" resultid="1717" heatid="2016" lane="5" entrytime="00:00:26.58" entrycourse="SCM" />
                <RESULT eventid="1195" points="322" swimtime="00:01:20.65" resultid="1718" heatid="2044" lane="3" entrytime="00:01:20.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="799" nation="BRA" region="PR" clubid="1777" name="Colégio Mater Dei, Maringá" shortname="Mrga-Mater Dei,C">
          <ATHLETES>
            <ATHLETE firstname="Andressa" lastname="Zamarian Gouvea" birthdate="2007-09-18" gender="F" nation="BRA" license="318503" swrid="5603929" athleteid="1778" externalid="318503">
              <RESULTS>
                <RESULT eventid="1077" points="376" swimtime="00:00:34.98" resultid="1779" heatid="1982" lane="7" entrytime="00:00:35.52" entrycourse="SCM" />
                <RESULT eventid="1135" points="362" swimtime="00:02:46.86" resultid="1780" heatid="2018" lane="3" entrytime="00:02:43.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                    <SPLIT distance="100" swimtime="00:01:20.48" />
                    <SPLIT distance="150" swimtime="00:02:03.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="385" swimtime="00:05:17.92" resultid="1781" heatid="2002" lane="7" entrytime="00:05:16.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.86" />
                    <SPLIT distance="100" swimtime="00:01:16.11" />
                    <SPLIT distance="150" swimtime="00:01:56.48" />
                    <SPLIT distance="200" swimtime="00:02:37.02" />
                    <SPLIT distance="250" swimtime="00:03:17.50" />
                    <SPLIT distance="300" swimtime="00:03:58.11" />
                    <SPLIT distance="350" swimtime="00:04:38.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Batista Sanchez" birthdate="2009-05-22" gender="M" nation="BRA" license="370668" swrid="5255779" athleteid="1782" externalid="370668">
              <RESULTS>
                <RESULT eventid="1097" points="384" swimtime="00:00:34.30" resultid="1783" heatid="1995" lane="4" entrytime="00:00:36.01" entrycourse="SCM" />
                <RESULT eventid="1123" points="394" swimtime="00:02:43.87" resultid="1784" heatid="2007" lane="7" entrytime="00:02:41.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.69" />
                    <SPLIT distance="100" swimtime="00:01:17.99" />
                    <SPLIT distance="150" swimtime="00:02:00.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="415" swimtime="00:01:14.09" resultid="1785" heatid="2044" lane="4" entrytime="00:01:16.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Garcia Cavalcante" birthdate="2008-08-11" gender="M" nation="BRA" license="369676" swrid="5603841" athleteid="1786" externalid="369676">
              <RESULTS>
                <RESULT eventid="1105" points="372" swimtime="00:19:37.24" resultid="1787" heatid="1999" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                    <SPLIT distance="100" swimtime="00:01:11.78" />
                    <SPLIT distance="150" swimtime="00:01:49.83" />
                    <SPLIT distance="200" swimtime="00:02:28.20" />
                    <SPLIT distance="250" swimtime="00:03:06.42" />
                    <SPLIT distance="300" swimtime="00:03:45.30" />
                    <SPLIT distance="350" swimtime="00:04:23.65" />
                    <SPLIT distance="400" swimtime="00:05:02.41" />
                    <SPLIT distance="450" swimtime="00:05:41.51" />
                    <SPLIT distance="500" swimtime="00:06:19.54" />
                    <SPLIT distance="550" swimtime="00:06:57.48" />
                    <SPLIT distance="600" swimtime="00:07:35.94" />
                    <SPLIT distance="650" swimtime="00:08:14.55" />
                    <SPLIT distance="700" swimtime="00:08:52.83" />
                    <SPLIT distance="750" swimtime="00:09:31.91" />
                    <SPLIT distance="800" swimtime="00:10:11.17" />
                    <SPLIT distance="850" swimtime="00:10:51.04" />
                    <SPLIT distance="900" swimtime="00:11:30.74" />
                    <SPLIT distance="950" swimtime="00:12:10.49" />
                    <SPLIT distance="1000" swimtime="00:12:50.73" />
                    <SPLIT distance="1050" swimtime="00:13:30.29" />
                    <SPLIT distance="1100" swimtime="00:14:10.50" />
                    <SPLIT distance="1150" swimtime="00:14:51.04" />
                    <SPLIT distance="1200" swimtime="00:15:30.92" />
                    <SPLIT distance="1250" swimtime="00:16:13.08" />
                    <SPLIT distance="1300" swimtime="00:16:54.49" />
                    <SPLIT distance="1350" swimtime="00:17:35.12" />
                    <SPLIT distance="1400" swimtime="00:18:15.69" />
                    <SPLIT distance="1450" swimtime="00:18:57.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1123" points="351" swimtime="00:02:50.25" resultid="1788" heatid="2007" lane="1" entrytime="00:02:41.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                    <SPLIT distance="100" swimtime="00:01:20.37" />
                    <SPLIT distance="150" swimtime="00:02:04.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6517" nation="BRA" region="PR" clubid="1813" name="Colégio Regina Mundi, Maringá" shortname="Mrga-Regina Mundi,C">
          <ATHLETES>
            <ATHLETE firstname="Theodoro" lastname="Marques Serra" birthdate="2009-11-24" gender="M" nation="BRA" license="370661" swrid="5603870" athleteid="1814" externalid="370661">
              <RESULTS>
                <RESULT eventid="1081" points="390" swimtime="00:01:01.36" resultid="1815" heatid="1986" lane="2" entrytime="00:01:00.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="318" swimtime="00:02:34.68" resultid="1816" heatid="2019" lane="5" entrytime="00:02:37.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:14.37" />
                    <SPLIT distance="150" swimtime="00:01:54.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="329" swimtime="00:01:09.99" resultid="1817" heatid="2033" lane="2" entrytime="00:01:09.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15552" nation="BRA" region="PR" clubid="1833" name="Colégio Positivo Master, Ponta Grossa" shortname="Pgro-Positivo.Mast,C">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Carolina Babiuki" birthdate="2007-02-06" gender="F" nation="BRA" license="316227" swrid="5600131" athleteid="1838" externalid="316227" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1077" points="501" swimtime="00:00:31.79" resultid="1839" heatid="1982" lane="3" entrytime="00:00:32.09" entrycourse="SCM" />
                <RESULT eventid="1127" points="519" swimtime="00:00:28.53" resultid="1840" heatid="2011" lane="4" entrytime="00:00:28.97" entrycourse="SCM" />
                <RESULT eventid="1167" points="437" swimtime="00:01:12.31" resultid="1841" heatid="2031" lane="3" entrytime="00:01:10.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Delinski" birthdate="2009-11-28" gender="F" nation="BRA" license="385190" swrid="5600150" athleteid="1842" externalid="385190">
              <RESULTS>
                <RESULT eventid="1101" points="305" swimtime="00:00:42.12" resultid="1843" heatid="1998" lane="2" entrytime="00:00:41.86" entrycourse="SCM" />
                <RESULT eventid="1119" points="255" swimtime="00:03:32.04" resultid="1844" heatid="2005" lane="2" entrytime="00:03:26.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.50" />
                    <SPLIT distance="100" swimtime="00:01:40.10" />
                    <SPLIT distance="150" swimtime="00:02:36.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="264" swimtime="00:01:25.51" resultid="1845" heatid="2030" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fegert" birthdate="2009-04-13" gender="M" nation="BRA" license="353813" swrid="5622279" athleteid="1846" externalid="353813">
              <RESULTS>
                <RESULT eventid="1147" points="390" swimtime="00:01:05.36" resultid="1847" heatid="2022" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" status="DNS" swimtime="00:00:00.00" resultid="1848" heatid="2016" lane="1" entrytime="00:00:27.72" entrycourse="SCM" />
                <RESULT eventid="1187" points="450" swimtime="00:00:28.38" resultid="1849" heatid="2040" lane="4" entrytime="00:00:30.46" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Gueiber Montes" birthdate="2009-03-09" gender="M" nation="BRA" license="342154" swrid="5600179" athleteid="1834" externalid="342154">
              <RESULTS>
                <RESULT eventid="1081" points="516" swimtime="00:00:55.87" resultid="1835" heatid="1987" lane="5" entrytime="00:00:54.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="488" swimtime="00:00:25.59" resultid="1836" heatid="2017" lane="6" entrytime="00:00:25.27" entrycourse="SCM" />
                <RESULT eventid="1171" points="491" swimtime="00:01:01.25" resultid="1837" heatid="2033" lane="5" entrytime="00:01:00.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="PGRO-POS.MASTER,C &apos;&apos;A&apos;&apos;" number="1">
              <RESULTS>
                <RESULT eventid="1109" points="441" swimtime="00:02:04.95" resultid="1850" heatid="2000" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="100" swimtime="00:01:12.23" />
                    <SPLIT distance="150" swimtime="00:01:40.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1838" number="1" />
                    <RELAYPOSITION athleteid="1842" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1846" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1834" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6485" nation="BRA" region="PR" clubid="1260" name="Colégio Integrado, Campo Mourão" shortname="Cmou-Integrado,C">
          <ATHLETES>
            <ATHLETE firstname="Guilherme" lastname="Stipp Silva" birthdate="2009-12-02" gender="M" nation="BRA" license="378462" swrid="5603918" athleteid="1261" externalid="378462">
              <RESULTS>
                <RESULT eventid="1081" points="377" swimtime="00:01:02.03" resultid="1262" heatid="1986" lane="8" entrytime="00:01:03.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" status="DSQ" swimtime="00:00:37.87" resultid="1263" heatid="1995" lane="5" entrytime="00:00:39.01" entrycourse="SCM" />
                <RESULT eventid="1131" points="393" swimtime="00:00:27.52" resultid="1264" heatid="2015" lane="3" entrytime="00:00:29.18" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15551" nation="BRA" region="PR" clubid="1540" name="Colégio Estadual Pedro Macedo, Curitiba" shortname="Ctba-Pedro Macedo,Ce">
          <ATHLETES>
            <ATHLETE firstname="Nicolas" lastname="Mingorance Martins" birthdate="2007-10-13" gender="M" nation="BRA" license="393920" swrid="5622295" athleteid="1549" externalid="393920">
              <RESULTS>
                <RESULT eventid="1081" points="460" swimtime="00:00:58.06" resultid="1550" heatid="1987" lane="8" entrytime="00:00:56.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="278" swimtime="00:00:38.22" resultid="1551" heatid="1994" lane="3" />
                <RESULT eventid="1131" points="437" swimtime="00:00:26.55" resultid="1552" heatid="2017" lane="7" entrytime="00:00:25.71" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="David Cella" birthdate="2008-02-17" gender="M" nation="BRA" license="341107" swrid="5634581" athleteid="1541" externalid="341107">
              <RESULTS>
                <RESULT eventid="1081" points="588" swimtime="00:00:53.52" resultid="1542" heatid="1987" lane="6" entrytime="00:00:54.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="499" swimtime="00:00:31.45" resultid="1543" heatid="1996" lane="5" entrytime="00:00:30.47" entrycourse="SCM" />
                <RESULT eventid="1131" points="549" swimtime="00:00:24.62" resultid="1544" heatid="2017" lane="4" entrytime="00:00:24.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Krupacz" birthdate="2008-04-18" gender="F" nation="BRA" license="329187" swrid="5634611" athleteid="1545" externalid="329187">
              <RESULTS>
                <RESULT eventid="1077" points="531" swimtime="00:00:31.17" resultid="1546" heatid="1982" lane="4" entrytime="00:00:30.70" entrycourse="SCM" />
                <RESULT eventid="1111" points="519" swimtime="00:04:47.80" resultid="1547" heatid="2002" lane="3" entrytime="00:04:47.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                    <SPLIT distance="100" swimtime="00:01:08.10" />
                    <SPLIT distance="150" swimtime="00:01:43.48" />
                    <SPLIT distance="200" swimtime="00:02:19.05" />
                    <SPLIT distance="250" swimtime="00:02:55.55" />
                    <SPLIT distance="300" swimtime="00:03:32.81" />
                    <SPLIT distance="350" swimtime="00:04:10.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="572" swimtime="00:01:06.11" resultid="1548" heatid="2031" lane="4" entrytime="00:01:06.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="10585" nation="BRA" region="PR" clubid="1615" name="Colégio Estadual Santa Cândida, Curitiba" shortname="Ctba-Stª. Candida,Ce">
          <ATHLETES>
            <ATHLETE firstname="Carlos" lastname="Alexandre Azevedo" birthdate="2008-05-20" gender="M" nation="BRA" license="398694" swrid="5717240" athleteid="1616" externalid="398694">
              <RESULTS>
                <RESULT eventid="1097" points="209" swimtime="00:00:41.99" resultid="1617" heatid="1995" lane="3" entrytime="00:00:43.48" entrycourse="SCM" />
                <RESULT eventid="1131" points="270" swimtime="00:00:31.18" resultid="1618" heatid="2015" lane="1" entrytime="00:00:30.98" entrycourse="SCM" />
                <RESULT eventid="1195" points="213" swimtime="00:01:32.44" resultid="1619" heatid="2044" lane="2" entrytime="00:01:35.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13348" nation="BRA" region="PR" clubid="1610" name="Colégio Sesi CIC, Curitiba" shortname="Ctba-Sesi CIC,C">
          <ATHLETES>
            <ATHLETE firstname="Giulia" lastname="Quignalia Goncalves" birthdate="2008-04-15" gender="F" nation="BRA" license="V414492" athleteid="1611" externalid="V414492">
              <RESULTS>
                <RESULT eventid="1061" points="218" swimtime="00:13:12.70" resultid="1612" heatid="1975" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                    <SPLIT distance="150" swimtime="00:02:13.69" />
                    <SPLIT distance="200" swimtime="00:03:03.57" />
                    <SPLIT distance="250" swimtime="00:03:54.40" />
                    <SPLIT distance="300" swimtime="00:04:45.52" />
                    <SPLIT distance="350" swimtime="00:05:37.24" />
                    <SPLIT distance="400" swimtime="00:06:28.64" />
                    <SPLIT distance="450" swimtime="00:07:19.77" />
                    <SPLIT distance="500" swimtime="00:08:11.45" />
                    <SPLIT distance="550" swimtime="00:09:02.38" />
                    <SPLIT distance="600" swimtime="00:09:53.40" />
                    <SPLIT distance="650" swimtime="00:10:43.50" />
                    <SPLIT distance="700" swimtime="00:11:34.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="220" swimtime="00:06:23.09" resultid="1613" heatid="2001" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:01:23.78" />
                    <SPLIT distance="150" swimtime="00:02:12.57" />
                    <SPLIT distance="200" swimtime="00:03:04.31" />
                    <SPLIT distance="250" swimtime="00:03:55.70" />
                    <SPLIT distance="300" swimtime="00:04:46.37" />
                    <SPLIT distance="350" swimtime="00:05:36.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1199" points="214" swimtime="00:25:16.43" resultid="1614" heatid="2047" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                    <SPLIT distance="100" swimtime="00:01:29.22" />
                    <SPLIT distance="150" swimtime="00:02:17.67" />
                    <SPLIT distance="200" swimtime="00:03:08.59" />
                    <SPLIT distance="250" swimtime="00:04:00.32" />
                    <SPLIT distance="300" swimtime="00:04:52.03" />
                    <SPLIT distance="350" swimtime="00:05:42.94" />
                    <SPLIT distance="400" swimtime="00:06:34.19" />
                    <SPLIT distance="450" swimtime="00:07:25.58" />
                    <SPLIT distance="500" swimtime="00:08:17.02" />
                    <SPLIT distance="550" swimtime="00:09:09.68" />
                    <SPLIT distance="600" swimtime="00:10:00.81" />
                    <SPLIT distance="650" swimtime="00:10:52.26" />
                    <SPLIT distance="700" swimtime="00:11:43.69" />
                    <SPLIT distance="750" swimtime="00:12:35.03" />
                    <SPLIT distance="800" swimtime="00:13:26.92" />
                    <SPLIT distance="850" swimtime="00:14:18.53" />
                    <SPLIT distance="900" swimtime="00:15:09.48" />
                    <SPLIT distance="950" swimtime="00:16:01.46" />
                    <SPLIT distance="1000" swimtime="00:16:52.64" />
                    <SPLIT distance="1050" swimtime="00:17:44.01" />
                    <SPLIT distance="1100" swimtime="00:18:35.71" />
                    <SPLIT distance="1150" swimtime="00:19:26.77" />
                    <SPLIT distance="1200" swimtime="00:20:17.91" />
                    <SPLIT distance="1250" swimtime="00:21:08.96" />
                    <SPLIT distance="1300" swimtime="00:21:59.79" />
                    <SPLIT distance="1350" swimtime="00:22:49.52" />
                    <SPLIT distance="1400" swimtime="00:23:39.52" />
                    <SPLIT distance="1450" swimtime="00:24:29.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18933" nation="BRA" region="PR" clubid="1645" name="Colégio Estadual Jardim Santa Cruz, Cascavel" shortname="Cvel-Jardim Santa,Ce">
          <ATHLETES>
            <ATHLETE firstname="Isis" lastname="Emanuele Balan Da Silva" birthdate="2009-01-30" gender="F" nation="BRA" license="V414483" athleteid="1646" externalid="V414483">
              <RESULTS>
                <RESULT eventid="1085" points="147" swimtime="00:01:35.14" resultid="1647" heatid="1988" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="127" reactiontime="+57" swimtime="00:00:50.17" resultid="1648" heatid="1981" lane="8" />
                <RESULT eventid="1127" points="168" swimtime="00:00:41.54" resultid="1649" heatid="2009" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17296" nation="BRA" region="PR" clubid="1250" name="Colégio Nossa Sra. Do Rosário, Colombo" shortname="Clbo-N.Sra.Rosário,C">
          <ATHLETES>
            <ATHLETE firstname="Jennifer" lastname="De Abreu" birthdate="2009-11-07" gender="F" nation="BRA" license="356212" swrid="5600144" athleteid="1251" externalid="356212">
              <RESULTS>
                <RESULT eventid="1069" points="377" swimtime="00:02:48.63" resultid="1252" heatid="1977" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="100" swimtime="00:01:18.13" />
                    <SPLIT distance="150" swimtime="00:02:08.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="440" swimtime="00:00:30.14" resultid="1253" heatid="2011" lane="7" entrytime="00:00:29.61" entrycourse="SCM" />
                <RESULT eventid="1183" points="434" swimtime="00:00:32.20" resultid="1254" heatid="2037" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3725" nation="BRA" region="PR" clubid="1738" name="Colégio Sagrada Família, Mandaguari" shortname="Mdri-Sagrada Fami.,C">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Isabel Henriques" birthdate="2007-09-05" gender="F" nation="BRA" license="V414491" athleteid="1739" externalid="V414491">
              <RESULTS>
                <RESULT eventid="1085" points="156" swimtime="00:01:33.16" resultid="1740" heatid="1988" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="127" swimtime="00:00:50.11" resultid="1741" heatid="1981" lane="1" />
                <RESULT eventid="1127" points="169" swimtime="00:00:41.40" resultid="1742" heatid="2008" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15595" nation="BRA" region="PR" clubid="1743" name="Colégio Adventista De Maringá" shortname="Mrga-Adventista,C">
          <ATHLETES>
            <ATHLETE firstname="Rafael" lastname="Quental De Meireles" birthdate="2008-11-20" gender="M" nation="BRA" license="392103" swrid="5603898" athleteid="1744" externalid="392103">
              <RESULTS>
                <RESULT eventid="1147" points="307" swimtime="00:01:10.79" resultid="1745" heatid="2022" lane="5" entrytime="00:01:08.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="339" swimtime="00:00:28.91" resultid="1746" heatid="2015" lane="5" entrytime="00:00:29.02" entrycourse="SCM" />
                <RESULT eventid="1179" points="371" swimtime="00:02:18.28" resultid="1747" heatid="2036" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                    <SPLIT distance="100" swimtime="00:01:04.41" />
                    <SPLIT distance="150" swimtime="00:01:41.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="14743" nation="BRA" region="PR" clubid="1818" name="Colégio Santo Inácio, Maringá" shortname="Mrga-Santo Inácio,C">
          <ATHLETES>
            <ATHLETE firstname="Hammon" lastname="Henrique Costa" birthdate="2008-09-19" gender="M" nation="BRA" license="408703" swrid="5726000" athleteid="1819" externalid="408703">
              <RESULTS>
                <RESULT eventid="1081" status="DNS" swimtime="00:00:00.00" resultid="1820" heatid="1985" lane="4" entrytime="00:01:05.42" entrycourse="SCM" />
                <RESULT eventid="1097" status="DNS" swimtime="00:00:00.00" resultid="1821" heatid="1993" lane="4" />
                <RESULT eventid="1131" status="DNS" swimtime="00:00:00.00" resultid="1822" heatid="2015" lane="2" entrytime="00:00:29.48" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6520" nation="BRA" region="PR" clubid="1876" name="Colégio Estadual Semiramis Barros Braga, Pinhais" shortname="Pin-Semira. Braga,Ce">
          <ATHLETES>
            <ATHLETE firstname="Enzo" lastname="Andreis Ramos" birthdate="2007-03-26" gender="M" nation="BRA" license="406719" swrid="5717243" athleteid="1877" externalid="406719">
              <RESULTS>
                <RESULT eventid="1081" points="360" swimtime="00:01:03.02" resultid="1878" heatid="1985" lane="5" entrytime="00:01:06.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1073" points="222" swimtime="00:00:36.50" resultid="1879" heatid="1979" lane="6" entrytime="00:00:36.91" entrycourse="SCM" />
                <RESULT eventid="1131" points="342" swimtime="00:00:28.81" resultid="1880" heatid="2015" lane="4" entrytime="00:00:28.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2611" nation="BRA" region="PR" clubid="1891" name="Colégio Estadual Hermínia Lupion, Ribeirão Pinhal" shortname="Rpin-Hermínia,Ce">
          <ATHLETES>
            <ATHLETE firstname="Yasmin" lastname="Karoline Gordiano" birthdate="2009-03-19" gender="F" nation="BRA" license="V414484" athleteid="1892" externalid="V414484">
              <RESULTS>
                <RESULT eventid="1135" status="DSQ" swimtime="00:00:00.00" resultid="1893" heatid="2018" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.47" />
                    <SPLIT distance="100" swimtime="00:02:39.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" status="DNS" swimtime="00:00:00.00" resultid="1894" heatid="2034" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6486" nation="BRA" region="PR" clubid="1446" name="Colégio Da Polícia Militar, Curitiba" shortname="Ctba-Cpmpr,C">
          <ATHLETES>
            <ATHLETE firstname="Bernardo" lastname="Casiano Andrade" birthdate="2008-09-22" gender="M" nation="BRA" license="V414512" athleteid="1478" externalid="V414512">
              <RESULTS>
                <RESULT eventid="1097" points="213" swimtime="00:00:41.73" resultid="1479" heatid="1994" lane="1" />
                <RESULT eventid="1131" points="281" swimtime="00:00:30.77" resultid="1480" heatid="2014" lane="7" />
                <RESULT eventid="1195" points="197" swimtime="00:01:34.91" resultid="1481" heatid="2043" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietra" lastname="Olandoski Demori" birthdate="2007-06-23" gender="F" nation="BRA" license="V384323" athleteid="1455" externalid="V384323">
              <RESULTS>
                <RESULT eventid="1085" points="181" swimtime="00:01:28.80" resultid="1456" heatid="1988" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="120" swimtime="00:00:57.48" resultid="1457" heatid="1998" lane="8" />
                <RESULT eventid="1127" points="184" swimtime="00:00:40.31" resultid="1458" heatid="2009" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Akira Oshima" birthdate="2008-08-26" gender="M" nation="BRA" license="V414510" athleteid="1471" externalid="V414510">
              <RESULTS>
                <RESULT eventid="1073" points="218" swimtime="00:00:36.70" resultid="1472" heatid="1978" lane="5" />
                <RESULT eventid="1131" points="309" swimtime="00:00:29.81" resultid="1473" heatid="2014" lane="2" />
                <RESULT eventid="1171" points="187" swimtime="00:01:24.41" resultid="1474" heatid="2032" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Andrianczik Corcini" birthdate="2008-07-19" gender="M" nation="BRA" license="406685" swrid="5736533" athleteid="1459" externalid="406685">
              <RESULTS>
                <RESULT eventid="1081" points="269" swimtime="00:01:09.40" resultid="1460" heatid="1983" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="225" swimtime="00:00:40.99" resultid="1461" heatid="1994" lane="5" />
                <RESULT eventid="1195" points="214" swimtime="00:01:32.35" resultid="1462" heatid="2044" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joshua" lastname="Gomide Capraro" birthdate="2009-01-18" gender="M" nation="BRA" license="339030" swrid="5600177" athleteid="1447" externalid="339030">
              <RESULTS>
                <RESULT eventid="1081" points="521" swimtime="00:00:55.71" resultid="1448" heatid="1987" lane="2" entrytime="00:00:55.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="498" swimtime="00:00:25.42" resultid="1449" heatid="2017" lane="5" entrytime="00:00:24.95" entrycourse="SCM" />
                <RESULT eventid="1179" points="538" swimtime="00:02:02.12" resultid="1450" heatid="2036" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                    <SPLIT distance="100" swimtime="00:00:58.06" />
                    <SPLIT distance="150" swimtime="00:01:29.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hannah" lastname="Do Vale Heinrichs" birthdate="2007-09-13" gender="F" nation="BRA" license="V414493" athleteid="1463" externalid="V414493">
              <RESULTS>
                <RESULT eventid="1077" points="250" swimtime="00:00:40.05" resultid="1464" heatid="1981" lane="2" />
                <RESULT eventid="1127" points="276" swimtime="00:00:35.20" resultid="1465" heatid="2009" lane="8" />
                <RESULT eventid="1167" points="212" swimtime="00:01:31.95" resultid="1466" heatid="2030" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabelly" lastname="Brodbeck Hawthorne" birthdate="2007-05-06" gender="F" nation="BRA" license="V384243" athleteid="1451" externalid="V384243">
              <RESULTS>
                <RESULT eventid="1101" points="169" swimtime="00:00:51.22" resultid="1452" heatid="1997" lane="6" />
                <RESULT eventid="1127" points="285" swimtime="00:00:34.83" resultid="1453" heatid="2009" lane="2" />
                <RESULT eventid="1183" status="WDR" swimtime="00:00:00.00" resultid="1454" heatid="2037" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Meneguete Toledo" birthdate="2009-10-05" gender="F" nation="BRA" license="V414494" athleteid="1467" externalid="V414494">
              <RESULTS>
                <RESULT eventid="1085" points="198" swimtime="00:01:26.20" resultid="1468" heatid="1988" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="115" swimtime="00:00:51.81" resultid="1469" heatid="1980" lane="3" />
                <RESULT eventid="1127" points="214" swimtime="00:00:38.29" resultid="1470" heatid="2009" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Dias Da Cruz Goncalves" birthdate="2007-03-25" gender="M" nation="BRA" license="V414511" athleteid="1475" externalid="V414511">
              <RESULTS>
                <RESULT eventid="1073" points="120" swimtime="00:00:44.71" resultid="1476" heatid="1978" lane="3" />
                <RESULT eventid="1131" points="226" swimtime="00:00:33.06" resultid="1477" heatid="2013" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CTBA-POL. MILITAR,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1161" points="373" swimtime="00:01:53.54" resultid="1484" heatid="2027" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                    <SPLIT distance="100" swimtime="00:00:59.51" />
                    <SPLIT distance="150" swimtime="00:01:28.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1459" number="1" />
                    <RELAYPOSITION athleteid="1471" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1478" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1447" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1203" points="297" swimtime="00:02:14.47" resultid="1485" heatid="2048" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                    <SPLIT distance="100" swimtime="00:01:15.58" />
                    <SPLIT distance="150" swimtime="00:01:45.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1471" number="1" />
                    <RELAYPOSITION athleteid="1459" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1447" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1478" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="CTBA-POL. MILITAR,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1159" points="250" swimtime="00:02:26.68" resultid="1482" heatid="2026" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                    <SPLIT distance="100" swimtime="00:01:18.07" />
                    <SPLIT distance="150" swimtime="00:01:52.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1455" number="1" />
                    <RELAYPOSITION athleteid="1467" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1463" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1451" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1205" points="176" swimtime="00:03:02.60" resultid="1483" heatid="2049" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.39" />
                    <SPLIT distance="100" swimtime="00:01:35.85" />
                    <SPLIT distance="150" swimtime="00:02:24.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1463" number="1" />
                    <RELAYPOSITION athleteid="1455" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1451" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1467" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="CTBA-POL. MILITAR,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1109" points="297" swimtime="00:02:22.53" resultid="1486" heatid="2000" lane="5">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:01:49.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1463" number="1" />
                    <RELAYPOSITION athleteid="1478" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1447" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1451" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="4574" nation="BRA" region="PR" clubid="1673" name="Colégio Estadual Almirante Tamandaré, Fozi" shortname="Fozi-Al.Tamandaré,Ce">
          <ATHLETES>
            <ATHLETE firstname="Matheus" lastname="Rogge" birthdate="2008-09-02" gender="M" nation="BRA" license="383387" swrid="4883279" athleteid="1674" externalid="383387" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1081" points="491" swimtime="00:00:56.80" resultid="1675" heatid="1986" lane="4" entrytime="00:00:56.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1131" points="466" swimtime="00:00:26.00" resultid="1676" heatid="2017" lane="2" entrytime="00:00:25.67" entrycourse="SCM" />
                <RESULT eventid="1171" points="313" swimtime="00:01:11.14" resultid="1677" heatid="2033" lane="6" entrytime="00:01:07.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Mattiello" birthdate="2009-04-11" gender="F" nation="BRA" license="367011" swrid="5596914" athleteid="1678" externalid="367011" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1085" points="392" swimtime="00:01:08.65" resultid="1679" heatid="1990" lane="3" entrytime="00:01:07.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="399" swimtime="00:00:31.14" resultid="1680" heatid="2010" lane="4" entrytime="00:00:30.48" entrycourse="SCM" />
                <RESULT eventid="1175" points="410" swimtime="00:02:28.42" resultid="1681" heatid="2034" lane="3" entrytime="00:02:31.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:13.15" />
                    <SPLIT distance="150" swimtime="00:01:51.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18932" nation="BRA" region="PR" clubid="1535" name="Colégio Estadual Paulo Leminski, Curitiba" shortname="Ctba-P. Leminski,Ce">
          <ATHLETES>
            <ATHLETE firstname="Herick" lastname="Dos Santos" birthdate="2009-06-11" gender="M" nation="BRA" license="406724" swrid="5717258" athleteid="1536" externalid="406724">
              <RESULTS>
                <RESULT eventid="1115" points="168" swimtime="00:06:24.53" resultid="1537" heatid="2003" lane="4" entrytime="00:07:14.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                    <SPLIT distance="100" swimtime="00:01:25.72" />
                    <SPLIT distance="150" swimtime="00:02:15.43" />
                    <SPLIT distance="200" swimtime="00:03:06.46" />
                    <SPLIT distance="250" swimtime="00:03:56.15" />
                    <SPLIT distance="300" swimtime="00:04:46.48" />
                    <SPLIT distance="350" swimtime="00:05:36.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1171" points="101" swimtime="00:01:43.45" resultid="1538" heatid="2032" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1163" points="151" swimtime="00:13:52.24" resultid="1539" heatid="2029" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                    <SPLIT distance="100" swimtime="00:01:28.64" />
                    <SPLIT distance="150" swimtime="00:02:18.88" />
                    <SPLIT distance="200" swimtime="00:03:10.15" />
                    <SPLIT distance="250" swimtime="00:04:03.24" />
                    <SPLIT distance="300" swimtime="00:04:55.87" />
                    <SPLIT distance="350" swimtime="00:05:49.88" />
                    <SPLIT distance="400" swimtime="00:06:44.56" />
                    <SPLIT distance="450" swimtime="00:07:37.73" />
                    <SPLIT distance="500" swimtime="00:08:31.11" />
                    <SPLIT distance="550" swimtime="00:09:24.79" />
                    <SPLIT distance="600" swimtime="00:10:18.10" />
                    <SPLIT distance="650" swimtime="00:11:11.58" />
                    <SPLIT distance="700" swimtime="00:12:06.91" />
                    <SPLIT distance="750" swimtime="00:13:00.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16000" nation="BRA" region="PR" clubid="1789" name="Colégio Nobel, Maringá" shortname="Mrga-Nobel,C">
          <ATHLETES>
            <ATHLETE firstname="Sophia" lastname="Donato De Morais" birthdate="2009-03-28" gender="F" nation="BRA" license="345588" swrid="5485198" athleteid="1790" externalid="345588">
              <RESULTS>
                <RESULT eventid="1077" points="362" swimtime="00:00:35.40" resultid="1791" heatid="1982" lane="2" entrytime="00:00:35.28" entrycourse="SCM" />
                <RESULT eventid="1135" points="362" swimtime="00:02:46.77" resultid="1792" heatid="2018" lane="5" entrytime="00:02:41.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.02" />
                    <SPLIT distance="100" swimtime="00:01:19.65" />
                    <SPLIT distance="150" swimtime="00:02:03.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="371" swimtime="00:01:16.35" resultid="1793" heatid="2031" lane="7" entrytime="00:01:16.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16303" nation="BRA" region="PR" clubid="1497" name="CCM Ermelino De Leão, Curitiba" shortname="Ctba-Ermeli.Leão,CCM">
          <ATHLETES>
            <ATHLETE firstname="Izabelly" lastname="Mendonca Bello" birthdate="2008-04-15" gender="F" nation="BRA" license="376996" swrid="5600217" athleteid="1498" externalid="376996" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1069" points="331" swimtime="00:02:55.99" resultid="1499" heatid="1977" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.65" />
                    <SPLIT distance="100" swimtime="00:01:25.68" />
                    <SPLIT distance="150" swimtime="00:02:14.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="352" swimtime="00:03:10.46" resultid="1500" heatid="2005" lane="6" entrytime="00:03:06.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                    <SPLIT distance="100" swimtime="00:01:30.35" />
                    <SPLIT distance="150" swimtime="00:02:20.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1191" points="398" swimtime="00:01:24.77" resultid="1501" heatid="2042" lane="2" entrytime="00:01:27.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15570" nation="BRA" region="PR" clubid="1379" name="Colégio Bom Jesus Seminário, Curitiba" shortname="Ctba-Bj Seminário,C">
          <ATHLETES>
            <ATHLETE firstname="Pedro" lastname="Servienski Silva" birthdate="2009-09-10" gender="M" nation="BRA" license="V383395" athleteid="1384" externalid="V383395">
              <RESULTS>
                <RESULT eventid="1097" points="214" swimtime="00:00:41.69" resultid="1385" heatid="1995" lane="2" entrytime="00:00:46.41" entrycourse="SCM" />
                <RESULT eventid="1131" points="254" swimtime="00:00:31.81" resultid="1386" heatid="2014" lane="4" entrytime="00:00:32.91" entrycourse="SCM" />
                <RESULT eventid="1195" status="DSQ" swimtime="00:01:37.24" resultid="1387" heatid="2044" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicole" lastname="Crestani Nunes" birthdate="2008-12-15" gender="F" nation="BRA" license="V414479" athleteid="1388" externalid="V414479">
              <RESULTS>
                <RESULT eventid="1085" status="DNS" swimtime="00:00:00.00" resultid="1389" heatid="1989" lane="8" />
                <RESULT eventid="1077" status="DNS" swimtime="00:00:00.00" resultid="1390" heatid="1980" lane="7" />
                <RESULT eventid="1127" status="DNS" swimtime="00:00:00.00" resultid="1391" heatid="2008" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ferreira Motta" birthdate="2008-10-24" gender="M" nation="BRA" license="378068" swrid="5600160" athleteid="1380" externalid="378068">
              <RESULTS>
                <RESULT eventid="1081" points="392" swimtime="00:01:01.23" resultid="1381" heatid="1986" lane="6" entrytime="00:01:00.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="372" swimtime="00:00:34.68" resultid="1382" heatid="1996" lane="1" entrytime="00:00:33.03" entrycourse="SCM" />
                <RESULT eventid="1131" points="364" swimtime="00:00:28.23" resultid="1383" heatid="2016" lane="8" entrytime="00:00:28.04" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="10546" nation="BRA" region="PR" clubid="1553" name="Colégio Positivo Jardim Ambiental, Curitiba" shortname="Ctba-Posi. Ambien.,C">
          <ATHLETES>
            <ATHLETE firstname="Marcus" lastname="Vinicius De Almeida" birthdate="2009-06-16" gender="M" nation="BRA" license="348099" swrid="5600272" athleteid="1554" externalid="348099">
              <RESULTS>
                <RESULT eventid="1097" points="455" swimtime="00:00:32.43" resultid="1555" heatid="1996" lane="7" entrytime="00:00:32.37" entrycourse="SCM" />
                <RESULT eventid="1123" points="436" swimtime="00:02:38.35" resultid="1556" heatid="2006" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:01:14.73" />
                    <SPLIT distance="150" swimtime="00:01:56.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="489" swimtime="00:01:10.13" resultid="1557" heatid="2045" lane="2" entrytime="00:01:11.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
