<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.79567">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Curitiba" name="Troféu Ossami Fukuda (Pré-Mirim/Petiz) 2024" course="LCM" deadline="2024-05-20" entrystartdate="2024-05-14" entrytype="INVITATION" hostclub="Clube Curitibano" hostclub.url="https://clubecuritibano.com.br/" number="38308" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/evento/natacao/38308/" startmethod="1" timing="AUTOMATIC" touchpad="BOTHSIDE" masters="F" withdrawuntil="2024-05-22" state="PR" nation="BRA">
      <AGEDATE value="2024-05-24" type="YEAR" />
      <POOL name="Parque Aquático do Clube Curitibano" lanemin="1" lanemax="8" />
      <FACILITY city="Curitiba" name="Parque Aquático do Clube Curitibano" nation="BRA" state="PR" street="Avenida Presidente Getúlio Vargas, 2857" street2="Água Verde" zip="80240-040" />
      <POINTTABLE pointtableid="3017" name="FINA Point Scoring" version="2024" />
      <QUALIFY from="2023-05-24" until="2024-05-23" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-05-24" daytime="08:40" endtime="12:02" number="1" officialmeeting="08:00" warmupfrom="07:30" warmupuntil="08:30">
          <EVENTS>
            <EVENT eventid="1062" daytime="08:40" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1063" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2566" />
                    <RANKING order="2" place="2" resultid="2377" />
                    <RANKING order="3" place="3" resultid="1867" />
                    <RANKING order="4" place="4" resultid="2367" />
                    <RANKING order="5" place="5" resultid="1937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1832" />
                    <RANKING order="2" place="2" resultid="1773" />
                    <RANKING order="3" place="3" resultid="1718" />
                    <RANKING order="4" place="4" resultid="1678" />
                    <RANKING order="5" place="5" resultid="1683" />
                    <RANKING order="6" place="6" resultid="1738" />
                    <RANKING order="7" place="7" resultid="1763" />
                    <RANKING order="8" place="8" resultid="1463" />
                    <RANKING order="9" place="9" resultid="2342" />
                    <RANKING order="10" place="-1" resultid="1246" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2733" daytime="08:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2734" daytime="08:48" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1065" daytime="08:56" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1066" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2616" />
                    <RANKING order="2" place="2" resultid="1817" />
                    <RANKING order="3" place="3" resultid="1857" />
                    <RANKING order="4" place="4" resultid="1623" />
                    <RANKING order="5" place="5" resultid="1510" />
                    <RANKING order="6" place="6" resultid="1862" />
                    <RANKING order="7" place="7" resultid="1807" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1505" />
                    <RANKING order="2" place="2" resultid="1708" />
                    <RANKING order="3" place="3" resultid="1673" />
                    <RANKING order="4" place="4" resultid="1693" />
                    <RANKING order="5" place="5" resultid="1743" />
                    <RANKING order="6" place="6" resultid="1417" />
                    <RANKING order="7" place="7" resultid="1453" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2735" daytime="08:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2736" daytime="09:02" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1068" daytime="09:10" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1069" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2500" />
                    <RANKING order="2" place="2" resultid="2042" />
                    <RANKING order="3" place="3" resultid="2067" />
                    <RANKING order="4" place="4" resultid="2509" />
                    <RANKING order="5" place="5" resultid="1633" />
                    <RANKING order="6" place="6" resultid="2082" />
                    <RANKING order="7" place="7" resultid="2087" />
                    <RANKING order="8" place="8" resultid="2022" />
                    <RANKING order="9" place="9" resultid="2137" />
                    <RANKING order="10" place="10" resultid="2077" />
                    <RANKING order="11" place="-1" resultid="2017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2541" />
                    <RANKING order="2" place="2" resultid="1892" />
                    <RANKING order="3" place="3" resultid="1638" />
                    <RANKING order="4" place="4" resultid="1520" />
                    <RANKING order="5" place="5" resultid="1957" />
                    <RANKING order="6" place="6" resultid="1992" />
                    <RANKING order="7" place="7" resultid="1977" />
                    <RANKING order="8" place="8" resultid="1379" />
                    <RANKING order="9" place="9" resultid="2697" />
                    <RANKING order="10" place="10" resultid="2641" />
                    <RANKING order="11" place="11" resultid="1241" />
                    <RANKING order="12" place="12" resultid="1932" />
                    <RANKING order="13" place="13" resultid="2514" />
                    <RANKING order="14" place="-1" resultid="1962" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2737" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2738" daytime="09:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2739" daytime="09:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2740" daytime="09:26" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1071" daytime="09:30" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1072" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2027" />
                    <RANKING order="2" place="2" resultid="2621" />
                    <RANKING order="3" place="3" resultid="1581" />
                    <RANKING order="4" place="4" resultid="2012" />
                    <RANKING order="5" place="5" resultid="2072" />
                    <RANKING order="6" place="6" resultid="2097" />
                    <RANKING order="7" place="7" resultid="2127" />
                    <RANKING order="8" place="8" resultid="2117" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1324" />
                    <RANKING order="2" place="2" resultid="1882" />
                    <RANKING order="3" place="3" resultid="1972" />
                    <RANKING order="4" place="4" resultid="1329" />
                    <RANKING order="5" place="5" resultid="2092" />
                    <RANKING order="6" place="6" resultid="2581" />
                    <RANKING order="7" place="7" resultid="2656" />
                    <RANKING order="8" place="8" resultid="2596" />
                    <RANKING order="9" place="9" resultid="1374" />
                    <RANKING order="10" place="10" resultid="2441" />
                    <RANKING order="11" place="11" resultid="2197" />
                    <RANKING order="12" place="-1" resultid="1902" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2741" daytime="09:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2742" daytime="09:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2743" daytime="09:40" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1074" daytime="09:46" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1075" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1359" />
                    <RANKING order="2" place="2" resultid="1758" />
                    <RANKING order="3" place="3" resultid="2157" />
                    <RANKING order="4" place="4" resultid="1587" />
                    <RANKING order="5" place="5" resultid="1261" />
                    <RANKING order="6" place="6" resultid="1768" />
                    <RANKING order="7" place="7" resultid="2386" />
                    <RANKING order="8" place="8" resultid="2352" />
                    <RANKING order="9" place="9" resultid="1917" />
                    <RANKING order="10" place="10" resultid="2303" />
                    <RANKING order="11" place="11" resultid="1987" />
                    <RANKING order="12" place="12" resultid="2631" />
                    <RANKING order="13" place="13" resultid="1567" />
                    <RANKING order="14" place="14" resultid="1787" />
                    <RANKING order="15" place="15" resultid="2488" />
                    <RANKING order="16" place="-1" resultid="1407" />
                    <RANKING order="17" place="-1" resultid="2702" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1076" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2322" />
                    <RANKING order="2" place="2" resultid="1713" />
                    <RANKING order="3" place="3" resultid="1723" />
                    <RANKING order="4" place="4" resultid="2307" />
                    <RANKING order="5" place="5" resultid="2142" />
                    <RANKING order="6" place="6" resultid="2536" />
                    <RANKING order="7" place="7" resultid="1309" />
                    <RANKING order="8" place="8" resultid="2667" />
                    <RANKING order="9" place="9" resultid="1877" />
                    <RANKING order="10" place="10" resultid="1576" />
                    <RANKING order="11" place="11" resultid="2343" />
                    <RANKING order="12" place="12" resultid="1427" />
                    <RANKING order="13" place="13" resultid="2522" />
                    <RANKING order="14" place="14" resultid="2678" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2744" daytime="09:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2745" daytime="09:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2746" daytime="09:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2747" daytime="09:52" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1077" daytime="09:54" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1078" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1624" />
                    <RANKING order="2" place="2" resultid="3375" />
                    <RANKING order="3" place="3" resultid="1511" />
                    <RANKING order="4" place="4" resultid="1458" />
                    <RANKING order="5" place="5" resultid="1339" />
                    <RANKING order="6" place="6" resultid="2601" />
                    <RANKING order="7" place="7" resultid="2611" />
                    <RANKING order="8" place="8" resultid="1852" />
                    <RANKING order="9" place="9" resultid="1837" />
                    <RANKING order="10" place="10" resultid="2673" />
                    <RANKING order="11" place="11" resultid="2428" />
                    <RANKING order="12" place="-1" resultid="1822" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1703" />
                    <RANKING order="2" place="2" resultid="2531" />
                    <RANKING order="3" place="3" resultid="1728" />
                    <RANKING order="4" place="4" resultid="1872" />
                    <RANKING order="5" place="5" resultid="2362" />
                    <RANKING order="6" place="6" resultid="1744" />
                    <RANKING order="7" place="7" resultid="1643" />
                    <RANKING order="8" place="8" resultid="1603" />
                    <RANKING order="9" place="9" resultid="1698" />
                    <RANKING order="10" place="10" resultid="2626" />
                    <RANKING order="11" place="11" resultid="1783" />
                    <RANKING order="12" place="12" resultid="1418" />
                    <RANKING order="13" place="13" resultid="1442" />
                    <RANKING order="14" place="-1" resultid="1847" />
                    <RANKING order="15" place="-1" resultid="1549" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2748" daytime="09:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2749" daytime="09:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2750" daytime="09:58" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2751" daytime="10:00" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1080" daytime="10:04" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1081" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2068" />
                    <RANKING order="2" place="2" resultid="2057" />
                    <RANKING order="3" place="3" resultid="1634" />
                    <RANKING order="4" place="4" resultid="1266" />
                    <RANKING order="5" place="5" resultid="2023" />
                    <RANKING order="6" place="6" resultid="2088" />
                    <RANKING order="7" place="7" resultid="2122" />
                    <RANKING order="8" place="8" resultid="1529" />
                    <RANKING order="9" place="9" resultid="2167" />
                    <RANKING order="10" place="10" resultid="2102" />
                    <RANKING order="11" place="11" resultid="2187" />
                    <RANKING order="12" place="12" resultid="2032" />
                    <RANKING order="13" place="13" resultid="1432" />
                    <RANKING order="14" place="14" resultid="2138" />
                    <RANKING order="15" place="15" resultid="2112" />
                    <RANKING order="16" place="-1" resultid="2018" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2542" />
                    <RANKING order="2" place="2" resultid="2332" />
                    <RANKING order="3" place="3" resultid="1893" />
                    <RANKING order="4" place="4" resultid="1628" />
                    <RANKING order="5" place="5" resultid="2002" />
                    <RANKING order="6" place="6" resultid="2698" />
                    <RANKING order="7" place="7" resultid="1571" />
                    <RANKING order="8" place="8" resultid="1251" />
                    <RANKING order="9" place="9" resultid="2357" />
                    <RANKING order="10" place="10" resultid="2007" />
                    <RANKING order="11" place="11" resultid="1521" />
                    <RANKING order="12" place="12" resultid="1319" />
                    <RANKING order="13" place="13" resultid="1993" />
                    <RANKING order="14" place="14" resultid="1481" />
                    <RANKING order="15" place="15" resultid="1897" />
                    <RANKING order="16" place="16" resultid="2688" />
                    <RANKING order="17" place="17" resultid="2438" />
                    <RANKING order="18" place="-1" resultid="2182" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2752" daytime="10:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2753" daytime="10:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2754" daytime="10:08" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2755" daytime="10:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2756" daytime="10:12" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1083" daytime="10:16" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1084" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2013" />
                    <RANKING order="2" place="2" resultid="2372" />
                    <RANKING order="3" place="3" resultid="2132" />
                    <RANKING order="4" place="4" resultid="2107" />
                    <RANKING order="5" place="5" resultid="1369" />
                    <RANKING order="6" place="6" resultid="1582" />
                    <RANKING order="7" place="7" resultid="2062" />
                    <RANKING order="8" place="8" resultid="2433" />
                    <RANKING order="9" place="9" resultid="2147" />
                    <RANKING order="10" place="10" resultid="2098" />
                    <RANKING order="11" place="11" resultid="2382" />
                    <RANKING order="12" place="12" resultid="2192" />
                    <RANKING order="13" place="13" resultid="2172" />
                    <RANKING order="14" place="14" resultid="1648" />
                    <RANKING order="15" place="15" resultid="2152" />
                    <RANKING order="16" place="16" resultid="2162" />
                    <RANKING order="17" place="17" resultid="2177" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1515" />
                    <RANKING order="2" place="2" resultid="1912" />
                    <RANKING order="3" place="3" resultid="2395" />
                    <RANKING order="4" place="4" resultid="2582" />
                    <RANKING order="5" place="5" resultid="2497" />
                    <RANKING order="6" place="6" resultid="1256" />
                    <RANKING order="7" place="7" resultid="1967" />
                    <RANKING order="8" place="8" resultid="1539" />
                    <RANKING order="9" place="9" resultid="1613" />
                    <RANKING order="10" place="10" resultid="1947" />
                    <RANKING order="11" place="11" resultid="1384" />
                    <RANKING order="12" place="12" resultid="2657" />
                    <RANKING order="13" place="13" resultid="1364" />
                    <RANKING order="14" place="14" resultid="1927" />
                    <RANKING order="15" place="15" resultid="1907" />
                    <RANKING order="16" place="16" resultid="2661" />
                    <RANKING order="17" place="17" resultid="1271" />
                    <RANKING order="18" place="18" resultid="1422" />
                    <RANKING order="19" place="19" resultid="1354" />
                    <RANKING order="20" place="20" resultid="1922" />
                    <RANKING order="21" place="21" resultid="2646" />
                    <RANKING order="22" place="22" resultid="2597" />
                    <RANKING order="23" place="23" resultid="2198" />
                    <RANKING order="24" place="24" resultid="2571" />
                    <RANKING order="25" place="25" resultid="1952" />
                    <RANKING order="26" place="25" resultid="2442" />
                    <RANKING order="27" place="27" resultid="1544" />
                    <RANKING order="28" place="-1" resultid="1942" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2757" daytime="10:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2758" daytime="10:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2759" daytime="10:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2760" daytime="10:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2761" daytime="10:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2762" daytime="10:26" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1086" daytime="10:28" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1087" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1753" />
                    <RANKING order="2" place="2" resultid="1802" />
                    <RANKING order="3" place="3" resultid="1797" />
                    <RANKING order="4" place="4" resultid="1812" />
                    <RANKING order="5" place="5" resultid="1448" />
                    <RANKING order="6" place="6" resultid="1887" />
                    <RANKING order="7" place="7" resultid="2347" />
                    <RANKING order="8" place="8" resultid="1412" />
                    <RANKING order="9" place="9" resultid="2302" />
                    <RANKING order="10" place="10" resultid="1279" />
                    <RANKING order="11" place="11" resultid="1289" />
                    <RANKING order="12" place="12" resultid="2420" />
                    <RANKING order="13" place="13" resultid="1566" />
                    <RANKING order="14" place="-1" resultid="2586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1833" />
                    <RANKING order="2" place="2" resultid="1774" />
                    <RANKING order="3" place="3" resultid="1982" />
                    <RANKING order="4" place="4" resultid="1764" />
                    <RANKING order="5" place="5" resultid="2561" />
                    <RANKING order="6" place="6" resultid="2666" />
                    <RANKING order="7" place="7" resultid="2415" />
                    <RANKING order="8" place="8" resultid="1247" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2763" daytime="10:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2764" daytime="10:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2765" daytime="10:36" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1089" daytime="10:40" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1090" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1236" />
                    <RANKING order="2" place="2" resultid="1608" />
                    <RANKING order="3" place="3" resultid="1748" />
                    <RANKING order="4" place="4" resultid="1997" />
                    <RANKING order="5" place="5" resultid="2551" />
                    <RANKING order="6" place="6" resultid="2591" />
                    <RANKING order="7" place="7" resultid="1792" />
                    <RANKING order="8" place="8" resultid="1344" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1299" />
                    <RANKING order="2" place="2" resultid="1663" />
                    <RANKING order="3" place="3" resultid="2483" />
                    <RANKING order="4" place="4" resultid="2327" />
                    <RANKING order="5" place="5" resultid="1668" />
                    <RANKING order="6" place="6" resultid="2317" />
                    <RANKING order="7" place="7" resultid="2556" />
                    <RANKING order="8" place="8" resultid="1284" />
                    <RANKING order="9" place="9" resultid="1304" />
                    <RANKING order="10" place="9" resultid="2651" />
                    <RANKING order="11" place="11" resultid="2400" />
                    <RANKING order="12" place="12" resultid="1437" />
                    <RANKING order="13" place="13" resultid="2683" />
                    <RANKING order="14" place="14" resultid="1334" />
                    <RANKING order="15" place="15" resultid="1827" />
                    <RANKING order="16" place="-1" resultid="1688" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2766" daytime="10:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2767" daytime="10:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2768" daytime="10:46" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1092" daytime="10:50" gender="X" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1093" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2242" />
                    <RANKING order="2" place="2" resultid="2266" />
                    <RANKING order="3" place="3" resultid="2290" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2769" daytime="10:50" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1094" daytime="10:56" gender="X" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1095" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2720" />
                    <RANKING order="2" place="2" resultid="2243" />
                    <RANKING order="3" place="3" resultid="1396" />
                    <RANKING order="4" place="4" resultid="1275" />
                    <RANKING order="5" place="5" resultid="1659" />
                    <RANKING order="6" place="6" resultid="2267" />
                    <RANKING order="7" place="7" resultid="2473" />
                    <RANKING order="8" place="8" resultid="2726" />
                    <RANKING order="9" place="9" resultid="2291" />
                    <RANKING order="10" place="10" resultid="1562" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2770" daytime="10:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2771" daytime="10:58" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1096" daytime="11:04" gender="X" number="13" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1097" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2240" />
                    <RANKING order="2" place="2" resultid="2288" />
                    <RANKING order="3" place="3" resultid="2718" />
                    <RANKING order="4" place="4" resultid="2264" />
                    <RANKING order="5" place="5" resultid="1394" />
                    <RANKING order="6" place="6" resultid="2724" />
                    <RANKING order="7" place="-1" resultid="2471" />
                    <RANKING order="8" place="-1" resultid="2730" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2772" daytime="11:04" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1098" daytime="11:08" gender="X" number="14" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1099" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2241" />
                    <RANKING order="2" place="2" resultid="2265" />
                    <RANKING order="3" place="3" resultid="2289" />
                    <RANKING order="4" place="4" resultid="1395" />
                    <RANKING order="5" place="5" resultid="2472" />
                    <RANKING order="6" place="6" resultid="2719" />
                    <RANKING order="7" place="7" resultid="2479" />
                    <RANKING order="8" place="8" resultid="2725" />
                    <RANKING order="9" place="-1" resultid="1496" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2773" daytime="11:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2774" daytime="11:12" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-05-24" daytime="15:40" endtime="18:33" number="2" officialmeeting="15:00" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1100" daytime="15:40" gender="F" number="15" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1101" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2354" />
                    <RANKING order="2" place="2" resultid="1799" />
                    <RANKING order="3" place="3" resultid="1759" />
                    <RANKING order="4" place="4" resultid="2379" />
                    <RANKING order="5" place="5" resultid="2369" />
                    <RANKING order="6" place="6" resultid="1939" />
                    <RANKING order="7" place="7" resultid="2608" />
                    <RANKING order="8" place="8" resultid="1316" />
                    <RANKING order="9" place="9" resultid="2314" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1835" />
                    <RANKING order="2" place="2" resultid="1725" />
                    <RANKING order="3" place="3" resultid="1685" />
                    <RANKING order="4" place="4" resultid="1739" />
                    <RANKING order="5" place="5" resultid="2340" />
                    <RANKING order="6" place="6" resultid="1404" />
                    <RANKING order="7" place="7" resultid="1465" />
                    <RANKING order="8" place="8" resultid="2411" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2775" daytime="15:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2776" daytime="15:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2777" daytime="15:46" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1103" daytime="15:50" gender="M" number="16" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1104" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1238" />
                    <RANKING order="2" place="2" resultid="1839" />
                    <RANKING order="3" place="3" resultid="1502" />
                    <RANKING order="4" place="4" resultid="1351" />
                    <RANKING order="5" place="5" resultid="3376" />
                    <RANKING order="6" place="6" resultid="1859" />
                    <RANKING order="7" place="-1" resultid="1750" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1665" />
                    <RANKING order="2" place="2" resultid="1508" />
                    <RANKING order="3" place="3" resultid="1734" />
                    <RANKING order="4" place="4" resultid="1874" />
                    <RANKING order="5" place="5" resultid="1455" />
                    <RANKING order="6" place="6" resultid="1605" />
                    <RANKING order="7" place="7" resultid="1644" />
                    <RANKING order="8" place="8" resultid="2628" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2778" daytime="15:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2779" daytime="15:52" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1106" daytime="15:56" gender="F" number="17" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1107" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2501" />
                    <RANKING order="2" place="2" resultid="2510" />
                    <RANKING order="3" place="3" resultid="2044" />
                    <RANKING order="4" place="4" resultid="2070" />
                    <RANKING order="5" place="5" resultid="1636" />
                    <RANKING order="6" place="6" resultid="2025" />
                    <RANKING order="7" place="7" resultid="2123" />
                    <RANKING order="8" place="8" resultid="2089" />
                    <RANKING order="9" place="9" resultid="2078" />
                    <RANKING order="10" place="10" resultid="2104" />
                    <RANKING order="11" place="-1" resultid="2019" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1108" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2333" />
                    <RANKING order="2" place="2" resultid="1895" />
                    <RANKING order="3" place="3" resultid="2636" />
                    <RANKING order="4" place="4" resultid="1380" />
                    <RANKING order="5" place="5" resultid="1959" />
                    <RANKING order="6" place="6" resultid="1979" />
                    <RANKING order="7" place="7" resultid="2047" />
                    <RANKING order="8" place="8" resultid="1630" />
                    <RANKING order="9" place="9" resultid="1899" />
                    <RANKING order="10" place="10" resultid="1252" />
                    <RANKING order="11" place="11" resultid="1573" />
                    <RANKING order="12" place="12" resultid="2689" />
                    <RANKING order="13" place="13" resultid="2519" />
                    <RANKING order="14" place="14" resultid="2008" />
                    <RANKING order="15" place="15" resultid="1933" />
                    <RANKING order="16" place="-1" resultid="1963" />
                    <RANKING order="17" place="-1" resultid="2183" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2780" daytime="15:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2781" daytime="15:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2782" daytime="16:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2783" daytime="16:04" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1109" daytime="16:06" gender="M" number="18" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1110" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2029" />
                    <RANKING order="2" place="2" resultid="1649" />
                    <RANKING order="3" place="3" resultid="2074" />
                    <RANKING order="4" place="4" resultid="1598" />
                    <RANKING order="5" place="5" resultid="2134" />
                    <RANKING order="6" place="6" resultid="2383" />
                    <RANKING order="7" place="7" resultid="2064" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1883" />
                    <RANKING order="2" place="2" resultid="1326" />
                    <RANKING order="3" place="3" resultid="1974" />
                    <RANKING order="4" place="4" resultid="1969" />
                    <RANKING order="5" place="5" resultid="1653" />
                    <RANKING order="6" place="6" resultid="1914" />
                    <RANKING order="7" place="7" resultid="1365" />
                    <RANKING order="8" place="8" resultid="1257" />
                    <RANKING order="9" place="9" resultid="2053" />
                    <RANKING order="10" place="10" resultid="2093" />
                    <RANKING order="11" place="11" resultid="1330" />
                    <RANKING order="12" place="12" resultid="2037" />
                    <RANKING order="13" place="13" resultid="1356" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2784" daytime="16:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2785" daytime="16:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2786" daytime="16:10" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1112" daytime="16:12" gender="F" number="19" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1113" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1114" daytime="16:12" gender="M" number="20" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1115" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1535" />
                    <RANKING order="2" place="2" resultid="2447" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2787" daytime="16:12" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1116" daytime="16:14" gender="F" number="21" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1117" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1804" />
                    <RANKING order="2" place="2" resultid="1755" />
                    <RANKING order="3" place="3" resultid="2388" />
                    <RANKING order="4" place="4" resultid="1869" />
                    <RANKING order="5" place="5" resultid="1814" />
                    <RANKING order="6" place="6" resultid="2349" />
                    <RANKING order="7" place="7" resultid="1415" />
                    <RANKING order="8" place="8" resultid="2304" />
                    <RANKING order="9" place="9" resultid="1556" />
                    <RANKING order="10" place="10" resultid="1262" />
                    <RANKING order="11" place="11" resultid="2490" />
                    <RANKING order="12" place="12" resultid="2422" />
                    <RANKING order="13" place="13" resultid="1569" />
                    <RANKING order="14" place="14" resultid="1788" />
                    <RANKING order="15" place="15" resultid="1409" />
                    <RANKING order="16" place="16" resultid="2704" />
                    <RANKING order="17" place="17" resultid="2632" />
                    <RANKING order="18" place="-1" resultid="2588" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1775" />
                    <RANKING order="2" place="2" resultid="1983" />
                    <RANKING order="3" place="3" resultid="2668" />
                    <RANKING order="4" place="4" resultid="1766" />
                    <RANKING order="5" place="5" resultid="2563" />
                    <RANKING order="6" place="6" resultid="2538" />
                    <RANKING order="7" place="7" resultid="1428" />
                    <RANKING order="8" place="8" resultid="1474" />
                    <RANKING order="9" place="9" resultid="2679" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2788" daytime="16:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2789" daytime="16:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2790" daytime="16:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2791" daytime="16:24" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1119" daytime="16:26" gender="M" number="22" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1120" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1610" />
                    <RANKING order="2" place="2" resultid="1844" />
                    <RANKING order="3" place="3" resultid="1999" />
                    <RANKING order="4" place="4" resultid="2553" />
                    <RANKING order="5" place="5" resultid="2593" />
                    <RANKING order="6" place="6" resultid="1860" />
                    <RANKING order="7" place="7" resultid="1794" />
                    <RANKING order="8" place="8" resultid="1864" />
                    <RANKING order="9" place="9" resultid="1492" />
                    <RANKING order="10" place="10" resultid="1346" />
                    <RANKING order="11" place="11" resultid="2613" />
                    <RANKING order="12" place="12" resultid="2494" />
                    <RANKING order="13" place="13" resultid="2578" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1301" />
                    <RANKING order="2" place="2" resultid="2485" />
                    <RANKING order="3" place="3" resultid="2329" />
                    <RANKING order="4" place="4" resultid="1666" />
                    <RANKING order="5" place="5" resultid="1296" />
                    <RANKING order="6" place="6" resultid="2319" />
                    <RANKING order="7" place="7" resultid="1710" />
                    <RANKING order="8" place="8" resultid="1745" />
                    <RANKING order="9" place="9" resultid="2653" />
                    <RANKING order="10" place="10" resultid="2558" />
                    <RANKING order="11" place="11" resultid="1306" />
                    <RANKING order="12" place="12" resultid="2402" />
                    <RANKING order="13" place="13" resultid="1286" />
                    <RANKING order="14" place="14" resultid="2459" />
                    <RANKING order="15" place="15" resultid="1699" />
                    <RANKING order="16" place="16" resultid="1595" />
                    <RANKING order="17" place="17" resultid="1439" />
                    <RANKING order="18" place="18" resultid="1784" />
                    <RANKING order="19" place="19" resultid="2685" />
                    <RANKING order="20" place="20" resultid="1551" />
                    <RANKING order="21" place="21" resultid="1336" />
                    <RANKING order="22" place="22" resultid="1829" />
                    <RANKING order="23" place="-1" resultid="1690" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2792" daytime="16:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2793" daytime="16:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2794" daytime="16:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2795" daytime="16:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2796" daytime="16:36" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1122" daytime="16:38" gender="F" number="23" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1123" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2503" />
                    <RANKING order="2" place="2" resultid="2084" />
                    <RANKING order="3" place="3" resultid="1434" />
                    <RANKING order="4" place="4" resultid="1268" />
                    <RANKING order="5" place="5" resultid="2060" />
                    <RANKING order="6" place="6" resultid="1531" />
                    <RANKING order="7" place="7" resultid="2125" />
                    <RANKING order="8" place="8" resultid="2140" />
                    <RANKING order="9" place="9" resultid="2080" />
                    <RANKING order="10" place="10" resultid="2114" />
                    <RANKING order="11" place="11" resultid="2189" />
                    <RANKING order="12" place="12" resultid="2034" />
                    <RANKING order="13" place="13" resultid="2169" />
                    <RANKING order="14" place="-1" resultid="2020" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1124" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2543" />
                    <RANKING order="2" place="2" resultid="1640" />
                    <RANKING order="3" place="3" resultid="2334" />
                    <RANKING order="4" place="4" resultid="2638" />
                    <RANKING order="5" place="5" resultid="1960" />
                    <RANKING order="6" place="6" resultid="1980" />
                    <RANKING order="7" place="7" resultid="1574" />
                    <RANKING order="8" place="8" resultid="1522" />
                    <RANKING order="9" place="9" resultid="2359" />
                    <RANKING order="10" place="10" resultid="1243" />
                    <RANKING order="11" place="11" resultid="1321" />
                    <RANKING order="12" place="12" resultid="2005" />
                    <RANKING order="13" place="13" resultid="2643" />
                    <RANKING order="14" place="14" resultid="2049" />
                    <RANKING order="15" place="15" resultid="1934" />
                    <RANKING order="16" place="16" resultid="2516" />
                    <RANKING order="17" place="17" resultid="2520" />
                    <RANKING order="18" place="18" resultid="1483" />
                    <RANKING order="19" place="-1" resultid="1965" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2797" daytime="16:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2798" daytime="16:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2799" daytime="16:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2800" daytime="16:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2801" daytime="16:50" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1125" daytime="16:54" gender="M" number="24" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1126" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2623" />
                    <RANKING order="2" place="2" resultid="2392" />
                    <RANKING order="3" place="3" resultid="2015" />
                    <RANKING order="4" place="4" resultid="1371" />
                    <RANKING order="5" place="5" resultid="2374" />
                    <RANKING order="6" place="6" resultid="2435" />
                    <RANKING order="7" place="7" resultid="2194" />
                    <RANKING order="8" place="8" resultid="2129" />
                    <RANKING order="9" place="9" resultid="2100" />
                    <RANKING order="10" place="10" resultid="2119" />
                    <RANKING order="11" place="11" resultid="2110" />
                    <RANKING order="12" place="12" resultid="2135" />
                    <RANKING order="13" place="13" resultid="2174" />
                    <RANKING order="14" place="14" resultid="2164" />
                    <RANKING order="15" place="15" resultid="2149" />
                    <RANKING order="16" place="16" resultid="2154" />
                    <RANKING order="17" place="17" resultid="2179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1884" />
                    <RANKING order="2" place="2" resultid="2454" />
                    <RANKING order="3" place="3" resultid="2095" />
                    <RANKING order="4" place="4" resultid="1517" />
                    <RANKING order="5" place="5" resultid="2583" />
                    <RANKING order="6" place="6" resultid="1615" />
                    <RANKING order="7" place="7" resultid="2055" />
                    <RANKING order="8" place="8" resultid="1273" />
                    <RANKING order="9" place="9" resultid="1909" />
                    <RANKING order="10" place="10" resultid="1915" />
                    <RANKING order="11" place="11" resultid="2598" />
                    <RANKING order="12" place="12" resultid="2397" />
                    <RANKING order="13" place="13" resultid="2573" />
                    <RANKING order="14" place="14" resultid="1655" />
                    <RANKING order="15" place="15" resultid="1386" />
                    <RANKING order="16" place="16" resultid="2658" />
                    <RANKING order="17" place="17" resultid="1376" />
                    <RANKING order="18" place="18" resultid="1949" />
                    <RANKING order="19" place="19" resultid="2648" />
                    <RANKING order="20" place="20" resultid="1424" />
                    <RANKING order="21" place="21" resultid="2039" />
                    <RANKING order="22" place="22" resultid="1970" />
                    <RANKING order="23" place="23" resultid="2443" />
                    <RANKING order="24" place="24" resultid="1929" />
                    <RANKING order="25" place="25" resultid="1541" />
                    <RANKING order="26" place="26" resultid="1924" />
                    <RANKING order="27" place="27" resultid="2663" />
                    <RANKING order="28" place="28" resultid="1546" />
                    <RANKING order="29" place="29" resultid="1526" />
                    <RANKING order="30" place="30" resultid="2199" />
                    <RANKING order="31" place="31" resultid="1954" />
                    <RANKING order="32" place="-1" resultid="1904" />
                    <RANKING order="33" place="-1" resultid="1944" />
                    <RANKING order="34" place="-1" resultid="2671" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2802" daytime="16:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2803" daytime="16:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2804" daytime="17:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2805" daytime="17:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2806" daytime="17:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2807" daytime="17:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2808" daytime="17:14" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1128" daytime="17:18" gender="F" number="25" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1129" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2210" />
                    <RANKING order="2" place="2" resultid="2221" />
                    <RANKING order="3" place="3" resultid="1477" />
                    <RANKING order="4" place="4" resultid="2217" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2809" daytime="17:18" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1130" daytime="17:20" gender="M" number="26" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1131" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1534" />
                    <RANKING order="2" place="2" resultid="1486" />
                    <RANKING order="3" place="3" resultid="2446" />
                    <RANKING order="4" place="4" resultid="2208" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2810" daytime="17:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1132" daytime="17:22" gender="F" number="27" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1133" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2568" />
                    <RANKING order="2" place="2" resultid="1360" />
                    <RANKING order="3" place="3" resultid="2158" />
                    <RANKING order="4" place="4" resultid="1450" />
                    <RANKING order="5" place="5" resultid="1769" />
                    <RANKING order="6" place="6" resultid="1803" />
                    <RANKING order="7" place="7" resultid="1589" />
                    <RANKING order="8" place="8" resultid="2547" />
                    <RANKING order="9" place="9" resultid="1813" />
                    <RANKING order="10" place="10" resultid="2348" />
                    <RANKING order="11" place="11" resultid="1889" />
                    <RANKING order="12" place="12" resultid="2607" />
                    <RANKING order="13" place="13" resultid="1281" />
                    <RANKING order="14" place="14" resultid="2387" />
                    <RANKING order="15" place="15" resultid="1568" />
                    <RANKING order="16" place="16" resultid="1918" />
                    <RANKING order="17" place="17" resultid="1315" />
                    <RANKING order="18" place="18" resultid="1291" />
                    <RANKING order="19" place="19" resultid="1988" />
                    <RANKING order="20" place="20" resultid="2489" />
                    <RANKING order="21" place="21" resultid="1555" />
                    <RANKING order="22" place="22" resultid="2421" />
                    <RANKING order="23" place="23" resultid="1408" />
                    <RANKING order="24" place="24" resultid="2703" />
                    <RANKING order="25" place="-1" resultid="2587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1134" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1680" />
                    <RANKING order="2" place="2" resultid="1720" />
                    <RANKING order="3" place="3" resultid="2562" />
                    <RANKING order="4" place="4" resultid="1765" />
                    <RANKING order="5" place="5" resultid="2339" />
                    <RANKING order="6" place="6" resultid="1403" />
                    <RANKING order="7" place="7" resultid="2417" />
                    <RANKING order="8" place="8" resultid="2308" />
                    <RANKING order="9" place="9" resultid="1310" />
                    <RANKING order="10" place="10" resultid="2525" />
                    <RANKING order="11" place="11" resultid="1249" />
                    <RANKING order="12" place="12" resultid="1878" />
                    <RANKING order="13" place="13" resultid="1473" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2811" daytime="17:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2812" daytime="17:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2813" daytime="17:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2814" daytime="17:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2815" daytime="17:32" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1135" daytime="17:36" gender="M" number="28" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1136" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1237" />
                    <RANKING order="2" place="2" resultid="1501" />
                    <RANKING order="3" place="3" resultid="1843" />
                    <RANKING order="4" place="4" resultid="2618" />
                    <RANKING order="5" place="5" resultid="1819" />
                    <RANKING order="6" place="6" resultid="1350" />
                    <RANKING order="7" place="7" resultid="2430" />
                    <RANKING order="8" place="8" resultid="2407" />
                    <RANKING order="9" place="9" resultid="1810" />
                    <RANKING order="10" place="10" resultid="2602" />
                    <RANKING order="11" place="11" resultid="2552" />
                    <RANKING order="12" place="12" resultid="1340" />
                    <RANKING order="13" place="13" resultid="2592" />
                    <RANKING order="14" place="14" resultid="2612" />
                    <RANKING order="15" place="15" resultid="1793" />
                    <RANKING order="16" place="16" resultid="1853" />
                    <RANKING order="17" place="17" resultid="1491" />
                    <RANKING order="18" place="18" resultid="2674" />
                    <RANKING order="19" place="19" resultid="2493" />
                    <RANKING order="20" place="20" resultid="2577" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1137" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1507" />
                    <RANKING order="2" place="2" resultid="1295" />
                    <RANKING order="3" place="3" resultid="1705" />
                    <RANKING order="4" place="4" resultid="2532" />
                    <RANKING order="5" place="5" resultid="1695" />
                    <RANKING order="6" place="6" resultid="1670" />
                    <RANKING order="7" place="6" resultid="1729" />
                    <RANKING order="8" place="8" resultid="1470" />
                    <RANKING order="9" place="9" resultid="1675" />
                    <RANKING order="10" place="10" resultid="2318" />
                    <RANKING order="11" place="11" resultid="1419" />
                    <RANKING order="12" place="12" resultid="1620" />
                    <RANKING order="13" place="13" resultid="2652" />
                    <RANKING order="14" place="14" resultid="1848" />
                    <RANKING order="15" place="15" resultid="2694" />
                    <RANKING order="16" place="16" resultid="1594" />
                    <RANKING order="17" place="17" resultid="1443" />
                    <RANKING order="18" place="18" resultid="2458" />
                    <RANKING order="19" place="19" resultid="1438" />
                    <RANKING order="20" place="20" resultid="2684" />
                    <RANKING order="21" place="21" resultid="1828" />
                    <RANKING order="22" place="-1" resultid="1550" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2816" daytime="17:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2817" daytime="17:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2818" daytime="17:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2819" daytime="17:44" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2820" daytime="17:46" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2821" daytime="17:48" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1138" daytime="17:52" gender="X" number="29" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1139" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2246" />
                    <RANKING order="2" place="2" resultid="2270" />
                    <RANKING order="3" place="3" resultid="2294" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2822" daytime="17:52" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1140" daytime="17:56" gender="X" number="30" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1141" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2245" />
                    <RANKING order="2" place="2" resultid="2728" />
                    <RANKING order="3" place="3" resultid="2269" />
                    <RANKING order="4" place="4" resultid="1398" />
                    <RANKING order="5" place="5" resultid="1660" />
                    <RANKING order="6" place="6" resultid="2475" />
                    <RANKING order="7" place="7" resultid="1276" />
                    <RANKING order="8" place="8" resultid="2293" />
                    <RANKING order="9" place="9" resultid="1563" />
                    <RANKING order="10" place="-1" resultid="2722" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2823" daytime="17:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2824" daytime="18:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1142" daytime="18:06" gender="X" number="31" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1143" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2271" />
                    <RANKING order="2" place="2" resultid="2247" />
                    <RANKING order="3" place="3" resultid="2295" />
                    <RANKING order="4" place="4" resultid="2723" />
                    <RANKING order="5" place="5" resultid="1399" />
                    <RANKING order="6" place="6" resultid="2476" />
                    <RANKING order="7" place="7" resultid="2729" />
                    <RANKING order="8" place="-1" resultid="2731" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2825" daytime="18:06" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1144" daytime="18:10" gender="X" number="32" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1145" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2244" />
                    <RANKING order="2" place="2" resultid="2268" />
                    <RANKING order="3" place="3" resultid="2292" />
                    <RANKING order="4" place="4" resultid="2474" />
                    <RANKING order="5" place="5" resultid="2721" />
                    <RANKING order="6" place="6" resultid="1397" />
                    <RANKING order="7" place="7" resultid="2480" />
                    <RANKING order="8" place="8" resultid="1497" />
                    <RANKING order="9" place="9" resultid="2727" />
                    <RANKING order="10" place="10" resultid="2528" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2826" daytime="18:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2827" daytime="18:14" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-05-25" daytime="08:40" endtime="11:35" number="3" officialmeeting="08:00" warmupfrom="07:30" warmupuntil="08:30">
          <EVENTS>
            <EVENT eventid="1146" daytime="08:40" gender="F" number="33" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1147" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2378" />
                    <RANKING order="2" place="2" resultid="2546" />
                    <RANKING order="3" place="3" resultid="1449" />
                    <RANKING order="4" place="4" resultid="1868" />
                    <RANKING order="5" place="5" resultid="1413" />
                    <RANKING order="6" place="6" resultid="2312" />
                    <RANKING order="7" place="7" resultid="1290" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1148" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1834" />
                    <RANKING order="2" place="2" resultid="1679" />
                    <RANKING order="3" place="3" resultid="1684" />
                    <RANKING order="4" place="4" resultid="2143" />
                    <RANKING order="5" place="5" resultid="2337" />
                    <RANKING order="6" place="6" resultid="1464" />
                    <RANKING order="7" place="7" resultid="2344" />
                    <RANKING order="8" place="8" resultid="1248" />
                    <RANKING order="9" place="9" resultid="2523" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2828" daytime="08:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2829" daytime="08:44" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1149" daytime="08:50" gender="M" number="34" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1150" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1838" />
                    <RANKING order="2" place="2" resultid="2617" />
                    <RANKING order="3" place="3" resultid="1818" />
                    <RANKING order="4" place="4" resultid="1512" />
                    <RANKING order="5" place="5" resultid="1609" />
                    <RANKING order="6" place="6" resultid="2405" />
                    <RANKING order="7" place="7" resultid="2429" />
                    <RANKING order="8" place="8" resultid="1808" />
                    <RANKING order="9" place="9" resultid="1863" />
                    <RANKING order="10" place="10" resultid="2492" />
                    <RANKING order="11" place="-1" resultid="1749" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1151" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1506" />
                    <RANKING order="2" place="2" resultid="1704" />
                    <RANKING order="3" place="3" resultid="1694" />
                    <RANKING order="4" place="4" resultid="1709" />
                    <RANKING order="5" place="5" resultid="1674" />
                    <RANKING order="6" place="6" resultid="1669" />
                    <RANKING order="7" place="7" resultid="1468" />
                    <RANKING order="8" place="8" resultid="1618" />
                    <RANKING order="9" place="9" resultid="2363" />
                    <RANKING order="10" place="10" resultid="1305" />
                    <RANKING order="11" place="11" resultid="2457" />
                    <RANKING order="12" place="12" resultid="2693" />
                    <RANKING order="13" place="13" resultid="2401" />
                    <RANKING order="14" place="-1" resultid="1689" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2830" daytime="08:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2831" daytime="08:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2832" daytime="08:58" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2833" daytime="09:04" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1152" daytime="09:08" gender="F" number="35" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1153" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2043" />
                    <RANKING order="2" place="2" resultid="2069" />
                    <RANKING order="3" place="3" resultid="1635" />
                    <RANKING order="4" place="4" resultid="2024" />
                    <RANKING order="5" place="5" resultid="2058" />
                    <RANKING order="6" place="6" resultid="2103" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1894" />
                    <RANKING order="2" place="2" resultid="1639" />
                    <RANKING order="3" place="3" resultid="1958" />
                    <RANKING order="4" place="4" resultid="1629" />
                    <RANKING order="5" place="5" resultid="1994" />
                    <RANKING order="6" place="6" resultid="2003" />
                    <RANKING order="7" place="7" resultid="1898" />
                    <RANKING order="8" place="8" resultid="1978" />
                    <RANKING order="9" place="9" resultid="1572" />
                    <RANKING order="10" place="10" resultid="1320" />
                    <RANKING order="11" place="11" resultid="2505" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2834" daytime="09:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2835" daytime="09:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2836" daytime="09:20" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1155" daytime="09:26" gender="M" number="36" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1156" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2028" />
                    <RANKING order="2" place="2" resultid="2622" />
                    <RANKING order="3" place="3" resultid="2014" />
                    <RANKING order="4" place="4" resultid="1370" />
                    <RANKING order="5" place="5" resultid="2073" />
                    <RANKING order="6" place="6" resultid="2063" />
                    <RANKING order="7" place="7" resultid="2108" />
                    <RANKING order="8" place="8" resultid="2133" />
                    <RANKING order="9" place="9" resultid="2128" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1325" />
                    <RANKING order="2" place="2" resultid="1973" />
                    <RANKING order="3" place="3" resultid="1913" />
                    <RANKING order="4" place="4" resultid="1516" />
                    <RANKING order="5" place="5" resultid="1968" />
                    <RANKING order="6" place="6" resultid="1385" />
                    <RANKING order="7" place="7" resultid="2052" />
                    <RANKING order="8" place="8" resultid="2647" />
                    <RANKING order="9" place="9" resultid="1355" />
                    <RANKING order="10" place="-1" resultid="1903" />
                    <RANKING order="11" place="-1" resultid="1943" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2837" daytime="09:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2838" daytime="09:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2839" daytime="09:36" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1158" daytime="09:42" gender="F" number="37" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1159" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2567" />
                    <RANKING order="2" place="2" resultid="2353" />
                    <RANKING order="3" place="3" resultid="2368" />
                    <RANKING order="4" place="4" resultid="1754" />
                    <RANKING order="5" place="5" resultid="1798" />
                    <RANKING order="6" place="6" resultid="1588" />
                    <RANKING order="7" place="7" resultid="2425" />
                    <RANKING order="8" place="8" resultid="1938" />
                    <RANKING order="9" place="9" resultid="1280" />
                    <RANKING order="10" place="10" resultid="1414" />
                    <RANKING order="11" place="11" resultid="2606" />
                    <RANKING order="12" place="12" resultid="2313" />
                    <RANKING order="13" place="13" resultid="1888" />
                    <RANKING order="14" place="14" resultid="1314" />
                    <RANKING order="15" place="15" resultid="1554" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1160" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1724" />
                    <RANKING order="2" place="2" resultid="2323" />
                    <RANKING order="3" place="3" resultid="1719" />
                    <RANKING order="4" place="4" resultid="2338" />
                    <RANKING order="5" place="5" resultid="2416" />
                    <RANKING order="6" place="6" resultid="1402" />
                    <RANKING order="7" place="7" resultid="1577" />
                    <RANKING order="8" place="8" resultid="2537" />
                    <RANKING order="9" place="9" resultid="2410" />
                    <RANKING order="10" place="10" resultid="2524" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2840" daytime="09:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2841" daytime="09:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2842" daytime="09:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2843" daytime="09:48" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1161" daytime="09:50" gender="M" number="38" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1162" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1500" />
                    <RANKING order="2" place="2" resultid="1459" />
                    <RANKING order="3" place="3" resultid="1842" />
                    <RANKING order="4" place="4" resultid="1823" />
                    <RANKING order="5" place="5" resultid="1349" />
                    <RANKING order="6" place="6" resultid="3377" />
                    <RANKING order="7" place="7" resultid="1998" />
                    <RANKING order="8" place="8" resultid="1858" />
                    <RANKING order="9" place="9" resultid="2406" />
                    <RANKING order="10" place="10" resultid="1809" />
                    <RANKING order="11" place="11" resultid="1345" />
                    <RANKING order="12" place="12" resultid="2576" />
                    <RANKING order="13" place="-1" resultid="1490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1163" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1664" />
                    <RANKING order="2" place="2" resultid="1300" />
                    <RANKING order="3" place="3" resultid="1294" />
                    <RANKING order="4" place="4" resultid="1733" />
                    <RANKING order="5" place="5" resultid="1454" />
                    <RANKING order="6" place="6" resultid="2328" />
                    <RANKING order="7" place="7" resultid="1873" />
                    <RANKING order="8" place="8" resultid="2557" />
                    <RANKING order="9" place="9" resultid="1469" />
                    <RANKING order="10" place="10" resultid="1619" />
                    <RANKING order="11" place="11" resultid="1604" />
                    <RANKING order="12" place="12" resultid="1285" />
                    <RANKING order="13" place="13" resultid="2627" />
                    <RANKING order="14" place="14" resultid="1335" />
                    <RANKING order="15" place="15" resultid="1593" />
                    <RANKING order="16" place="-1" resultid="2484" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2844" daytime="09:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2845" daytime="09:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2846" daytime="09:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2847" daytime="09:56" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1164" daytime="09:58" gender="F" number="39" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1165" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2502" />
                    <RANKING order="2" place="2" resultid="2511" />
                    <RANKING order="3" place="3" resultid="2083" />
                    <RANKING order="4" place="4" resultid="1530" />
                    <RANKING order="5" place="5" resultid="1267" />
                    <RANKING order="6" place="6" resultid="2124" />
                    <RANKING order="7" place="7" resultid="2105" />
                    <RANKING order="8" place="8" resultid="2113" />
                    <RANKING order="9" place="9" resultid="1433" />
                    <RANKING order="10" place="10" resultid="2168" />
                    <RANKING order="11" place="11" resultid="2079" />
                    <RANKING order="12" place="12" resultid="2033" />
                    <RANKING order="13" place="13" resultid="2059" />
                    <RANKING order="14" place="14" resultid="2188" />
                    <RANKING order="15" place="15" resultid="2139" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1381" />
                    <RANKING order="2" place="2" resultid="2637" />
                    <RANKING order="3" place="3" resultid="2699" />
                    <RANKING order="4" place="4" resultid="2048" />
                    <RANKING order="5" place="5" resultid="2642" />
                    <RANKING order="6" place="6" resultid="1242" />
                    <RANKING order="7" place="7" resultid="1631" />
                    <RANKING order="8" place="8" resultid="1253" />
                    <RANKING order="9" place="9" resultid="2358" />
                    <RANKING order="10" place="10" resultid="2009" />
                    <RANKING order="11" place="11" resultid="1900" />
                    <RANKING order="12" place="12" resultid="2004" />
                    <RANKING order="13" place="13" resultid="2450" />
                    <RANKING order="14" place="14" resultid="2515" />
                    <RANKING order="15" place="15" resultid="1482" />
                    <RANKING order="16" place="16" resultid="2690" />
                    <RANKING order="17" place="17" resultid="2506" />
                    <RANKING order="18" place="-1" resultid="1964" />
                    <RANKING order="19" place="-1" resultid="2184" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2848" daytime="09:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2849" daytime="10:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2850" daytime="10:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2851" daytime="10:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2852" daytime="10:10" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1167" daytime="10:12" gender="M" number="40" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1168" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2030" />
                    <RANKING order="2" place="2" resultid="1650" />
                    <RANKING order="3" place="3" resultid="2373" />
                    <RANKING order="4" place="4" resultid="1599" />
                    <RANKING order="5" place="5" resultid="2193" />
                    <RANKING order="6" place="6" resultid="1583" />
                    <RANKING order="7" place="7" resultid="2075" />
                    <RANKING order="8" place="8" resultid="2065" />
                    <RANKING order="9" place="9" resultid="2434" />
                    <RANKING order="10" place="10" resultid="2148" />
                    <RANKING order="11" place="11" resultid="2109" />
                    <RANKING order="12" place="12" resultid="2178" />
                    <RANKING order="13" place="13" resultid="2099" />
                    <RANKING order="14" place="14" resultid="2118" />
                    <RANKING order="15" place="15" resultid="2173" />
                    <RANKING order="16" place="16" resultid="2163" />
                    <RANKING order="17" place="17" resultid="2153" />
                    <RANKING order="18" place="-1" resultid="2391" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1258" />
                    <RANKING order="2" place="2" resultid="2094" />
                    <RANKING order="3" place="3" resultid="2453" />
                    <RANKING order="4" place="4" resultid="1614" />
                    <RANKING order="5" place="5" resultid="1948" />
                    <RANKING order="6" place="6" resultid="2054" />
                    <RANKING order="7" place="7" resultid="1272" />
                    <RANKING order="8" place="8" resultid="1654" />
                    <RANKING order="9" place="9" resultid="1423" />
                    <RANKING order="10" place="10" resultid="2572" />
                    <RANKING order="11" place="11" resultid="2396" />
                    <RANKING order="12" place="12" resultid="2038" />
                    <RANKING order="13" place="13" resultid="1375" />
                    <RANKING order="14" place="14" resultid="2662" />
                    <RANKING order="15" place="15" resultid="1331" />
                    <RANKING order="16" place="16" resultid="1923" />
                    <RANKING order="17" place="17" resultid="1928" />
                    <RANKING order="18" place="18" resultid="1540" />
                    <RANKING order="19" place="19" resultid="1953" />
                    <RANKING order="20" place="20" resultid="1525" />
                    <RANKING order="21" place="21" resultid="1545" />
                    <RANKING order="22" place="-1" resultid="1366" />
                    <RANKING order="23" place="-1" resultid="1908" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2853" daytime="10:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2854" daytime="10:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2855" daytime="10:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2856" daytime="10:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2857" daytime="10:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2858" daytime="10:26" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1170" daytime="10:30" gender="F" number="41" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1171" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1361" />
                    <RANKING order="2" place="2" resultid="1760" />
                    <RANKING order="3" place="3" resultid="1263" />
                    <RANKING order="4" place="4" resultid="2159" />
                    <RANKING order="5" place="5" resultid="1590" />
                    <RANKING order="6" place="6" resultid="1770" />
                    <RANKING order="7" place="7" resultid="1989" />
                    <RANKING order="8" place="8" resultid="1919" />
                    <RANKING order="9" place="9" resultid="2633" />
                    <RANKING order="10" place="10" resultid="1789" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2324" />
                    <RANKING order="2" place="2" resultid="1714" />
                    <RANKING order="3" place="3" resultid="1740" />
                    <RANKING order="4" place="4" resultid="1984" />
                    <RANKING order="5" place="5" resultid="2144" />
                    <RANKING order="6" place="6" resultid="2309" />
                    <RANKING order="7" place="7" resultid="1311" />
                    <RANKING order="8" place="8" resultid="1879" />
                    <RANKING order="9" place="9" resultid="2345" />
                    <RANKING order="10" place="10" resultid="1429" />
                    <RANKING order="11" place="11" resultid="2680" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2859" daytime="10:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2860" daytime="10:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2861" daytime="10:36" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3396" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1173" daytime="10:38" gender="M" number="42" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1174" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1625" />
                    <RANKING order="2" place="2" resultid="1513" />
                    <RANKING order="3" place="3" resultid="2603" />
                    <RANKING order="4" place="4" resultid="1341" />
                    <RANKING order="5" place="5" resultid="1854" />
                    <RANKING order="6" place="6" resultid="2675" />
                    <RANKING order="7" place="-1" resultid="1824" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1706" />
                    <RANKING order="2" place="2" resultid="2533" />
                    <RANKING order="3" place="3" resultid="1730" />
                    <RANKING order="4" place="4" resultid="1875" />
                    <RANKING order="5" place="5" resultid="2364" />
                    <RANKING order="6" place="6" resultid="1746" />
                    <RANKING order="7" place="7" resultid="1645" />
                    <RANKING order="8" place="8" resultid="1700" />
                    <RANKING order="9" place="9" resultid="2629" />
                    <RANKING order="10" place="10" resultid="1785" />
                    <RANKING order="11" place="-1" resultid="1849" />
                    <RANKING order="12" place="-1" resultid="1444" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2862" daytime="10:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2863" daytime="10:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2864" daytime="10:46" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1176" daytime="10:48" gender="F" number="43" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1177" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2226" />
                    <RANKING order="2" place="2" resultid="2250" />
                    <RANKING order="3" place="3" resultid="2274" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2865" daytime="10:48" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1178" daytime="10:54" gender="F" number="44" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1179" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2706" />
                    <RANKING order="2" place="2" resultid="2224" />
                    <RANKING order="3" place="3" resultid="2461" />
                    <RANKING order="4" place="4" resultid="2526" />
                    <RANKING order="5" place="-1" resultid="2248" />
                    <RANKING order="6" place="-1" resultid="2272" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2866" daytime="10:54" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1180" daytime="10:58" gender="M" number="45" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1181" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2234" />
                    <RANKING order="2" place="2" resultid="2467" />
                    <RANKING order="3" place="3" resultid="2258" />
                    <RANKING order="4" place="4" resultid="2282" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2867" daytime="10:58" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1182" daytime="11:02" gender="M" number="46" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1183" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2232" />
                    <RANKING order="2" place="2" resultid="1390" />
                    <RANKING order="3" place="3" resultid="2712" />
                    <RANKING order="4" place="4" resultid="2256" />
                    <RANKING order="5" place="5" resultid="1558" />
                    <RANKING order="6" place="6" resultid="2280" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2868" daytime="11:02" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1184" daytime="11:08" gender="F" number="47" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1185" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2225" />
                    <RANKING order="2" place="2" resultid="2249" />
                    <RANKING order="3" place="3" resultid="2462" />
                    <RANKING order="4" place="4" resultid="1388" />
                    <RANKING order="5" place="5" resultid="2707" />
                    <RANKING order="6" place="6" resultid="2273" />
                    <RANKING order="7" place="-1" resultid="2477" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2869" daytime="11:08" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1186" daytime="11:12" gender="F" number="48" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1187" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2227" />
                    <RANKING order="2" place="2" resultid="2251" />
                    <RANKING order="3" place="3" resultid="2463" />
                    <RANKING order="4" place="4" resultid="2275" />
                    <RANKING order="5" place="5" resultid="2708" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2870" daytime="11:12" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1188" daytime="11:16" gender="M" number="49" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1189" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2233" />
                    <RANKING order="2" place="2" resultid="2257" />
                    <RANKING order="3" place="3" resultid="2713" />
                    <RANKING order="4" place="4" resultid="2281" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2871" daytime="11:16" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1190" daytime="11:20" gender="M" number="50" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1191" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2235" />
                    <RANKING order="2" place="2" resultid="2259" />
                    <RANKING order="3" place="3" resultid="1391" />
                    <RANKING order="4" place="4" resultid="2283" />
                    <RANKING order="5" place="5" resultid="2468" />
                    <RANKING order="6" place="6" resultid="1559" />
                    <RANKING order="7" place="7" resultid="1494" />
                    <RANKING order="8" place="8" resultid="2714" />
                    <RANKING order="9" place="9" resultid="1657" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2872" daytime="11:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2873" daytime="11:24" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-05-25" daytime="15:40" endtime="18:18" number="4" officialmeeting="15:00" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1192" daytime="15:40" gender="F" number="51" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1193" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2569" />
                    <RANKING order="2" place="2" resultid="2380" />
                    <RANKING order="3" place="3" resultid="1761" />
                    <RANKING order="4" place="4" resultid="2355" />
                    <RANKING order="5" place="5" resultid="1800" />
                    <RANKING order="6" place="6" resultid="2548" />
                    <RANKING order="7" place="7" resultid="2370" />
                    <RANKING order="8" place="8" resultid="1890" />
                    <RANKING order="9" place="9" resultid="1282" />
                    <RANKING order="10" place="10" resultid="1940" />
                    <RANKING order="11" place="11" resultid="1292" />
                    <RANKING order="12" place="12" resultid="1317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1686" />
                    <RANKING order="2" place="2" resultid="1726" />
                    <RANKING order="3" place="3" resultid="1721" />
                    <RANKING order="4" place="4" resultid="1741" />
                    <RANKING order="5" place="5" resultid="1715" />
                    <RANKING order="6" place="6" resultid="2564" />
                    <RANKING order="7" place="7" resultid="2325" />
                    <RANKING order="8" place="8" resultid="2418" />
                    <RANKING order="9" place="9" resultid="1578" />
                    <RANKING order="10" place="10" resultid="2298" />
                    <RANKING order="11" place="-1" resultid="2412" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2874" daytime="15:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2875" daytime="15:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2876" daytime="15:50" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1195" daytime="15:56" gender="M" number="52" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1196" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1626" />
                    <RANKING order="2" place="2" resultid="1840" />
                    <RANKING order="3" place="3" resultid="1825" />
                    <RANKING order="4" place="4" resultid="1611" />
                    <RANKING order="5" place="5" resultid="2619" />
                    <RANKING order="6" place="6" resultid="1820" />
                    <RANKING order="7" place="7" resultid="2408" />
                    <RANKING order="8" place="8" resultid="1855" />
                    <RANKING order="9" place="9" resultid="1795" />
                    <RANKING order="10" place="-1" resultid="1461" />
                    <RANKING order="11" place="-1" resultid="2000" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1197" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1731" />
                    <RANKING order="2" place="2" resultid="1736" />
                    <RANKING order="3" place="3" resultid="2365" />
                    <RANKING order="4" place="4" resultid="2486" />
                    <RANKING order="5" place="5" resultid="1606" />
                    <RANKING order="6" place="6" resultid="1621" />
                    <RANKING order="7" place="7" resultid="1646" />
                    <RANKING order="8" place="8" resultid="1701" />
                    <RANKING order="9" place="-1" resultid="2330" />
                    <RANKING order="10" place="-1" resultid="1691" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2877" daytime="15:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2878" daytime="16:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2879" daytime="16:06" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1198" daytime="16:10" gender="F" number="53" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1199" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2212" />
                    <RANKING order="2" place="2" resultid="2223" />
                    <RANKING order="3" place="3" resultid="1479" />
                    <RANKING order="4" place="4" resultid="2206" />
                    <RANKING order="5" place="5" resultid="2219" />
                    <RANKING order="6" place="6" resultid="2215" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2880" daytime="16:10" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1200" daytime="16:14" gender="M" number="54" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1201" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1488" />
                    <RANKING order="2" place="2" resultid="1537" />
                    <RANKING order="3" place="3" resultid="2203" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2881" daytime="16:14" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1202" daytime="16:16" gender="F" number="55" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1203" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2090" />
                    <RANKING order="2" place="2" resultid="2045" />
                    <RANKING order="3" place="3" resultid="2085" />
                    <RANKING order="4" place="4" resultid="2512" />
                    <RANKING order="5" place="5" resultid="1269" />
                    <RANKING order="6" place="6" resultid="1532" />
                    <RANKING order="7" place="7" resultid="1435" />
                    <RANKING order="8" place="8" resultid="2115" />
                    <RANKING order="9" place="9" resultid="2190" />
                    <RANKING order="10" place="10" resultid="2170" />
                    <RANKING order="11" place="11" resultid="2035" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1204" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2544" />
                    <RANKING order="2" place="2" resultid="2335" />
                    <RANKING order="3" place="3" resultid="2639" />
                    <RANKING order="4" place="4" resultid="1641" />
                    <RANKING order="5" place="5" resultid="2360" />
                    <RANKING order="6" place="6" resultid="1523" />
                    <RANKING order="7" place="7" resultid="1244" />
                    <RANKING order="8" place="8" resultid="1254" />
                    <RANKING order="9" place="9" resultid="2700" />
                    <RANKING order="10" place="10" resultid="2050" />
                    <RANKING order="11" place="11" resultid="2644" />
                    <RANKING order="12" place="12" resultid="2010" />
                    <RANKING order="13" place="13" resultid="1382" />
                    <RANKING order="14" place="14" resultid="1995" />
                    <RANKING order="15" place="15" resultid="1935" />
                    <RANKING order="16" place="16" resultid="1322" />
                    <RANKING order="17" place="17" resultid="2507" />
                    <RANKING order="18" place="18" resultid="2517" />
                    <RANKING order="19" place="19" resultid="2451" />
                    <RANKING order="20" place="20" resultid="2439" />
                    <RANKING order="21" place="21" resultid="1484" />
                    <RANKING order="22" place="22" resultid="2691" />
                    <RANKING order="23" place="23" resultid="2185" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2882" daytime="16:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2883" daytime="16:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2884" daytime="16:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2885" daytime="16:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2886" daytime="16:24" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1205" daytime="16:26" gender="M" number="56" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1206" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2624" />
                    <RANKING order="2" place="2" resultid="1651" />
                    <RANKING order="3" place="3" resultid="1600" />
                    <RANKING order="4" place="4" resultid="2375" />
                    <RANKING order="5" place="5" resultid="1584" />
                    <RANKING order="6" place="6" resultid="2393" />
                    <RANKING order="7" place="7" resultid="1372" />
                    <RANKING order="8" place="8" resultid="2195" />
                    <RANKING order="9" place="9" resultid="2436" />
                    <RANKING order="10" place="10" resultid="2384" />
                    <RANKING order="11" place="11" resultid="2130" />
                    <RANKING order="12" place="12" resultid="2120" />
                    <RANKING order="13" place="13" resultid="2165" />
                    <RANKING order="14" place="14" resultid="2150" />
                    <RANKING order="15" place="15" resultid="2175" />
                    <RANKING order="16" place="16" resultid="2155" />
                    <RANKING order="17" place="17" resultid="2180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1327" />
                    <RANKING order="2" place="2" resultid="1885" />
                    <RANKING order="3" place="3" resultid="1518" />
                    <RANKING order="4" place="4" resultid="1975" />
                    <RANKING order="5" place="5" resultid="1367" />
                    <RANKING order="6" place="6" resultid="2455" />
                    <RANKING order="7" place="7" resultid="1259" />
                    <RANKING order="8" place="8" resultid="2584" />
                    <RANKING order="9" place="9" resultid="1274" />
                    <RANKING order="10" place="10" resultid="2040" />
                    <RANKING order="11" place="11" resultid="2599" />
                    <RANKING order="12" place="12" resultid="2398" />
                    <RANKING order="13" place="13" resultid="1616" />
                    <RANKING order="14" place="14" resultid="1332" />
                    <RANKING order="15" place="15" resultid="1656" />
                    <RANKING order="16" place="16" resultid="2498" />
                    <RANKING order="17" place="17" resultid="1387" />
                    <RANKING order="18" place="18" resultid="2659" />
                    <RANKING order="19" place="19" resultid="1425" />
                    <RANKING order="20" place="20" resultid="2574" />
                    <RANKING order="21" place="21" resultid="1950" />
                    <RANKING order="22" place="22" resultid="1377" />
                    <RANKING order="23" place="23" resultid="2649" />
                    <RANKING order="24" place="24" resultid="2444" />
                    <RANKING order="25" place="25" resultid="1930" />
                    <RANKING order="26" place="26" resultid="1542" />
                    <RANKING order="27" place="27" resultid="2664" />
                    <RANKING order="28" place="28" resultid="1357" />
                    <RANKING order="29" place="29" resultid="1925" />
                    <RANKING order="30" place="30" resultid="1527" />
                    <RANKING order="31" place="31" resultid="2200" />
                    <RANKING order="32" place="32" resultid="1547" />
                    <RANKING order="33" place="33" resultid="1955" />
                    <RANKING order="34" place="-1" resultid="1905" />
                    <RANKING order="35" place="-1" resultid="1910" />
                    <RANKING order="36" place="-1" resultid="1945" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2887" daytime="16:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2888" daytime="16:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2889" daytime="16:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2890" daytime="16:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2891" daytime="16:36" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2892" daytime="16:38" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2893" daytime="16:40" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1208" daytime="16:42" gender="F" number="57" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1209" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1362" />
                    <RANKING order="2" place="2" resultid="2160" />
                    <RANKING order="3" place="3" resultid="1805" />
                    <RANKING order="4" place="4" resultid="1870" />
                    <RANKING order="5" place="5" resultid="1451" />
                    <RANKING order="6" place="6" resultid="1591" />
                    <RANKING order="7" place="7" resultid="1756" />
                    <RANKING order="8" place="8" resultid="1771" />
                    <RANKING order="9" place="9" resultid="2350" />
                    <RANKING order="10" place="10" resultid="2389" />
                    <RANKING order="11" place="11" resultid="1815" />
                    <RANKING order="12" place="12" resultid="2426" />
                    <RANKING order="13" place="13" resultid="2549" />
                    <RANKING order="14" place="14" resultid="1557" />
                    <RANKING order="15" place="15" resultid="1920" />
                    <RANKING order="16" place="16" resultid="1264" />
                    <RANKING order="17" place="17" resultid="2609" />
                    <RANKING order="18" place="18" resultid="2305" />
                    <RANKING order="19" place="19" resultid="2315" />
                    <RANKING order="20" place="20" resultid="1410" />
                    <RANKING order="21" place="21" resultid="1990" />
                    <RANKING order="22" place="22" resultid="2423" />
                    <RANKING order="23" place="23" resultid="1790" />
                    <RANKING order="24" place="24" resultid="2705" />
                    <RANKING order="25" place="25" resultid="2634" />
                    <RANKING order="26" place="-1" resultid="2589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1210" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1776" />
                    <RANKING order="2" place="2" resultid="1681" />
                    <RANKING order="3" place="3" resultid="2145" />
                    <RANKING order="4" place="4" resultid="1985" />
                    <RANKING order="5" place="5" resultid="2539" />
                    <RANKING order="6" place="6" resultid="2669" />
                    <RANKING order="7" place="7" resultid="1716" />
                    <RANKING order="8" place="8" resultid="1312" />
                    <RANKING order="9" place="9" resultid="1466" />
                    <RANKING order="10" place="10" resultid="2310" />
                    <RANKING order="11" place="11" resultid="1579" />
                    <RANKING order="12" place="12" resultid="2299" />
                    <RANKING order="13" place="13" resultid="2413" />
                    <RANKING order="14" place="14" resultid="1880" />
                    <RANKING order="15" place="15" resultid="1430" />
                    <RANKING order="16" place="16" resultid="2681" />
                    <RANKING order="17" place="17" resultid="1475" />
                    <RANKING order="18" place="-1" resultid="1405" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2894" daytime="16:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2895" daytime="16:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2896" daytime="16:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2897" daytime="16:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2898" daytime="16:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2899" daytime="16:52" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1211" daytime="16:54" gender="M" number="58" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1212" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1239" />
                    <RANKING order="2" place="2" resultid="1503" />
                    <RANKING order="3" place="3" resultid="1460" />
                    <RANKING order="4" place="4" resultid="1845" />
                    <RANKING order="5" place="5" resultid="2554" />
                    <RANKING order="6" place="6" resultid="1352" />
                    <RANKING order="7" place="7" resultid="2604" />
                    <RANKING order="8" place="8" resultid="1751" />
                    <RANKING order="9" place="9" resultid="1342" />
                    <RANKING order="10" place="10" resultid="3378" />
                    <RANKING order="11" place="11" resultid="2431" />
                    <RANKING order="12" place="12" resultid="2594" />
                    <RANKING order="13" place="13" resultid="1865" />
                    <RANKING order="14" place="14" resultid="1347" />
                    <RANKING order="15" place="15" resultid="1493" />
                    <RANKING order="16" place="16" resultid="2614" />
                    <RANKING order="17" place="17" resultid="2676" />
                    <RANKING order="18" place="18" resultid="2579" />
                    <RANKING order="19" place="19" resultid="2495" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1213" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1297" />
                    <RANKING order="2" place="2" resultid="1302" />
                    <RANKING order="3" place="3" resultid="1471" />
                    <RANKING order="4" place="4" resultid="2534" />
                    <RANKING order="5" place="5" resultid="1696" />
                    <RANKING order="6" place="6" resultid="2320" />
                    <RANKING order="7" place="7" resultid="1671" />
                    <RANKING order="8" place="8" resultid="1676" />
                    <RANKING order="9" place="8" resultid="1711" />
                    <RANKING order="10" place="10" resultid="1735" />
                    <RANKING order="11" place="11" resultid="1287" />
                    <RANKING order="12" place="12" resultid="1456" />
                    <RANKING order="13" place="13" resultid="1850" />
                    <RANKING order="14" place="14" resultid="1420" />
                    <RANKING order="15" place="15" resultid="2559" />
                    <RANKING order="16" place="16" resultid="1307" />
                    <RANKING order="17" place="17" resultid="2695" />
                    <RANKING order="18" place="18" resultid="2460" />
                    <RANKING order="19" place="19" resultid="2654" />
                    <RANKING order="20" place="20" resultid="1596" />
                    <RANKING order="21" place="21" resultid="1440" />
                    <RANKING order="22" place="22" resultid="2403" />
                    <RANKING order="23" place="23" resultid="1445" />
                    <RANKING order="24" place="24" resultid="1337" />
                    <RANKING order="25" place="25" resultid="1552" />
                    <RANKING order="26" place="26" resultid="2686" />
                    <RANKING order="27" place="27" resultid="1830" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2900" daytime="16:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2901" daytime="16:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2902" daytime="16:58" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2903" daytime="17:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2904" daytime="17:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2905" daytime="17:02" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1214" daytime="17:04" gender="F" number="59" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1215" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2211" />
                    <RANKING order="2" place="2" resultid="2222" />
                    <RANKING order="3" place="3" resultid="1478" />
                    <RANKING order="4" place="4" resultid="2218" />
                    <RANKING order="5" place="5" resultid="2205" />
                    <RANKING order="6" place="6" resultid="2214" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2906" daytime="17:04" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1216" daytime="17:06" gender="M" number="60" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1217" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1536" />
                    <RANKING order="2" place="2" resultid="1487" />
                    <RANKING order="3" place="3" resultid="2448" />
                    <RANKING order="4" place="4" resultid="2202" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2907" daytime="17:06" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1218" daytime="17:08" gender="F" number="61" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1219" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2229" />
                    <RANKING order="2" place="2" resultid="2253" />
                    <RANKING order="3" place="3" resultid="2277" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2908" daytime="17:08" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1220" daytime="17:14" gender="F" number="62" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1221" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2710" />
                    <RANKING order="2" place="2" resultid="2230" />
                    <RANKING order="3" place="3" resultid="2254" />
                    <RANKING order="4" place="4" resultid="2465" />
                    <RANKING order="5" place="5" resultid="2527" />
                    <RANKING order="6" place="-1" resultid="2278" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2909" daytime="17:14" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1222" daytime="17:20" gender="M" number="63" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1223" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2237" />
                    <RANKING order="2" place="2" resultid="2470" />
                    <RANKING order="3" place="3" resultid="2261" />
                    <RANKING order="4" place="4" resultid="2285" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2910" daytime="17:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1224" daytime="17:24" gender="M" number="64" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1225" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2238" />
                    <RANKING order="2" place="2" resultid="1393" />
                    <RANKING order="3" place="3" resultid="2262" />
                    <RANKING order="4" place="4" resultid="1561" />
                    <RANKING order="5" place="5" resultid="2286" />
                    <RANKING order="6" place="-1" resultid="2716" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2911" daytime="17:24" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1226" daytime="17:30" gender="F" number="65" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1227" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2228" />
                    <RANKING order="2" place="2" resultid="2464" />
                    <RANKING order="3" place="3" resultid="2252" />
                    <RANKING order="4" place="4" resultid="1389" />
                    <RANKING order="5" place="5" resultid="2709" />
                    <RANKING order="6" place="6" resultid="2276" />
                    <RANKING order="7" place="7" resultid="2478" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2912" daytime="17:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1228" daytime="17:34" gender="F" number="66" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1229" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2231" />
                    <RANKING order="2" place="2" resultid="2255" />
                    <RANKING order="3" place="3" resultid="2466" />
                    <RANKING order="4" place="4" resultid="2279" />
                    <RANKING order="5" place="5" resultid="2711" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2913" daytime="17:34" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1230" daytime="17:38" gender="M" number="67" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1231" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2239" />
                    <RANKING order="2" place="2" resultid="2263" />
                    <RANKING order="3" place="3" resultid="2717" />
                    <RANKING order="4" place="4" resultid="2287" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2914" daytime="17:38" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1232" daytime="17:44" gender="M" number="68" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1233" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2236" />
                    <RANKING order="2" place="2" resultid="2260" />
                    <RANKING order="3" place="3" resultid="1392" />
                    <RANKING order="4" place="4" resultid="2469" />
                    <RANKING order="5" place="5" resultid="2715" />
                    <RANKING order="6" place="6" resultid="1560" />
                    <RANKING order="7" place="7" resultid="2284" />
                    <RANKING order="8" place="8" resultid="1658" />
                    <RANKING order="9" place="9" resultid="1495" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2915" daytime="17:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2916" daytime="17:48" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="2539" nation="BRA" region="PR" clubid="1564" swrid="93771" name="Círculo Militar Do Paraná" shortname="Círculo Militar">
          <ATHLETES>
            <ATHLETE firstname="Rafael" lastname="Cavalcante Pierin" birthdate="2015-03-31" gender="M" nation="BRA" license="408082" swrid="5725986" athleteid="1580" externalid="408082">
              <RESULTS>
                <RESULT eventid="1071" points="116" swimtime="00:03:28.87" resultid="1581" heatid="2742" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                    <SPLIT distance="100" swimtime="00:01:39.36" />
                    <SPLIT distance="150" swimtime="00:02:34.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="83" swimtime="00:00:59.29" resultid="1582" heatid="2759" lane="5" />
                <RESULT eventid="1167" points="98" reactiontime="+70" swimtime="00:00:50.92" resultid="1583" heatid="2854" lane="4" />
                <RESULT eventid="1205" points="110" swimtime="00:00:43.57" resultid="1584" heatid="2888" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Cavalcante Pierin" birthdate="2012-10-30" gender="F" nation="BRA" license="406952" swrid="5717250" athleteid="1575" externalid="406952">
              <RESULTS>
                <RESULT eventid="1074" points="218" swimtime="00:00:48.38" resultid="1576" heatid="2745" lane="2" />
                <RESULT eventid="1158" points="193" swimtime="00:00:42.20" resultid="1577" heatid="2841" lane="7" />
                <RESULT eventid="1192" points="258" swimtime="00:03:18.01" resultid="1578" heatid="2874" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.48" />
                    <SPLIT distance="100" swimtime="00:01:35.89" />
                    <SPLIT distance="150" swimtime="00:02:31.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="285" swimtime="00:00:35.86" resultid="1579" heatid="2894" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Vieira Coelho" birthdate="2014-09-28" gender="F" nation="BRA" license="406951" swrid="5717301" athleteid="1570" externalid="406951">
              <RESULTS>
                <RESULT eventid="1080" points="158" swimtime="00:00:53.92" resultid="1571" heatid="2753" lane="4" />
                <RESULT eventid="1152" points="144" swimtime="00:04:00.12" resultid="1572" heatid="2835" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.49" />
                    <SPLIT distance="100" swimtime="00:02:00.93" />
                    <SPLIT distance="150" swimtime="00:03:08.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1106" points="96" swimtime="00:00:53.23" resultid="1573" heatid="2782" lane="1" />
                <RESULT eventid="1122" points="178" swimtime="00:01:31.81" resultid="1574" heatid="2799" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arya" lastname="Zgoda De Brito Afonso" birthdate="2013-01-03" gender="F" nation="BRA" license="378331" swrid="5588976" athleteid="1565" externalid="378331">
              <RESULTS>
                <RESULT eventid="1086" points="143" swimtime="00:01:49.47" resultid="1566" heatid="2764" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="143" swimtime="00:00:55.71" resultid="1567" heatid="2746" lane="6" entrytime="00:00:52.92" entrycourse="LCM" />
                <RESULT eventid="1132" points="190" swimtime="00:01:29.82" resultid="1568" heatid="2814" lane="2" entrytime="00:01:26.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="181" swimtime="00:00:47.46" resultid="1569" heatid="2790" lane="5" entrytime="00:00:45.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2416" nation="BRA" region="PR" clubid="1277" swrid="93758" name="Apan/Maringá">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Luiza Rampasi" birthdate="2013-10-16" gender="F" nation="BRA" license="382209" swrid="5603866" athleteid="1313" externalid="382209">
              <RESULTS>
                <RESULT eventid="1158" points="100" swimtime="00:00:52.61" resultid="1314" heatid="2842" lane="1" entrytime="00:00:55.79" entrycourse="LCM" />
                <RESULT eventid="1132" points="186" swimtime="00:01:30.56" resultid="1315" heatid="2812" lane="5" entrytime="00:01:43.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="111" swimtime="00:01:55.14" resultid="1316" heatid="2775" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="165" swimtime="00:03:49.83" resultid="1317" heatid="2874" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.78" />
                    <SPLIT distance="100" swimtime="00:02:01.89" />
                    <SPLIT distance="150" swimtime="00:03:02.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Constantino" birthdate="2012-06-02" gender="F" nation="BRA" license="382208" swrid="5420069" athleteid="1308" externalid="382208">
              <RESULTS>
                <RESULT eventid="1074" points="261" swimtime="00:00:45.59" resultid="1309" heatid="2747" lane="8" entrytime="00:00:49.19" entrycourse="LCM" />
                <RESULT eventid="1132" points="260" swimtime="00:01:21.01" resultid="1310" heatid="2814" lane="6" entrytime="00:01:24.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="226" swimtime="00:01:45.19" resultid="1311" heatid="2860" lane="4" entrytime="00:01:56.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="351" swimtime="00:00:33.44" resultid="1312" heatid="2897" lane="4" entrytime="00:00:37.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Baldo De França" birthdate="2014-04-21" gender="M" nation="BRA" license="393773" swrid="5507467" athleteid="1353" externalid="393773">
              <RESULTS>
                <RESULT eventid="1083" points="85" swimtime="00:00:58.88" resultid="1354" heatid="2761" lane="2" entrytime="00:01:04.04" entrycourse="LCM" />
                <RESULT eventid="1155" points="89" swimtime="00:04:14.55" resultid="1355" heatid="2837" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.92" />
                    <SPLIT distance="100" swimtime="00:02:04.24" />
                    <SPLIT distance="150" swimtime="00:03:13.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="77" swimtime="00:00:52.33" resultid="1356" heatid="2785" lane="6" entrytime="00:01:12.84" entrycourse="LCM" />
                <RESULT eventid="1205" points="87" swimtime="00:00:47.13" resultid="1357" heatid="2891" lane="5" entrytime="00:00:46.26" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Otavio Luz" birthdate="2013-07-27" gender="M" nation="BRA" license="392111" swrid="5603882" athleteid="1348" externalid="392111">
              <RESULTS>
                <RESULT eventid="1161" points="172" swimtime="00:00:40.01" resultid="1349" heatid="2845" lane="4" entrytime="00:00:47.30" entrycourse="LCM" />
                <RESULT eventid="1135" points="200" swimtime="00:01:20.06" resultid="1350" heatid="2819" lane="3" entrytime="00:01:29.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="153" swimtime="00:01:32.37" resultid="1351" heatid="2778" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="217" swimtime="00:00:34.79" resultid="1352" heatid="2903" lane="1" entrytime="00:00:38.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Bernardo Padua" birthdate="2013-07-15" gender="M" nation="BRA" license="392108" swrid="5305422" athleteid="1338" externalid="392108">
              <RESULTS>
                <RESULT eventid="1077" points="178" swimtime="00:00:46.05" resultid="1339" heatid="2750" lane="2" entrytime="00:00:51.48" entrycourse="LCM" />
                <RESULT eventid="1135" points="165" swimtime="00:01:25.38" resultid="1340" heatid="2819" lane="6" entrytime="00:01:29.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="159" swimtime="00:01:44.90" resultid="1341" heatid="2862" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="195" swimtime="00:00:36.01" resultid="1342" heatid="2902" lane="1" entrytime="00:00:43.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Pacheco" birthdate="2012-10-03" gender="M" nation="BRA" license="370663" swrid="5603883" athleteid="1283" externalid="370663">
              <RESULTS>
                <RESULT eventid="1089" points="193" swimtime="00:01:29.17" resultid="1284" heatid="2766" lane="5" />
                <RESULT eventid="1161" points="146" swimtime="00:00:42.26" resultid="1285" heatid="2847" lane="8" entrytime="00:00:41.05" entrycourse="LCM" />
                <RESULT eventid="1119" points="157" swimtime="00:00:43.61" resultid="1286" heatid="2794" lane="4" entrytime="00:00:45.86" entrycourse="LCM" />
                <RESULT eventid="1211" points="253" swimtime="00:00:33.03" resultid="1287" heatid="2904" lane="3" entrytime="00:00:33.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Pastre" birthdate="2014-03-10" gender="F" nation="BRA" license="403760" swrid="5684593" athleteid="1378" externalid="403760">
              <RESULTS>
                <RESULT eventid="1068" points="170" swimtime="00:03:23.35" resultid="1379" heatid="2739" lane="5" />
                <RESULT eventid="1106" points="154" swimtime="00:00:45.51" resultid="1380" heatid="2781" lane="2" />
                <RESULT eventid="1164" points="247" reactiontime="+65" swimtime="00:00:42.78" resultid="1381" heatid="2851" lane="5" entrytime="00:00:57.72" entrycourse="LCM" />
                <RESULT eventid="1202" points="170" swimtime="00:00:42.57" resultid="1382" heatid="2885" lane="2" entrytime="00:00:48.47" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raphael" lastname="Piai Pellegrini" birthdate="2012-03-24" gender="M" nation="BRA" license="377261" swrid="5603894" athleteid="1293" externalid="377261">
              <RESULTS>
                <RESULT eventid="1161" points="254" swimtime="00:00:35.16" resultid="1294" heatid="2847" lane="6" entrytime="00:00:37.50" entrycourse="LCM" />
                <RESULT eventid="1135" points="345" swimtime="00:01:06.79" resultid="1295" heatid="2821" lane="7" entrytime="00:01:13.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="251" swimtime="00:00:37.31" resultid="1296" heatid="2793" lane="8" />
                <RESULT eventid="1211" points="353" swimtime="00:00:29.58" resultid="1297" heatid="2905" lane="6" entrytime="00:00:32.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrielle" lastname="Borba" birthdate="2014-06-15" gender="F" nation="BRA" license="385705" swrid="5323267" athleteid="1318" externalid="385705">
              <RESULTS>
                <RESULT eventid="1080" points="130" swimtime="00:00:57.42" resultid="1319" heatid="2756" lane="8" entrytime="00:00:59.67" entrycourse="LCM" />
                <RESULT eventid="1152" points="135" swimtime="00:04:05.72" resultid="1320" heatid="2836" lane="1" entrytime="00:04:22.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.83" />
                    <SPLIT distance="100" swimtime="00:02:01.07" />
                    <SPLIT distance="150" swimtime="00:03:09.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1122" points="159" swimtime="00:01:35.42" resultid="1321" heatid="2801" lane="8" entrytime="00:01:46.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="164" swimtime="00:00:43.13" resultid="1322" heatid="2886" lane="1" entrytime="00:00:44.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Novak Pinho" birthdate="2012-11-14" gender="M" nation="BRA" license="378199" swrid="5603879" athleteid="1303" externalid="378199">
              <RESULTS>
                <RESULT eventid="1089" points="181" swimtime="00:01:31.14" resultid="1304" heatid="2768" lane="1" entrytime="00:01:33.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1149" points="186" swimtime="00:02:58.48" resultid="1305" heatid="2832" lane="6" entrytime="00:03:01.74" entrycourse="LCM" />
                <RESULT eventid="1119" points="174" swimtime="00:00:42.17" resultid="1306" heatid="2795" lane="2" entrytime="00:00:44.06" entrycourse="LCM" />
                <RESULT eventid="1211" points="206" swimtime="00:00:35.36" resultid="1307" heatid="2903" lane="2" entrytime="00:00:36.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Peroni Passafaro" birthdate="2013-09-17" gender="F" nation="BRA" license="370659" swrid="5603893" athleteid="1278" externalid="370659">
              <RESULTS>
                <RESULT eventid="1086" points="179" swimtime="00:01:41.67" resultid="1279" heatid="2764" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="162" swimtime="00:00:44.78" resultid="1280" heatid="2842" lane="4" entrytime="00:00:47.47" entrycourse="LCM" />
                <RESULT eventid="1132" points="212" swimtime="00:01:26.70" resultid="1281" heatid="2814" lane="8" entrytime="00:01:28.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="192" swimtime="00:03:38.54" resultid="1282" heatid="2874" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.16" />
                    <SPLIT distance="100" swimtime="00:01:43.17" />
                    <SPLIT distance="150" swimtime="00:02:53.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Catarina" lastname="Wendt Jesus" birthdate="2013-07-09" gender="F" nation="BRA" license="393778" swrid="5641780" athleteid="1358" externalid="393778">
              <RESULTS>
                <RESULT eventid="1074" points="320" swimtime="00:00:42.60" resultid="1359" heatid="2747" lane="7" entrytime="00:00:46.28" entrycourse="LCM" />
                <RESULT eventid="1132" points="367" swimtime="00:01:12.16" resultid="1360" heatid="2811" lane="6" />
                <RESULT eventid="1170" points="312" swimtime="00:01:34.54" resultid="1361" heatid="2860" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="386" swimtime="00:00:32.41" resultid="1362" heatid="2899" lane="1" entrytime="00:00:35.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lavinia" lastname="Bossoni" birthdate="2013-11-03" gender="F" nation="BRA" license="377260" swrid="5343093" athleteid="1288" externalid="377260">
              <RESULTS>
                <RESULT eventid="1086" points="166" swimtime="00:01:44.27" resultid="1289" heatid="2764" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="175" swimtime="00:03:21.55" resultid="1290" heatid="2828" lane="2" />
                <RESULT eventid="1132" points="184" swimtime="00:01:30.90" resultid="1291" heatid="2813" lane="7" entrytime="00:01:38.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="170" swimtime="00:03:47.32" resultid="1292" heatid="2875" lane="7" entrytime="00:04:13.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.86" />
                    <SPLIT distance="150" swimtime="00:02:56.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Dos Reis Monteiro" birthdate="2014-08-05" gender="M" nation="BRA" license="392095" swrid="5697226" athleteid="1323" externalid="392095">
              <RESULTS>
                <RESULT eventid="1071" points="219" swimtime="00:02:49.12" resultid="1324" heatid="2741" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.31" />
                    <SPLIT distance="150" swimtime="00:02:05.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="203" swimtime="00:03:13.83" resultid="1325" heatid="2839" lane="5" entrytime="00:03:25.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                    <SPLIT distance="100" swimtime="00:01:35.26" />
                    <SPLIT distance="150" swimtime="00:02:32.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="168" swimtime="00:00:40.32" resultid="1326" heatid="2786" lane="5" entrytime="00:00:40.97" entrycourse="LCM" />
                <RESULT eventid="1205" points="257" swimtime="00:00:32.86" resultid="1327" heatid="2893" lane="4" entrytime="00:00:34.36" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Muniz" birthdate="2012-09-03" gender="M" nation="BRA" license="392106" swrid="5603877" athleteid="1333" externalid="392106">
              <RESULTS>
                <RESULT eventid="1089" points="91" swimtime="00:01:54.43" resultid="1334" heatid="2767" lane="6" />
                <RESULT eventid="1161" points="101" swimtime="00:00:47.68" resultid="1335" heatid="2845" lane="3" entrytime="00:01:00.29" entrycourse="LCM" />
                <RESULT eventid="1119" points="84" swimtime="00:00:53.75" resultid="1336" heatid="2792" lane="3" />
                <RESULT eventid="1211" points="163" swimtime="00:00:38.26" resultid="1337" heatid="2902" lane="7" entrytime="00:00:43.26" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Rafael Padial" birthdate="2014-03-07" gender="M" nation="BRA" license="397331" swrid="5641774" athleteid="1363" externalid="397331">
              <RESULTS>
                <RESULT eventid="1083" points="108" swimtime="00:00:54.40" resultid="1364" heatid="2762" lane="1" entrytime="00:00:56.92" entrycourse="LCM" />
                <RESULT eventid="1109" points="110" swimtime="00:00:46.39" resultid="1365" heatid="2786" lane="7" entrytime="00:00:49.48" entrycourse="LCM" />
                <RESULT eventid="1167" status="DNS" swimtime="00:00:00.00" resultid="1366" heatid="2857" lane="4" entrytime="00:00:51.94" entrycourse="LCM" />
                <RESULT eventid="1205" points="202" swimtime="00:00:35.62" resultid="1367" heatid="2893" lane="6" entrytime="00:00:38.32" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="De Correa" birthdate="2014-12-03" gender="M" nation="BRA" license="403387" swrid="5676286" athleteid="1373" externalid="403387">
              <RESULTS>
                <RESULT eventid="1071" points="108" swimtime="00:03:33.68" resultid="1374" heatid="2741" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.66" />
                    <SPLIT distance="150" swimtime="00:02:36.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="109" reactiontime="+75" swimtime="00:00:49.22" resultid="1375" heatid="2857" lane="2" entrytime="00:00:54.97" entrycourse="LCM" />
                <RESULT eventid="1125" points="118" swimtime="00:01:35.34" resultid="1376" heatid="2808" lane="1" entrytime="00:01:39.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="120" swimtime="00:00:42.30" resultid="1377" heatid="2892" lane="7" entrytime="00:00:43.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Tomazeli" birthdate="2013-02-05" gender="M" nation="BRA" license="392109" swrid="5614097" athleteid="1343" externalid="392109">
              <RESULTS>
                <RESULT eventid="1089" points="113" swimtime="00:01:46.60" resultid="1344" heatid="2767" lane="1" />
                <RESULT eventid="1161" points="94" swimtime="00:00:48.86" resultid="1345" heatid="2845" lane="5" entrytime="00:00:51.17" entrycourse="LCM" />
                <RESULT eventid="1119" points="119" swimtime="00:00:47.76" resultid="1346" heatid="2794" lane="3" entrytime="00:00:47.54" entrycourse="LCM" />
                <RESULT eventid="1211" points="159" swimtime="00:00:38.54" resultid="1347" heatid="2902" lane="5" entrytime="00:00:39.94" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Santos Carraro" birthdate="2014-06-04" gender="M" nation="BRA" license="392097" swrid="5603908" athleteid="1328" externalid="392097">
              <RESULTS>
                <RESULT eventid="1071" points="174" swimtime="00:03:02.36" resultid="1329" heatid="2743" lane="2" entrytime="00:03:25.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="100" swimtime="00:01:26.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="86" swimtime="00:00:50.31" resultid="1330" heatid="2786" lane="1" entrytime="00:00:51.62" entrycourse="LCM" />
                <RESULT eventid="1167" points="93" reactiontime="+65" swimtime="00:00:51.93" resultid="1331" heatid="2858" lane="1" entrytime="00:00:50.25" entrycourse="LCM" />
                <RESULT eventid="1205" points="146" swimtime="00:00:39.69" resultid="1332" heatid="2893" lane="8" entrytime="00:00:39.82" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Ayres" birthdate="2012-05-05" gender="M" nation="BRA" license="378035" swrid="5208079" athleteid="1298" externalid="378035">
              <RESULTS>
                <RESULT eventid="1089" points="302" swimtime="00:01:16.84" resultid="1299" heatid="2766" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="293" swimtime="00:00:33.52" resultid="1300" heatid="2847" lane="3" entrytime="00:00:35.32" entrycourse="LCM" />
                <RESULT eventid="1119" points="283" swimtime="00:00:35.83" resultid="1301" heatid="2796" lane="6" entrytime="00:00:39.02" entrycourse="LCM" />
                <RESULT eventid="1211" points="324" swimtime="00:00:30.44" resultid="1302" heatid="2905" lane="3" entrytime="00:00:31.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Yukio Tacaiama" birthdate="2014-06-29" gender="M" nation="BRA" license="407184" swrid="5718894" athleteid="1383" externalid="407184">
              <RESULTS>
                <RESULT eventid="1083" points="115" swimtime="00:00:53.23" resultid="1384" heatid="2758" lane="4" />
                <RESULT eventid="1155" points="124" swimtime="00:03:48.60" resultid="1385" heatid="2837" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.39" />
                    <SPLIT distance="100" swimtime="00:01:55.32" />
                    <SPLIT distance="150" swimtime="00:03:00.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="133" swimtime="00:01:31.78" resultid="1386" heatid="2803" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="143" swimtime="00:00:39.97" resultid="1387" heatid="2887" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Arthur Da Silva Ortiz" birthdate="2015-04-20" gender="M" nation="BRA" license="399733" swrid="5676285" athleteid="1368" externalid="399733">
              <RESULTS>
                <RESULT eventid="1083" points="85" swimtime="00:00:58.90" resultid="1369" heatid="2760" lane="2" entrytime="00:01:12.11" entrycourse="LCM" />
                <RESULT eventid="1155" points="96" swimtime="00:04:08.88" resultid="1370" heatid="2838" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.54" />
                    <SPLIT distance="150" swimtime="00:03:12.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="98" swimtime="00:01:41.53" resultid="1371" heatid="2804" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="103" swimtime="00:00:44.51" resultid="1372" heatid="2890" lane="2" entrytime="00:01:21.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1182" points="172" swimtime="00:02:32.41" resultid="1390" heatid="2868" lane="3" entrytime="00:02:30.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1373" number="1" />
                    <RELAYPOSITION athleteid="1328" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1383" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1323" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1224" points="146" reactiontime="+66" swimtime="00:02:56.90" resultid="1393" heatid="2911" lane="3" entrytime="00:02:59.10">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:17.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1363" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="1323" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1328" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1383" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1190" points="280" swimtime="00:02:09.63" resultid="1391" heatid="2873" lane="2" entrytime="00:02:12.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1283" number="1" />
                    <RELAYPOSITION athleteid="1303" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1293" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1298" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1232" points="224" reactiontime="+82" swimtime="00:02:33.34" resultid="1392" heatid="2916" lane="6" entrytime="00:02:32.67">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1298" number="1" reactiontime="+82" />
                    <RELAYPOSITION athleteid="1283" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1293" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1303" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="F" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1184" points="252" swimtime="00:02:30.75" resultid="1388" heatid="2869" lane="2" entrytime="00:02:45.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.20" />
                    <SPLIT distance="100" swimtime="00:01:20.88" />
                    <SPLIT distance="150" swimtime="00:01:58.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1288" number="1" />
                    <RELAYPOSITION athleteid="1313" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1278" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1358" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1226" points="215" reactiontime="+72" swimtime="00:02:56.27" resultid="1389" heatid="2912" lane="2" entrytime="00:03:08.05">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1288" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="1358" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1278" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1313" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1096" swimtime="00:02:29.53" resultid="1394" heatid="2772" lane="2" entrytime="00:02:17.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                    <SPLIT distance="100" swimtime="00:01:17.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1288" number="1" />
                    <RELAYPOSITION athleteid="1278" number="2" />
                    <RELAYPOSITION athleteid="1343" number="3" />
                    <RELAYPOSITION athleteid="1348" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1142" swimtime="00:02:56.33" resultid="1399" heatid="2825" lane="2" entrytime="00:02:44.54">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1278" number="1" />
                    <RELAYPOSITION athleteid="1338" number="2" />
                    <RELAYPOSITION athleteid="1348" number="3" />
                    <RELAYPOSITION athleteid="1288" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1098" swimtime="00:02:07.10" resultid="1395" heatid="2774" lane="3" entrytime="00:02:10.32">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1293" number="1" />
                    <RELAYPOSITION athleteid="1308" number="2" />
                    <RELAYPOSITION athleteid="1358" number="3" />
                    <RELAYPOSITION athleteid="1298" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1144" swimtime="00:02:33.39" resultid="1397" heatid="2827" lane="3" entrytime="00:02:23.78">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1298" number="1" />
                    <RELAYPOSITION athleteid="1308" number="2" />
                    <RELAYPOSITION athleteid="1293" number="3" />
                    <RELAYPOSITION athleteid="1358" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1094" swimtime="00:02:33.73" resultid="1396" heatid="2771" lane="2" entrytime="00:02:31.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.28" />
                    <SPLIT distance="100" swimtime="00:01:18.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1363" number="1" />
                    <RELAYPOSITION athleteid="1378" number="2" />
                    <RELAYPOSITION athleteid="1318" number="3" />
                    <RELAYPOSITION athleteid="1323" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1140" swimtime="00:02:58.73" resultid="1398" heatid="2824" lane="2" entrytime="00:02:54.67">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1378" number="1" />
                    <RELAYPOSITION athleteid="1323" number="2" />
                    <RELAYPOSITION athleteid="1328" number="3" />
                    <RELAYPOSITION athleteid="1318" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="16131" nation="BRA" region="PR" clubid="2296" swrid="93766" name="Associação Nadar Colombo" shortname="Equipe Nadar">
          <ATHLETES>
            <ATHLETE firstname="Tayna" lastname="Macedo Gabardo" birthdate="2012-12-01" gender="F" nation="BRA" license="406704" swrid="5717281" athleteid="2297" externalid="406704">
              <RESULTS>
                <RESULT eventid="1192" points="192" swimtime="00:03:38.52" resultid="2298" heatid="2874" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.59" />
                    <SPLIT distance="100" swimtime="00:01:48.57" />
                    <SPLIT distance="150" swimtime="00:02:49.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="254" swimtime="00:00:37.23" resultid="2299" heatid="2894" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13068" nation="BRA" region="PR" clubid="2481" swrid="93787" name="Sociedade Morgenau" shortname="Morgenau">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Fernanda De Lima" birthdate="2013-09-26" gender="F" nation="BRA" license="378290" swrid="5588693" athleteid="2487" externalid="378290">
              <RESULTS>
                <RESULT eventid="1074" points="107" swimtime="00:01:01.33" resultid="2488" heatid="2745" lane="7" />
                <RESULT eventid="1132" points="169" swimtime="00:01:33.38" resultid="2489" heatid="2812" lane="4" entrytime="00:01:40.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="185" swimtime="00:00:47.12" resultid="2490" heatid="2790" lane="1" entrytime="00:00:49.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Paes Pereira" birthdate="2013-03-11" gender="M" nation="BRA" license="391137" swrid="5602567" athleteid="2491" externalid="391137">
              <RESULTS>
                <RESULT eventid="1149" points="91" swimtime="00:03:46.13" resultid="2492" heatid="2831" lane="2" />
                <RESULT eventid="1135" points="91" swimtime="00:01:44.10" resultid="2493" heatid="2818" lane="2" entrytime="00:01:44.28" entrycourse="LCM" />
                <RESULT eventid="1119" points="98" swimtime="00:00:51.05" resultid="2494" heatid="2794" lane="1" entrytime="00:00:51.71" entrycourse="LCM" />
                <RESULT eventid="1211" points="110" swimtime="00:00:43.52" resultid="2495" heatid="2901" lane="4" entrytime="00:00:45.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Tomaz Zmievski" birthdate="2012-09-20" gender="F" nation="BRA" license="406725" swrid="5717300" athleteid="2521" externalid="406725">
              <RESULTS>
                <RESULT eventid="1074" points="128" swimtime="00:00:57.83" resultid="2522" heatid="2744" lane="4" />
                <RESULT eventid="1146" points="173" swimtime="00:03:22.37" resultid="2523" heatid="2828" lane="8" />
                <RESULT eventid="1158" points="103" swimtime="00:00:52.06" resultid="2524" heatid="2841" lane="2" />
                <RESULT eventid="1132" points="211" swimtime="00:01:26.76" resultid="2525" heatid="2812" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Felipe Kuhn" birthdate="2014-03-22" gender="M" nation="BRA" license="392121" swrid="5602536" athleteid="2496" externalid="392121">
              <RESULTS>
                <RESULT eventid="1083" points="138" swimtime="00:00:50.20" resultid="2497" heatid="2758" lane="2" />
                <RESULT eventid="1205" points="143" swimtime="00:00:39.93" resultid="2498" heatid="2888" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Alves" birthdate="2012-10-12" gender="M" nation="BRA" license="369324" swrid="5588674" athleteid="2482" externalid="369324">
              <RESULTS>
                <RESULT eventid="1089" points="268" swimtime="00:01:19.94" resultid="2483" heatid="2768" lane="3" entrytime="00:01:28.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" status="DSQ" swimtime="00:00:35.95" resultid="2484" heatid="2846" lane="6" entrytime="00:00:42.45" entrycourse="LCM" />
                <RESULT eventid="1119" points="281" swimtime="00:00:35.95" resultid="2485" heatid="2796" lane="2" entrytime="00:00:39.31" entrycourse="LCM" />
                <RESULT eventid="1195" points="209" swimtime="00:03:11.81" resultid="2486" heatid="2877" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                    <SPLIT distance="100" swimtime="00:01:28.03" />
                    <SPLIT distance="150" swimtime="00:02:31.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Melo" birthdate="2015-02-07" gender="F" nation="BRA" license="406717" swrid="5717280" athleteid="2508" externalid="406717">
              <RESULTS>
                <RESULT eventid="1068" points="140" swimtime="00:03:37.05" resultid="2509" heatid="2738" lane="7" />
                <RESULT eventid="1106" points="113" swimtime="00:00:50.43" resultid="2510" heatid="2780" lane="6" />
                <RESULT eventid="1164" points="167" swimtime="00:00:48.72" resultid="2511" heatid="2848" lane="5" />
                <RESULT eventid="1202" points="150" swimtime="00:00:44.38" resultid="2512" heatid="2884" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Nitz Costa" birthdate="2015-02-09" gender="F" nation="BRA" license="397328" swrid="5641773" athleteid="2499" externalid="397328">
              <RESULTS>
                <RESULT eventid="1068" points="178" swimtime="00:03:20.33" resultid="2500" heatid="2738" lane="5" />
                <RESULT eventid="1106" points="140" swimtime="00:00:47.00" resultid="2501" heatid="2783" lane="7" entrytime="00:00:59.23" entrycourse="LCM" />
                <RESULT eventid="1164" points="189" reactiontime="+39" swimtime="00:00:46.75" resultid="2502" heatid="2852" lane="5" entrytime="00:00:49.70" entrycourse="LCM" />
                <RESULT eventid="1122" points="174" swimtime="00:01:32.45" resultid="2503" heatid="2799" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maryana" lastname="Lemos Carvalho" birthdate="2014-02-10" gender="F" nation="BRA" license="406718" swrid="5717278" athleteid="2513" externalid="406718">
              <RESULTS>
                <RESULT eventid="1068" points="91" swimtime="00:04:10.43" resultid="2514" heatid="2739" lane="7" />
                <RESULT eventid="1164" points="107" reactiontime="+65" swimtime="00:00:56.54" resultid="2515" heatid="2850" lane="3" />
                <RESULT eventid="1122" points="119" swimtime="00:01:45.04" resultid="2516" heatid="2800" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="145" swimtime="00:00:44.87" resultid="2517" heatid="2884" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cecilia Carstens" birthdate="2014-02-22" gender="F" nation="BRA" license="406721" swrid="5717251" athleteid="2518" externalid="406721">
              <RESULTS>
                <RESULT eventid="1106" points="81" swimtime="00:00:56.35" resultid="2519" heatid="2780" lane="3" />
                <RESULT eventid="1122" points="114" swimtime="00:01:46.50" resultid="2520" heatid="2797" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Lara" birthdate="2014-09-02" gender="F" nation="BRA" license="406686" swrid="5717259" athleteid="2504" externalid="406686">
              <RESULTS>
                <RESULT eventid="1152" points="96" swimtime="00:04:34.55" resultid="2505" heatid="2835" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.36" />
                    <SPLIT distance="100" swimtime="00:02:12.83" />
                    <SPLIT distance="150" swimtime="00:03:37.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="86" reactiontime="+82" swimtime="00:01:00.73" resultid="2506" heatid="2850" lane="1" />
                <RESULT eventid="1202" points="151" swimtime="00:00:44.24" resultid="2507" heatid="2883" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="F" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1178" points="156" swimtime="00:02:57.02" resultid="2526" heatid="2866" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                    <SPLIT distance="100" swimtime="00:01:26.52" />
                    <SPLIT distance="150" swimtime="00:02:12.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2499" number="1" />
                    <RELAYPOSITION athleteid="2504" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2508" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2513" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1220" points="108" reactiontime="+63" swimtime="00:03:41.57" resultid="2527" heatid="2909" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.80" />
                    <SPLIT distance="100" swimtime="00:02:15.56" />
                    <SPLIT distance="150" swimtime="00:02:53.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2513" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="2508" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2499" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2504" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="X" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1144" swimtime="00:03:07.17" resultid="2528" heatid="2826" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2491" number="1" />
                    <RELAYPOSITION athleteid="2521" number="2" />
                    <RELAYPOSITION athleteid="2482" number="3" />
                    <RELAYPOSITION athleteid="2487" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="36" nation="BRA" region="PR" clubid="1601" swrid="93753" name="Associação Atlética Comercial" shortname="Comercial Cascavel">
          <ATHLETES>
            <ATHLETE firstname="Marianna" lastname="Galvao Oliveira" birthdate="2014-03-18" gender="F" nation="BRA" license="390835" swrid="5596902" athleteid="1627" externalid="390835">
              <RESULTS>
                <RESULT eventid="1080" points="206" swimtime="00:00:49.32" resultid="1628" heatid="2756" lane="2" entrytime="00:00:56.53" entrycourse="LCM" />
                <RESULT eventid="1152" points="165" swimtime="00:03:49.57" resultid="1629" heatid="2836" lane="6" entrytime="00:04:12.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:54.83" />
                    <SPLIT distance="150" swimtime="00:02:58.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1106" points="108" swimtime="00:00:51.21" resultid="1630" heatid="2783" lane="2" entrytime="00:00:56.30" entrycourse="LCM" />
                <RESULT eventid="1164" points="153" swimtime="00:00:50.15" resultid="1631" heatid="2851" lane="6" entrytime="00:00:59.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Pedro Serafini" birthdate="2012-05-15" gender="M" nation="BRA" license="365488" swrid="5596924" athleteid="1617" externalid="365488">
              <RESULTS>
                <RESULT eventid="1149" points="214" swimtime="00:02:50.42" resultid="1618" heatid="2832" lane="2" entrytime="00:03:01.79" entrycourse="LCM" />
                <RESULT eventid="1161" points="161" swimtime="00:00:40.86" resultid="1619" heatid="2845" lane="2" />
                <RESULT eventid="1135" points="201" swimtime="00:01:19.94" resultid="1620" heatid="2820" lane="1" entrytime="00:01:20.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="182" swimtime="00:03:20.98" resultid="1621" heatid="2878" lane="6" entrytime="00:03:26.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.65" />
                    <SPLIT distance="100" swimtime="00:01:39.74" />
                    <SPLIT distance="150" swimtime="00:02:40.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose" lastname="Eliziario Filho" birthdate="2014-03-27" gender="M" nation="BRA" license="406696" swrid="4979701" athleteid="1652" externalid="406696">
              <RESULTS>
                <RESULT eventid="1109" points="120" swimtime="00:00:45.10" resultid="1653" heatid="2784" lane="6" />
                <RESULT eventid="1167" points="116" reactiontime="+48" swimtime="00:00:48.25" resultid="1654" heatid="2854" lane="3" />
                <RESULT eventid="1125" points="134" swimtime="00:01:31.44" resultid="1655" heatid="2803" lane="8" />
                <RESULT eventid="1205" points="144" swimtime="00:00:39.89" resultid="1656" heatid="2887" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Vieira Rohnelt" birthdate="2012-05-03" gender="M" nation="BRA" license="365692" swrid="5588952" athleteid="1602" externalid="365692">
              <RESULTS>
                <RESULT eventid="1077" points="160" swimtime="00:00:47.72" resultid="1603" heatid="2750" lane="6" entrytime="00:00:49.85" entrycourse="LCM" />
                <RESULT eventid="1161" points="151" swimtime="00:00:41.79" resultid="1604" heatid="2845" lane="7" />
                <RESULT eventid="1103" points="149" swimtime="00:01:33.11" resultid="1605" heatid="2779" lane="2" entrytime="00:01:43.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="203" swimtime="00:03:13.89" resultid="1606" heatid="2879" lane="1" entrytime="00:03:20.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.65" />
                    <SPLIT distance="100" swimtime="00:01:36.34" />
                    <SPLIT distance="150" swimtime="00:02:31.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Henrique Marca Dos Santos" birthdate="2015-03-28" gender="M" nation="BRA" license="406695" swrid="4991165" athleteid="1647" externalid="406695">
              <RESULTS>
                <RESULT eventid="1083" points="34" swimtime="00:01:19.45" resultid="1648" heatid="2759" lane="8" />
                <RESULT eventid="1109" points="114" swimtime="00:00:45.87" resultid="1649" heatid="2785" lane="8" />
                <RESULT eventid="1167" points="137" reactiontime="+74" swimtime="00:00:45.66" resultid="1650" heatid="2856" lane="2" />
                <RESULT eventid="1205" points="157" swimtime="00:00:38.76" resultid="1651" heatid="2889" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Macedo Medeiros" birthdate="2012-05-12" gender="M" nation="BRA" license="392015" swrid="4697574" athleteid="1642" externalid="392015">
              <RESULTS>
                <RESULT eventid="1077" points="166" swimtime="00:00:47.19" resultid="1643" heatid="2749" lane="5" entrytime="00:00:54.05" entrycourse="LCM" />
                <RESULT eventid="1103" points="97" swimtime="00:01:47.56" resultid="1644" heatid="2778" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="162" swimtime="00:01:44.13" resultid="1645" heatid="2864" lane="8" entrytime="00:01:59.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="176" swimtime="00:03:23.10" resultid="1646" heatid="2878" lane="7" entrytime="00:03:34.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.57" />
                    <SPLIT distance="100" swimtime="00:01:43.59" />
                    <SPLIT distance="150" swimtime="00:02:38.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabelle" lastname="Cordeiro Silva" birthdate="2015-06-14" gender="F" nation="BRA" license="390839" swrid="5596878" athleteid="1632" externalid="390839">
              <RESULTS>
                <RESULT eventid="1068" points="138" swimtime="00:03:38.19" resultid="1633" heatid="2737" lane="5" />
                <RESULT eventid="1080" points="136" swimtime="00:00:56.68" resultid="1634" heatid="2756" lane="7" entrytime="00:00:58.60" entrycourse="LCM" />
                <RESULT eventid="1152" points="148" swimtime="00:03:58.35" resultid="1635" heatid="2835" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:58.79" />
                    <SPLIT distance="150" swimtime="00:03:04.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1106" points="75" swimtime="00:00:57.70" resultid="1636" heatid="2783" lane="3" entrytime="00:00:55.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Vargas Moreira" birthdate="2014-03-09" gender="F" nation="BRA" license="392014" swrid="4904290" athleteid="1637" externalid="392014">
              <RESULTS>
                <RESULT eventid="1068" points="265" swimtime="00:02:55.65" resultid="1638" heatid="2740" lane="5" entrytime="00:03:11.37" entrycourse="LCM" />
                <RESULT eventid="1152" points="205" swimtime="00:03:33.58" resultid="1639" heatid="2836" lane="5" entrytime="00:03:43.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.38" />
                    <SPLIT distance="100" swimtime="00:01:43.89" />
                    <SPLIT distance="150" swimtime="00:02:50.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1122" points="239" swimtime="00:01:23.26" resultid="1640" heatid="2801" lane="5" entrytime="00:01:27.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="231" swimtime="00:00:38.43" resultid="1641" heatid="2886" lane="3" entrytime="00:00:40.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Bonamigo" birthdate="2013-06-25" gender="M" nation="BRA" license="365484" swrid="5588558" athleteid="1622" externalid="365484">
              <RESULTS>
                <RESULT eventid="1065" points="223" swimtime="00:06:02.71" resultid="1623" heatid="2735" lane="6" />
                <RESULT eventid="1077" points="223" swimtime="00:00:42.73" resultid="1624" heatid="2751" lane="3" entrytime="00:00:41.56" entrycourse="LCM" />
                <RESULT eventid="1173" points="242" swimtime="00:01:31.25" resultid="1625" heatid="2863" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="240" swimtime="00:03:03.21" resultid="1626" heatid="2879" lane="3" entrytime="00:03:11.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.14" />
                    <SPLIT distance="100" swimtime="00:01:29.58" />
                    <SPLIT distance="150" swimtime="00:02:21.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Bezerra Sedlacek" birthdate="2014-02-26" gender="M" nation="BRA" license="380663" swrid="4300166" athleteid="1612" externalid="380663">
              <RESULTS>
                <RESULT eventid="1083" points="121" swimtime="00:00:52.41" resultid="1613" heatid="2760" lane="8" />
                <RESULT eventid="1167" points="137" reactiontime="+75" swimtime="00:00:45.62" resultid="1614" heatid="2855" lane="1" />
                <RESULT eventid="1125" points="157" swimtime="00:01:26.78" resultid="1615" heatid="2805" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="155" swimtime="00:00:38.89" resultid="1616" heatid="2888" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Emanuel Rech" birthdate="2013-12-02" gender="M" nation="BRA" license="380660" swrid="5588679" athleteid="1607" externalid="380660">
              <RESULTS>
                <RESULT eventid="1089" points="239" swimtime="00:01:23.10" resultid="1608" heatid="2767" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1149" points="205" swimtime="00:02:52.85" resultid="1609" heatid="2830" lane="3" />
                <RESULT eventid="1119" points="237" swimtime="00:00:38.01" resultid="1610" heatid="2796" lane="5" entrytime="00:00:38.73" entrycourse="LCM" />
                <RESULT eventid="1195" points="206" swimtime="00:03:12.76" resultid="1611" heatid="2879" lane="6" entrytime="00:03:15.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.98" />
                    <SPLIT distance="100" swimtime="00:01:32.53" />
                    <SPLIT distance="150" swimtime="00:02:29.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1190" points="208" swimtime="00:02:23.18" resultid="1657" heatid="2873" lane="4" entrytime="00:01:59.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:11.65" />
                    <SPLIT distance="150" swimtime="00:01:48.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1602" number="1" />
                    <RELAYPOSITION athleteid="1617" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1642" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1622" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1232" points="188" reactiontime="+63" swimtime="00:02:42.68" resultid="1658" heatid="2916" lane="4" entrytime="00:02:14.57">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.51" />
                    <SPLIT distance="150" swimtime="00:02:07.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1607" number="1" reactiontime="+63" />
                    <RELAYPOSITION athleteid="1642" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1617" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1602" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="X" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1094" swimtime="00:02:36.71" resultid="1659" heatid="2771" lane="3" entrytime="00:02:27.49">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1652" number="1" />
                    <RELAYPOSITION athleteid="1627" number="2" />
                    <RELAYPOSITION athleteid="1612" number="3" />
                    <RELAYPOSITION athleteid="1637" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1140" swimtime="00:03:02.66" resultid="1660" heatid="2824" lane="5" entrytime="00:02:45.09">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1612" number="1" />
                    <RELAYPOSITION athleteid="1627" number="2" />
                    <RELAYPOSITION athleteid="1652" number="3" />
                    <RELAYPOSITION athleteid="1637" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="2300" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Bruna" lastname="Scalise Drapzichinski" birthdate="2012-03-07" gender="F" nation="BRA" license="378349" swrid="5603909" athleteid="2321" externalid="378349">
              <RESULTS>
                <RESULT eventid="1074" points="459" swimtime="00:00:37.79" resultid="2322" heatid="2747" lane="5" entrytime="00:00:40.61" entrycourse="LCM" />
                <RESULT eventid="1158" points="300" swimtime="00:00:36.49" resultid="2323" heatid="2841" lane="6" />
                <RESULT eventid="1170" points="421" swimtime="00:01:25.51" resultid="2324" heatid="2861" lane="3" entrytime="00:01:35.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="301" swimtime="00:03:08.15" resultid="2325" heatid="2874" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                    <SPLIT distance="100" swimtime="00:01:30.41" />
                    <SPLIT distance="150" swimtime="00:02:23.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Stephany" birthdate="2012-07-27" gender="F" nation="BRA" license="382210" swrid="5603917" athleteid="2409" externalid="382210">
              <RESULTS>
                <RESULT eventid="1158" points="155" swimtime="00:00:45.41" resultid="2410" heatid="2843" lane="8" entrytime="00:00:46.23" entrycourse="LCM" />
                <RESULT eventid="1100" points="123" swimtime="00:01:51.33" resultid="2411" heatid="2777" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" status="DSQ" swimtime="00:03:47.93" resultid="2412" heatid="2874" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.56" />
                    <SPLIT distance="150" swimtime="00:03:00.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="247" swimtime="00:00:37.59" resultid="2413" heatid="2897" lane="3" entrytime="00:00:40.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Guidin Madureira" birthdate="2015-01-10" gender="M" nation="BRA" license="402116" swrid="5661347" athleteid="2390" externalid="402116">
              <RESULTS>
                <RESULT eventid="1167" status="DNS" swimtime="00:00:00.00" resultid="2391" heatid="2857" lane="6" entrytime="00:00:54.88" entrycourse="LCM" />
                <RESULT eventid="1125" points="109" swimtime="00:01:38.02" resultid="2392" heatid="2804" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="106" swimtime="00:00:44.09" resultid="2393" heatid="2891" lane="8" entrytime="00:00:52.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Bilemjian Leszczynski" birthdate="2014-02-22" gender="M" nation="BRA" license="406924" swrid="5631285" athleteid="2440" externalid="406924">
              <RESULTS>
                <RESULT eventid="1071" points="106" swimtime="00:03:35.00" resultid="2441" heatid="2741" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.76" />
                    <SPLIT distance="150" swimtime="00:02:40.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="73" swimtime="00:01:02.04" resultid="2442" heatid="2758" lane="6" />
                <RESULT eventid="1125" points="103" swimtime="00:01:39.68" resultid="2443" heatid="2803" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="113" swimtime="00:00:43.25" resultid="2444" heatid="2888" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Lima Coelho" birthdate="2012-12-12" gender="M" nation="BRA" license="393775" swrid="5615959" athleteid="2399" externalid="393775">
              <RESULTS>
                <RESULT eventid="1089" points="152" swimtime="00:01:36.60" resultid="2400" heatid="2766" lane="1" />
                <RESULT eventid="1149" points="122" swimtime="00:03:25.43" resultid="2401" heatid="2831" lane="5" />
                <RESULT eventid="1119" points="173" swimtime="00:00:42.25" resultid="2402" heatid="2792" lane="4" />
                <RESULT eventid="1211" points="166" swimtime="00:00:38.04" resultid="2403" heatid="2900" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Gevaerd Verssutti Garcia" birthdate="2013-10-15" gender="F" nation="BRA" license="378404" swrid="5588723" athleteid="2346" externalid="378404">
              <RESULTS>
                <RESULT eventid="1086" points="216" swimtime="00:01:35.45" resultid="2347" heatid="2763" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="241" swimtime="00:01:23.05" resultid="2348" heatid="2814" lane="7" entrytime="00:01:27.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="226" swimtime="00:00:44.06" resultid="2349" heatid="2790" lane="4" entrytime="00:00:44.87" entrycourse="LCM" />
                <RESULT eventid="1208" points="293" swimtime="00:00:35.54" resultid="2350" heatid="2897" lane="5" entrytime="00:00:39.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eloah" lastname="Frasson" birthdate="2012-06-14" gender="F" nation="BRA" license="378338" swrid="5577016" athleteid="2306" externalid="378338">
              <RESULTS>
                <RESULT eventid="1074" points="291" swimtime="00:00:43.99" resultid="2307" heatid="2747" lane="3" entrytime="00:00:42.42" entrycourse="LCM" />
                <RESULT eventid="1132" points="263" swimtime="00:01:20.70" resultid="2308" heatid="2815" lane="8" entrytime="00:01:21.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="256" swimtime="00:01:40.96" resultid="2309" heatid="2861" lane="5" entrytime="00:01:35.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="287" swimtime="00:00:35.78" resultid="2310" heatid="2898" lane="8" entrytime="00:00:37.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabel" lastname="Rezende" birthdate="2013-12-13" gender="F" nation="BRA" license="370657" swrid="5603900" athleteid="2301" externalid="370657">
              <RESULTS>
                <RESULT eventid="1086" points="180" swimtime="00:01:41.38" resultid="2302" heatid="2763" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="164" swimtime="00:00:53.19" resultid="2303" heatid="2745" lane="1" />
                <RESULT eventid="1116" points="207" swimtime="00:00:45.39" resultid="2304" heatid="2789" lane="4" entrytime="00:00:50.41" entrycourse="LCM" />
                <RESULT eventid="1208" points="225" swimtime="00:00:38.78" resultid="2305" heatid="2897" lane="7" entrytime="00:00:41.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Britto" birthdate="2012-10-04" gender="M" nation="BRA" license="378350" swrid="5588566" athleteid="2326" externalid="378350">
              <RESULTS>
                <RESULT eventid="1089" points="242" swimtime="00:01:22.79" resultid="2327" heatid="2768" lane="5" entrytime="00:01:25.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="221" swimtime="00:00:36.83" resultid="2328" heatid="2844" lane="4" />
                <RESULT eventid="1119" points="272" swimtime="00:00:36.34" resultid="2329" heatid="2796" lane="3" entrytime="00:00:38.87" entrycourse="LCM" />
                <RESULT eventid="1195" status="DSQ" swimtime="00:03:09.84" resultid="2330" heatid="2878" lane="3" entrytime="00:03:24.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                    <SPLIT distance="100" swimtime="00:01:27.62" />
                    <SPLIT distance="150" swimtime="00:02:27.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Sprengel Betim" birthdate="2012-08-17" gender="F" nation="BRA" license="385011" swrid="5588922" athleteid="2414" externalid="385011">
              <RESULTS>
                <RESULT eventid="1086" points="218" swimtime="00:01:35.12" resultid="2415" heatid="2765" lane="1" entrytime="00:01:38.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="230" swimtime="00:00:39.84" resultid="2416" heatid="2843" lane="7" entrytime="00:00:44.35" entrycourse="LCM" />
                <RESULT eventid="1132" points="270" swimtime="00:01:20.00" resultid="2417" heatid="2812" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="272" swimtime="00:03:14.61" resultid="2418" heatid="2875" lane="4" entrytime="00:03:37.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.15" />
                    <SPLIT distance="100" swimtime="00:01:37.70" />
                    <SPLIT distance="150" swimtime="00:02:34.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Schneider Yazbek" birthdate="2013-03-07" gender="F" nation="BRA" license="378329" swrid="5588907" athleteid="2376" externalid="378329">
              <RESULTS>
                <RESULT eventid="1062" points="320" swimtime="00:05:44.10" resultid="2377" heatid="2733" lane="5" />
                <RESULT eventid="1146" points="337" swimtime="00:02:42.07" resultid="2378" heatid="2829" lane="3" entrytime="00:02:44.04" entrycourse="LCM" />
                <RESULT eventid="1100" points="191" swimtime="00:01:36.23" resultid="2379" heatid="2775" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="292" swimtime="00:03:09.91" resultid="2380" heatid="2876" lane="7" entrytime="00:03:17.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                    <SPLIT distance="100" swimtime="00:01:34.23" />
                    <SPLIT distance="150" swimtime="00:02:29.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="De Ormeno" birthdate="2014-04-02" gender="M" nation="BRA" license="408702" athleteid="2452" externalid="408702">
              <RESULTS>
                <RESULT eventid="1167" points="153" reactiontime="+69" swimtime="00:00:43.94" resultid="2453" heatid="2855" lane="3" />
                <RESULT eventid="1125" points="189" swimtime="00:01:21.54" resultid="2454" heatid="2805" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="192" swimtime="00:00:36.20" resultid="2455" heatid="2889" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Ribeiro Melo" birthdate="2013-02-25" gender="M" nation="BRA" license="406921" swrid="5717293" athleteid="2427" externalid="406921">
              <RESULTS>
                <RESULT eventid="1077" points="111" swimtime="00:00:53.85" resultid="2428" heatid="2748" lane="5" />
                <RESULT eventid="1149" points="182" swimtime="00:02:59.97" resultid="2429" heatid="2830" lane="4" />
                <RESULT eventid="1135" points="193" swimtime="00:01:20.96" resultid="2430" heatid="2817" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="184" swimtime="00:00:36.74" resultid="2431" heatid="2900" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Bagatim" birthdate="2014-05-27" gender="F" nation="BRA" license="378353" swrid="5236649" athleteid="2331" externalid="378353">
              <RESULTS>
                <RESULT eventid="1080" points="221" swimtime="00:00:48.19" resultid="2332" heatid="2756" lane="5" entrytime="00:00:52.53" entrycourse="LCM" />
                <RESULT eventid="1106" points="238" swimtime="00:00:39.40" resultid="2333" heatid="2783" lane="4" entrytime="00:00:44.27" entrycourse="LCM" />
                <RESULT eventid="1122" points="230" swimtime="00:01:24.28" resultid="2334" heatid="2801" lane="3" entrytime="00:01:28.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="303" swimtime="00:00:35.12" resultid="2335" heatid="2886" lane="5" entrytime="00:00:37.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Zanatta Duda" birthdate="2013-08-28" gender="F" nation="BRA" license="406914" swrid="5717306" athleteid="2419" externalid="406914">
              <RESULTS>
                <RESULT eventid="1086" points="147" swimtime="00:01:48.45" resultid="2420" heatid="2764" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="141" swimtime="00:01:39.14" resultid="2421" heatid="2811" lane="5" />
                <RESULT eventid="1116" points="183" swimtime="00:00:47.26" resultid="2422" heatid="2788" lane="3" />
                <RESULT eventid="1208" points="166" swimtime="00:00:42.89" resultid="2423" heatid="2895" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dante" lastname="Gabriel Rossi" birthdate="2016-01-19" gender="M" nation="BRA" license="406928" swrid="5718627" athleteid="2445" externalid="406928">
              <RESULTS>
                <RESULT eventid="1130" points="50" swimtime="00:01:03.77" resultid="2446" heatid="2810" lane="3" />
                <RESULT eventid="1114" points="35" swimtime="00:01:07.92" resultid="2447" heatid="2787" lane="5" />
                <RESULT eventid="1216" points="51" swimtime="00:00:56.32" resultid="2448" heatid="2907" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Ognibeni Paupitz" birthdate="2014-08-08" gender="F" nation="BRA" license="406923" swrid="5718889" athleteid="2437" externalid="406923">
              <RESULTS>
                <RESULT eventid="1080" points="102" swimtime="00:01:02.31" resultid="2438" heatid="2754" lane="2" />
                <RESULT eventid="1202" points="128" swimtime="00:00:46.84" resultid="2439" heatid="2883" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robsson" lastname="Tows Oliveira" birthdate="2014-03-05" gender="M" nation="BRA" license="392107" swrid="5603922" athleteid="2394" externalid="392107">
              <RESULTS>
                <RESULT eventid="1083" points="158" swimtime="00:00:47.97" resultid="2395" heatid="2762" lane="3" entrytime="00:00:51.67" entrycourse="LCM" />
                <RESULT eventid="1167" points="111" swimtime="00:00:48.97" resultid="2396" heatid="2858" lane="6" entrytime="00:00:49.85" entrycourse="LCM" />
                <RESULT eventid="1125" points="138" swimtime="00:01:30.61" resultid="2397" heatid="2808" lane="2" entrytime="00:01:31.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="162" swimtime="00:00:38.33" resultid="2398" heatid="2892" lane="4" entrytime="00:00:40.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="De Andrade" birthdate="2015-12-24" gender="M" nation="BRA" license="406922" athleteid="2432" externalid="406922">
              <RESULTS>
                <RESULT eventid="1083" points="73" swimtime="00:01:02.01" resultid="2433" heatid="2758" lane="5" />
                <RESULT eventid="1167" points="80" reactiontime="+51" swimtime="00:00:54.51" resultid="2434" heatid="2855" lane="2" />
                <RESULT eventid="1125" points="90" swimtime="00:01:44.50" resultid="2435" heatid="2806" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="90" swimtime="00:00:46.55" resultid="2436" heatid="2890" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marco" lastname="Manzotti Marchi" birthdate="2015-06-26" gender="M" nation="BRA" license="396849" swrid="5641769" athleteid="2381" externalid="396849">
              <RESULTS>
                <RESULT eventid="1083" points="58" swimtime="00:01:06.92" resultid="2382" heatid="2758" lane="8" />
                <RESULT eventid="1109" points="52" swimtime="00:00:59.51" resultid="2383" heatid="2785" lane="5" entrytime="00:01:02.73" entrycourse="LCM" />
                <RESULT eventid="1205" points="83" swimtime="00:00:47.93" resultid="2384" heatid="2890" lane="3" entrytime="00:01:00.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Valentina Gozaga" birthdate="2014-06-28" gender="F" nation="BRA" license="385709" swrid="5603924" athleteid="2356" externalid="385709">
              <RESULTS>
                <RESULT eventid="1080" points="146" swimtime="00:00:55.33" resultid="2357" heatid="2755" lane="8" entrytime="00:01:09.40" entrycourse="LCM" />
                <RESULT eventid="1164" points="153" swimtime="00:00:50.21" resultid="2358" heatid="2852" lane="2" entrytime="00:00:51.94" entrycourse="LCM" />
                <RESULT eventid="1122" points="163" swimtime="00:01:34.64" resultid="2359" heatid="2801" lane="7" entrytime="00:01:41.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="220" swimtime="00:00:39.09" resultid="2360" heatid="2885" lane="4" entrytime="00:00:45.82" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benicio" lastname="Alves" birthdate="2012-04-26" gender="M" nation="BRA" license="370588" athleteid="2456" externalid="370588">
              <RESULTS>
                <RESULT eventid="1149" points="147" swimtime="00:03:13.01" resultid="2457" heatid="2831" lane="3" />
                <RESULT eventid="1135" points="152" swimtime="00:01:27.75" resultid="2458" heatid="2816" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="147" swimtime="00:00:44.57" resultid="2459" heatid="2793" lane="1" />
                <RESULT eventid="1211" points="185" swimtime="00:00:36.66" resultid="2460" heatid="2900" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Moreschi" birthdate="2012-08-09" gender="M" nation="BRA" license="385715" swrid="5603876" athleteid="2361" externalid="385715">
              <RESULTS>
                <RESULT eventid="1077" points="200" swimtime="00:00:44.32" resultid="2362" heatid="2751" lane="1" entrytime="00:00:45.64" entrycourse="LCM" />
                <RESULT eventid="1149" points="202" swimtime="00:02:53.79" resultid="2363" heatid="2831" lane="7" />
                <RESULT eventid="1173" points="191" swimtime="00:01:38.64" resultid="2364" heatid="2864" lane="6" entrytime="00:01:41.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="220" swimtime="00:03:08.80" resultid="2365" heatid="2879" lane="7" entrytime="00:03:20.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                    <SPLIT distance="100" swimtime="00:01:35.19" />
                    <SPLIT distance="150" swimtime="00:02:26.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Tiemi Yamaguchi" birthdate="2013-02-28" gender="F" nation="BRA" license="385707" swrid="5603920" athleteid="2351" externalid="385707">
              <RESULTS>
                <RESULT eventid="1074" points="246" swimtime="00:00:46.53" resultid="2352" heatid="2746" lane="1" entrytime="00:00:58.44" entrycourse="LCM" />
                <RESULT eventid="1158" points="248" swimtime="00:00:38.87" resultid="2353" heatid="2843" lane="6" entrytime="00:00:43.20" entrycourse="LCM" />
                <RESULT eventid="1100" points="223" swimtime="00:01:31.40" resultid="2354" heatid="2776" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="276" swimtime="00:03:13.48" resultid="2355" heatid="2876" lane="8" entrytime="00:03:37.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Rezende" birthdate="2012-01-23" gender="F" nation="BRA" license="370669" swrid="5603899" athleteid="2341" externalid="370669">
              <RESULTS>
                <RESULT eventid="1062" points="223" swimtime="00:06:28.10" resultid="2342" heatid="2733" lane="1" />
                <RESULT eventid="1074" points="169" swimtime="00:00:52.66" resultid="2343" heatid="2746" lane="2" entrytime="00:00:57.36" entrycourse="LCM" />
                <RESULT eventid="1146" points="227" swimtime="00:03:04.76" resultid="2344" heatid="2828" lane="5" entrytime="00:03:20.31" entrycourse="LCM" />
                <RESULT eventid="1170" points="175" swimtime="00:01:54.47" resultid="2345" heatid="2860" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Posser" birthdate="2013-02-07" gender="F" nation="BRA" license="378343" swrid="5603896" athleteid="2311" externalid="378343">
              <RESULTS>
                <RESULT eventid="1146" points="179" swimtime="00:03:20.02" resultid="2312" heatid="2828" lane="3" entrytime="00:03:40.21" entrycourse="LCM" />
                <RESULT eventid="1158" points="118" swimtime="00:00:49.77" resultid="2313" heatid="2841" lane="4" entrytime="00:00:56.24" entrycourse="LCM" />
                <RESULT eventid="1100" points="111" swimtime="00:01:55.22" resultid="2314" heatid="2775" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="213" swimtime="00:00:39.49" resultid="2315" heatid="2896" lane="7" entrytime="00:00:45.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Borges Duarte" birthdate="2014-02-10" gender="F" nation="BRA" license="408688" swrid="5725985" athleteid="2449" externalid="408688">
              <RESULTS>
                <RESULT eventid="1164" points="120" swimtime="00:00:54.40" resultid="2450" heatid="2850" lane="6" />
                <RESULT eventid="1202" points="138" swimtime="00:00:45.67" resultid="2451" heatid="2883" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Drapzichinski" birthdate="2015-08-21" gender="M" nation="BRA" license="391848" swrid="5603890" athleteid="2371" externalid="391848">
              <RESULTS>
                <RESULT eventid="1083" points="104" swimtime="00:00:55.12" resultid="2372" heatid="2760" lane="3" entrytime="00:01:09.84" entrycourse="LCM" />
                <RESULT eventid="1167" points="121" swimtime="00:00:47.49" resultid="2373" heatid="2856" lane="6" entrytime="00:01:08.17" entrycourse="LCM" />
                <RESULT eventid="1125" points="97" swimtime="00:01:41.68" resultid="2374" heatid="2805" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="118" swimtime="00:00:42.55" resultid="2375" heatid="2890" lane="5" entrytime="00:00:53.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monique" lastname="Istake" birthdate="2012-04-03" gender="F" nation="BRA" license="372023" swrid="5603857" athleteid="2336" externalid="372023">
              <RESULTS>
                <RESULT eventid="1146" points="302" swimtime="00:02:48.06" resultid="2337" heatid="2829" lane="2" entrytime="00:02:58.30" entrycourse="LCM" />
                <RESULT eventid="1158" points="258" swimtime="00:00:38.34" resultid="2338" heatid="2843" lane="5" entrytime="00:00:38.84" entrycourse="LCM" />
                <RESULT eventid="1132" points="298" swimtime="00:01:17.37" resultid="2339" heatid="2814" lane="4" entrytime="00:01:22.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="232" swimtime="00:01:30.19" resultid="2340" heatid="2777" lane="6" entrytime="00:01:39.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Paes Schemiko" birthdate="2013-02-25" gender="F" nation="BRA" license="406918" swrid="5725995" athleteid="2424" externalid="406918">
              <RESULTS>
                <RESULT eventid="1158" points="193" swimtime="00:00:42.23" resultid="2425" heatid="2840" lane="4" />
                <RESULT eventid="1208" points="258" swimtime="00:00:37.06" resultid="2426" heatid="2894" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Rossi" birthdate="2012-05-21" gender="M" nation="BRA" license="378346" swrid="5603901" athleteid="2316" externalid="378346">
              <RESULTS>
                <RESULT eventid="1089" points="212" swimtime="00:01:26.49" resultid="2317" heatid="2768" lane="2" entrytime="00:01:31.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="258" swimtime="00:01:13.54" resultid="2318" heatid="2820" lane="5" entrytime="00:01:17.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="239" swimtime="00:00:37.92" resultid="2319" heatid="2795" lane="3" entrytime="00:00:43.07" entrycourse="LCM" />
                <RESULT eventid="1211" points="286" swimtime="00:00:31.72" resultid="2320" heatid="2904" lane="6" entrytime="00:00:34.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Jupi Takaki" birthdate="2013-03-26" gender="F" nation="BRA" license="391845" swrid="5603861" athleteid="2366" externalid="391845">
              <RESULTS>
                <RESULT eventid="1062" points="224" swimtime="00:06:27.05" resultid="2367" heatid="2734" lane="1" />
                <RESULT eventid="1158" points="240" swimtime="00:00:39.29" resultid="2368" heatid="2842" lane="7" entrytime="00:00:51.75" entrycourse="LCM" />
                <RESULT eventid="1100" points="168" swimtime="00:01:40.36" resultid="2369" heatid="2776" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="202" swimtime="00:03:34.85" resultid="2370" heatid="2875" lane="1" entrytime="00:04:23.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.46" />
                    <SPLIT distance="100" swimtime="00:01:42.16" />
                    <SPLIT distance="150" swimtime="00:02:47.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Souza" birthdate="2013-09-11" gender="M" nation="BRA" license="382211" swrid="5603916" athleteid="2404" externalid="382211">
              <RESULTS>
                <RESULT eventid="1149" points="183" swimtime="00:02:59.45" resultid="2405" heatid="2832" lane="7" entrytime="00:03:04.07" entrycourse="LCM" />
                <RESULT eventid="1161" points="127" swimtime="00:00:44.25" resultid="2406" heatid="2846" lane="8" entrytime="00:00:47.24" entrycourse="LCM" />
                <RESULT eventid="1135" points="193" swimtime="00:01:21.01" resultid="2407" heatid="2819" lane="4" entrytime="00:01:23.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="163" swimtime="00:03:28.41" resultid="2408" heatid="2877" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.61" />
                    <SPLIT distance="100" swimtime="00:01:37.56" />
                    <SPLIT distance="150" swimtime="00:02:45.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Schmeiske Ruivo" birthdate="2013-10-21" gender="F" nation="BRA" license="402006" swrid="5661354" athleteid="2385" externalid="402006">
              <RESULTS>
                <RESULT eventid="1074" points="253" swimtime="00:00:46.09" resultid="2386" heatid="2744" lane="3" />
                <RESULT eventid="1132" points="196" swimtime="00:01:28.90" resultid="2387" heatid="2812" lane="3" entrytime="00:01:43.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="273" swimtime="00:00:41.36" resultid="2388" heatid="2790" lane="2" entrytime="00:00:48.91" entrycourse="LCM" />
                <RESULT eventid="1208" points="287" swimtime="00:00:35.76" resultid="2389" heatid="2896" lane="2" entrytime="00:00:44.82" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="9" agemin="9" agetotalmax="-1" agetotalmin="-1" gender="M" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1180" points="103" swimtime="00:03:00.95" resultid="2467" heatid="2867" lane="6">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2390" number="1" />
                    <RELAYPOSITION athleteid="2381" number="2" />
                    <RELAYPOSITION athleteid="2371" number="3" />
                    <RELAYPOSITION athleteid="2432" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1222" points="76" swimtime="00:03:39.35" resultid="2470" heatid="2910" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.83" />
                    <SPLIT distance="100" swimtime="00:01:56.55" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2432" number="1" />
                    <RELAYPOSITION athleteid="2371" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2381" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2390" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="M" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1190" points="241" swimtime="00:02:16.38" resultid="2468" heatid="2873" lane="6" entrytime="00:02:11.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                    <SPLIT distance="150" swimtime="00:01:44.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2326" number="1" />
                    <RELAYPOSITION athleteid="2456" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2361" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2316" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1232" points="222" reactiontime="+65" swimtime="00:02:33.98" resultid="2469" heatid="2916" lane="2" entrytime="00:02:36.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                    <SPLIT distance="100" swimtime="00:01:23.10" />
                    <SPLIT distance="150" swimtime="00:01:58.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2316" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2361" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2326" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2456" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="F" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1178" points="185" swimtime="00:02:47.11" resultid="2461" heatid="2866" lane="5" entrytime="00:02:30.85">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.89" />
                    <SPLIT distance="150" swimtime="00:02:02.63" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2356" number="1" />
                    <RELAYPOSITION athleteid="2449" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2331" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2437" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1220" points="135" reactiontime="+78" swimtime="00:03:25.64" resultid="2465" heatid="2909" lane="3" entrytime="00:03:03.29">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.83" />
                    <SPLIT distance="100" swimtime="00:01:52.15" />
                    <SPLIT distance="150" swimtime="00:02:37.30" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2449" number="1" reactiontime="+78" />
                    <RELAYPOSITION athleteid="2356" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2331" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2437" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="F" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1184" points="293" swimtime="00:02:23.44" resultid="2462" heatid="2869" lane="6" entrytime="00:02:28.41">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.31" />
                    <SPLIT distance="150" swimtime="00:01:48.73" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2376" number="1" />
                    <RELAYPOSITION athleteid="2424" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2366" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2351" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1226" points="301" reactiontime="+65" swimtime="00:02:37.44" resultid="2464" heatid="2912" lane="3" entrytime="00:02:43.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.21" />
                    <SPLIT distance="100" swimtime="00:01:24.76" />
                    <SPLIT distance="150" swimtime="00:02:03.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2385" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2351" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2366" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2376" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="F" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1186" points="337" swimtime="00:02:16.98" resultid="2463" heatid="2870" lane="3" entrytime="00:02:24.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                    <SPLIT distance="150" swimtime="00:01:41.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2321" number="1" />
                    <RELAYPOSITION athleteid="2336" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2306" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2414" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1228" points="314" reactiontime="+70" swimtime="00:02:35.28" resultid="2466" heatid="2913" lane="3" entrytime="00:02:49.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.84" />
                    <SPLIT distance="100" swimtime="00:01:23.41" />
                    <SPLIT distance="150" swimtime="00:02:00.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2414" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="2321" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2336" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2306" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="F" name="FÁBRICA DE NADADORES &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1184" status="DSQ" swimtime="00:02:29.93" resultid="2477" heatid="2869" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2419" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2385" number="2" reactiontime="+3276" status="DSQ" />
                    <RELAYPOSITION athleteid="2301" number="3" reactiontime="+3276" status="DSQ" />
                    <RELAYPOSITION athleteid="2346" number="4" reactiontime="+3276" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1226" points="184" reactiontime="+68" swimtime="00:03:05.57" resultid="2478" heatid="2912" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.84" />
                    <SPLIT distance="100" swimtime="00:01:39.38" />
                    <SPLIT distance="150" swimtime="00:02:23.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2346" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="2301" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2424" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2419" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="X" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1096" status="DSQ" swimtime="00:02:24.32" resultid="2471" heatid="2772" lane="6" entrytime="00:02:17.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                    <SPLIT distance="150" swimtime="00:01:49.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2427" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2404" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="2351" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="2376" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1142" swimtime="00:02:59.60" resultid="2476" heatid="2825" lane="6" entrytime="00:02:35.14">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2427" number="1" />
                    <RELAYPOSITION athleteid="2404" number="2" />
                    <RELAYPOSITION athleteid="2351" number="3" />
                    <RELAYPOSITION athleteid="2376" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="X" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1098" swimtime="00:02:08.65" resultid="2472" heatid="2774" lane="2" entrytime="00:02:13.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:04.47" />
                    <SPLIT distance="150" swimtime="00:01:35.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2321" number="1" />
                    <RELAYPOSITION athleteid="2336" number="2" />
                    <RELAYPOSITION athleteid="2316" number="3" />
                    <RELAYPOSITION athleteid="2326" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1144" swimtime="00:02:27.15" resultid="2474" heatid="2827" lane="7" entrytime="00:02:39.44">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2326" number="1" />
                    <RELAYPOSITION athleteid="2321" number="2" />
                    <RELAYPOSITION athleteid="2336" number="3" />
                    <RELAYPOSITION athleteid="2316" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="X" name="FÁBRICA DE NADADORES &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1094" swimtime="00:02:41.28" resultid="2473" heatid="2770" lane="3">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:05.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2356" number="1" />
                    <RELAYPOSITION athleteid="2394" number="2" />
                    <RELAYPOSITION athleteid="2440" number="3" />
                    <RELAYPOSITION athleteid="2331" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1140" swimtime="00:03:10.10" resultid="2475" heatid="2823" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2356" number="1" />
                    <RELAYPOSITION athleteid="2394" number="2" />
                    <RELAYPOSITION athleteid="2331" number="3" />
                    <RELAYPOSITION athleteid="2440" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="X" name="FÁBRICA DE NADADORES &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1098" swimtime="00:02:23.72" resultid="2479" heatid="2773" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:01:09.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2361" number="1" />
                    <RELAYPOSITION athleteid="2306" number="2" />
                    <RELAYPOSITION athleteid="2399" number="3" />
                    <RELAYPOSITION athleteid="2414" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1144" swimtime="00:02:42.24" resultid="2480" heatid="2826" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2399" number="1" />
                    <RELAYPOSITION athleteid="2306" number="2" />
                    <RELAYPOSITION athleteid="2414" number="3" />
                    <RELAYPOSITION athleteid="2361" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="11303" nation="BRA" region="PR" clubid="1446" swrid="93760" name="Associação De Talentos Da Natação" shortname="Atn/Curitiba">
          <ATHLETES>
            <ATHLETE firstname="Maximilian" lastname="Hock" birthdate="2016-11-20" gender="M" nation="DEU" license="408352" athleteid="1485" externalid="408352">
              <RESULTS>
                <RESULT eventid="1130" points="60" swimtime="00:01:00.03" resultid="1486" heatid="2810" lane="6" />
                <RESULT eventid="1216" points="77" swimtime="00:00:49.13" resultid="1487" heatid="2907" lane="3" />
                <RESULT eventid="1200" points="71" swimtime="00:01:02.48" resultid="1488" heatid="2881" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Goncalves Ghion" birthdate="2014-10-15" gender="F" nation="BRA" license="406912" swrid="5717269" athleteid="1480" externalid="406912">
              <RESULTS>
                <RESULT eventid="1080" points="113" swimtime="00:01:00.28" resultid="1481" heatid="2752" lane="5" />
                <RESULT eventid="1164" points="100" reactiontime="+61" swimtime="00:00:57.84" resultid="1482" heatid="2850" lane="2" />
                <RESULT eventid="1122" points="110" swimtime="00:01:47.71" resultid="1483" heatid="2800" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="126" swimtime="00:00:47.02" resultid="1484" heatid="2884" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Lemes Luis" birthdate="2013-10-14" gender="M" nation="BRA" license="410105" athleteid="1489" externalid="410105">
              <RESULTS>
                <RESULT eventid="1161" status="DNS" swimtime="00:00:00.00" resultid="1490" heatid="2844" lane="5" />
                <RESULT eventid="1135" points="135" swimtime="00:01:31.33" resultid="1491" heatid="2817" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="122" swimtime="00:00:47.37" resultid="1492" heatid="2792" lane="5" />
                <RESULT eventid="1211" points="147" swimtime="00:00:39.54" resultid="1493" heatid="2901" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Duarte De Almeida" birthdate="2013-12-09" gender="M" nation="BRA" license="385711" swrid="5588666" athleteid="1457" externalid="385711">
              <RESULTS>
                <RESULT eventid="1077" points="179" swimtime="00:00:45.96" resultid="1458" heatid="2748" lane="3" />
                <RESULT eventid="1161" points="213" swimtime="00:00:37.28" resultid="1459" heatid="2846" lane="2" entrytime="00:00:42.54" entrycourse="LCM" />
                <RESULT eventid="1211" points="258" swimtime="00:00:32.81" resultid="1460" heatid="2903" lane="5" entrytime="00:00:36.06" entrycourse="LCM" />
                <RESULT eventid="1195" status="DSQ" swimtime="00:03:08.05" resultid="1461" heatid="2878" lane="2" entrytime="00:03:26.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                    <SPLIT distance="100" swimtime="00:01:32.34" />
                    <SPLIT distance="150" swimtime="00:02:27.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Leal Kuss" birthdate="2012-10-20" gender="M" nation="BRA" license="385085" swrid="5588768" athleteid="1452" externalid="385085">
              <RESULTS>
                <RESULT eventid="1065" points="174" swimtime="00:06:33.68" resultid="1453" heatid="2736" lane="1" />
                <RESULT eventid="1161" points="232" swimtime="00:00:36.21" resultid="1454" heatid="2847" lane="2" entrytime="00:00:39.20" entrycourse="LCM" />
                <RESULT eventid="1103" points="169" swimtime="00:01:29.41" resultid="1455" heatid="2778" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="224" swimtime="00:00:34.42" resultid="1456" heatid="2903" lane="6" entrytime="00:00:36.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isis" lastname="De Miranda" birthdate="2012-01-10" gender="F" nation="BRA" license="397278" swrid="5652886" athleteid="1462" externalid="397278">
              <RESULTS>
                <RESULT eventid="1062" points="271" swimtime="00:06:03.34" resultid="1463" heatid="2734" lane="7" entrytime="00:06:18.97" entrycourse="LCM" />
                <RESULT eventid="1146" points="288" swimtime="00:02:50.71" resultid="1464" heatid="2829" lane="7" entrytime="00:03:00.52" entrycourse="LCM" />
                <RESULT eventid="1100" points="159" swimtime="00:01:42.30" resultid="1465" heatid="2777" lane="2" entrytime="00:01:52.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="308" swimtime="00:00:34.96" resultid="1466" heatid="2898" lane="1" entrytime="00:00:36.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Guedes Braga" birthdate="2013-04-09" gender="F" nation="BRA" license="385009" swrid="5602534" athleteid="1447" externalid="385009">
              <RESULTS>
                <RESULT eventid="1086" points="229" swimtime="00:01:33.67" resultid="1448" heatid="2764" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="269" swimtime="00:02:54.77" resultid="1449" heatid="2829" lane="1" entrytime="00:03:03.17" entrycourse="LCM" />
                <RESULT eventid="1132" points="328" swimtime="00:01:14.94" resultid="1450" heatid="2814" lane="5" entrytime="00:01:23.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="333" swimtime="00:00:34.05" resultid="1451" heatid="2898" lane="2" entrytime="00:00:36.22" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Vinicius Zonta" birthdate="2012-11-14" gender="M" nation="BRA" license="399517" swrid="5652903" athleteid="1467" externalid="399517">
              <RESULTS>
                <RESULT eventid="1149" points="258" swimtime="00:02:40.17" resultid="1468" heatid="2830" lane="5" />
                <RESULT eventid="1161" points="208" swimtime="00:00:37.58" resultid="1469" heatid="2844" lane="3" />
                <RESULT eventid="1135" points="282" swimtime="00:01:11.40" resultid="1470" heatid="2820" lane="3" entrytime="00:01:17.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="313" swimtime="00:00:30.79" resultid="1471" heatid="2904" lane="2" entrytime="00:00:34.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yohanna" lastname="Vitoria Sena" birthdate="2012-01-20" gender="F" nation="BRA" license="406710" swrid="5717302" athleteid="1472" externalid="406710">
              <RESULTS>
                <RESULT eventid="1132" points="128" swimtime="00:01:42.36" resultid="1473" heatid="2811" lane="7" />
                <RESULT eventid="1116" points="139" swimtime="00:00:51.74" resultid="1474" heatid="2789" lane="8" />
                <RESULT eventid="1208" points="170" swimtime="00:00:42.60" resultid="1475" heatid="2895" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Manuela Souza" birthdate="2016-07-07" gender="F" nation="BRA" license="406759" swrid="5717282" athleteid="1476" externalid="406759">
              <RESULTS>
                <RESULT eventid="1128" points="79" swimtime="00:01:02.34" resultid="1477" heatid="2809" lane="5" />
                <RESULT eventid="1214" points="83" swimtime="00:00:53.99" resultid="1478" heatid="2906" lane="6" />
                <RESULT eventid="1198" points="82" swimtime="00:01:06.88" resultid="1479" heatid="2880" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="M" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1190" points="236" swimtime="00:02:17.22" resultid="1494" heatid="2872" lane="4" entrytime="00:02:21.89">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                    <SPLIT distance="100" swimtime="00:01:13.97" />
                    <SPLIT distance="150" swimtime="00:01:43.60" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1489" number="1" />
                    <RELAYPOSITION athleteid="1467" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1457" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1452" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1232" points="185" reactiontime="+65" swimtime="00:02:43.62" resultid="1495" heatid="2915" lane="4" entrytime="00:02:52.19">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1489" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="1457" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1452" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1467" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="X" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1098" status="WDR" swimtime="00:00:00.00" resultid="1496" heatid="2774" lane="7" entrytime="00:02:16.46" />
                <RESULT eventid="1144" swimtime="00:02:54.00" resultid="1497" heatid="2827" lane="2" entrytime="00:02:38.19">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1472" number="1" />
                    <RELAYPOSITION athleteid="1467" number="2" />
                    <RELAYPOSITION athleteid="1462" number="3" />
                    <RELAYPOSITION athleteid="1452" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="13038" nation="BRA" region="PR" clubid="1400" swrid="93759" name="Associação De Pais E Atletas De Natação Ws/Crb" shortname="Apan/Ws">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Dos Santos" birthdate="2013-06-26" gender="F" nation="BRA" license="387512" swrid="5588662" athleteid="1411" externalid="387512">
              <RESULTS>
                <RESULT eventid="1086" points="199" swimtime="00:01:38.17" resultid="1412" heatid="2764" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="226" swimtime="00:03:05.03" resultid="1413" heatid="2828" lane="6" entrytime="00:03:49.81" entrycourse="LCM" />
                <RESULT eventid="1158" points="130" swimtime="00:00:48.13" resultid="1414" heatid="2841" lane="3" />
                <RESULT eventid="1116" points="222" swimtime="00:00:44.32" resultid="1415" heatid="2789" lane="3" entrytime="00:00:51.05" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leon" lastname="Bernardo Bello" birthdate="2014-11-23" gender="M" nation="BRA" license="400324" swrid="5717246" athleteid="1421" externalid="400324">
              <RESULTS>
                <RESULT eventid="1083" points="102" swimtime="00:00:55.43" resultid="1422" heatid="2760" lane="1" />
                <RESULT eventid="1167" points="115" reactiontime="+70" swimtime="00:00:48.42" resultid="1423" heatid="2854" lane="2" />
                <RESULT eventid="1125" points="113" swimtime="00:01:36.77" resultid="1424" heatid="2804" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="138" swimtime="00:00:40.45" resultid="1425" heatid="2890" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Bobko Ganacim" birthdate="2013-08-02" gender="F" nation="BRA" license="397332" swrid="5641754" athleteid="1406" externalid="397332">
              <RESULTS>
                <RESULT eventid="1074" status="DSQ" swimtime="00:01:02.11" resultid="1407" heatid="2745" lane="3" />
                <RESULT eventid="1132" points="131" swimtime="00:01:41.73" resultid="1408" heatid="2812" lane="2" entrytime="00:01:53.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="133" swimtime="00:00:52.49" resultid="1409" heatid="2789" lane="6" entrytime="00:00:54.06" entrycourse="LCM" />
                <RESULT eventid="1208" points="178" swimtime="00:00:41.95" resultid="1410" heatid="2896" lane="8" entrytime="00:00:48.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Gramms Dallarosa" birthdate="2015-01-14" gender="F" nation="BRA" license="406868" swrid="5717270" athleteid="1431" externalid="406868">
              <RESULTS>
                <RESULT eventid="1080" points="71" swimtime="00:01:10.36" resultid="1432" heatid="2752" lane="4" />
                <RESULT eventid="1164" points="101" reactiontime="+69" swimtime="00:00:57.61" resultid="1433" heatid="2849" lane="4" />
                <RESULT eventid="1122" points="106" swimtime="00:01:49.17" resultid="1434" heatid="2799" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="120" swimtime="00:00:47.79" resultid="1435" heatid="2882" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Da Reginalda" birthdate="2012-11-09" gender="M" nation="BRA" license="400275" swrid="5717253" athleteid="1416" externalid="400275">
              <RESULTS>
                <RESULT eventid="1065" points="203" swimtime="00:06:14.12" resultid="1417" heatid="2735" lane="4" />
                <RESULT eventid="1077" points="121" swimtime="00:00:52.43" resultid="1418" heatid="2749" lane="7" />
                <RESULT eventid="1135" points="215" swimtime="00:01:18.12" resultid="1419" heatid="2817" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="210" swimtime="00:00:35.15" resultid="1420" heatid="2901" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Cravcenco Marcondes" birthdate="2012-06-23" gender="F" nation="BRA" license="406866" swrid="5725987" athleteid="1426" externalid="406866">
              <RESULTS>
                <RESULT eventid="1074" points="164" swimtime="00:00:53.19" resultid="1427" heatid="2744" lane="5" />
                <RESULT eventid="1116" points="215" swimtime="00:00:44.79" resultid="1428" heatid="2788" lane="4" />
                <RESULT eventid="1170" points="156" swimtime="00:01:58.91" resultid="1429" heatid="2859" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="202" swimtime="00:00:40.20" resultid="1430" heatid="2895" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Ferreira" birthdate="2012-12-29" gender="F" nation="BRA" license="382235" swrid="5602538" athleteid="1401" externalid="382235">
              <RESULTS>
                <RESULT eventid="1158" points="205" swimtime="00:00:41.41" resultid="1402" heatid="2842" lane="5" entrytime="00:00:48.60" entrycourse="LCM" />
                <RESULT eventid="1132" points="274" swimtime="00:01:19.54" resultid="1403" heatid="2813" lane="4" entrytime="00:01:30.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="163" swimtime="00:01:41.46" resultid="1404" heatid="2777" lane="7" entrytime="00:01:53.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" status="DSQ" swimtime="00:00:35.55" resultid="1405" heatid="2897" lane="6" entrytime="00:00:40.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Bernardi Iurk" birthdate="2012-04-14" gender="M" nation="BRA" license="408687" swrid="5725984" athleteid="1441" externalid="408687">
              <RESULTS>
                <RESULT eventid="1077" points="108" swimtime="00:00:54.35" resultid="1442" heatid="2749" lane="1" />
                <RESULT eventid="1135" points="152" swimtime="00:01:27.74" resultid="1443" heatid="2816" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" status="DSQ" swimtime="00:01:58.21" resultid="1444" heatid="2863" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="165" swimtime="00:00:38.11" resultid="1445" heatid="2900" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Bernardi Iurk" birthdate="2012-04-14" gender="M" nation="BRA" license="406940" swrid="5717245" athleteid="1436" externalid="406940">
              <RESULTS>
                <RESULT eventid="1089" points="125" swimtime="00:01:43.04" resultid="1437" heatid="2766" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="151" swimtime="00:01:27.99" resultid="1438" heatid="2817" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="124" swimtime="00:00:47.12" resultid="1439" heatid="2793" lane="6" />
                <RESULT eventid="1211" points="167" swimtime="00:00:37.93" resultid="1440" heatid="2900" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1007" nation="BRA" region="PR" clubid="2529" swrid="93785" name="Santa Mônica Clube De Campo" shortname="Santa Mônica">
          <ATHLETES>
            <ATHLETE firstname="Davi" lastname="Luiz Cruz" birthdate="2012-10-13" gender="M" nation="BRA" license="393209" swrid="5616447" athleteid="2625" externalid="393209">
              <RESULTS>
                <RESULT eventid="1077" points="130" swimtime="00:00:51.13" resultid="2626" heatid="2748" lane="4" />
                <RESULT eventid="1161" points="125" swimtime="00:00:44.48" resultid="2627" heatid="2846" lane="3" entrytime="00:00:42.41" entrycourse="LCM" />
                <RESULT eventid="1103" points="88" swimtime="00:01:51.10" resultid="2628" heatid="2779" lane="7" entrytime="00:01:48.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="122" swimtime="00:01:54.59" resultid="2629" heatid="2862" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tais" lastname="Feltrin Martins" birthdate="2013-01-17" gender="F" nation="BRA" license="406840" swrid="5717262" athleteid="2701" externalid="406840">
              <RESULTS>
                <RESULT eventid="1074" status="DSQ" swimtime="00:01:04.70" resultid="2702" heatid="2745" lane="8" />
                <RESULT eventid="1132" points="95" swimtime="00:01:53.17" resultid="2703" heatid="2811" lane="3" />
                <RESULT eventid="1116" points="85" swimtime="00:01:01.05" resultid="2704" heatid="2789" lane="1" />
                <RESULT eventid="1208" points="135" swimtime="00:00:46.02" resultid="2705" heatid="2895" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mathias" lastname="Bernardo" birthdate="2014-05-17" gender="M" nation="BRA" license="387376" swrid="5652880" athleteid="2595" externalid="387376">
              <RESULTS>
                <RESULT eventid="1071" points="138" swimtime="00:03:16.91" resultid="2596" heatid="2742" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.27" />
                    <SPLIT distance="150" swimtime="00:02:25.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="75" swimtime="00:01:01.30" resultid="2597" heatid="2758" lane="3" />
                <RESULT eventid="1125" points="139" swimtime="00:01:30.30" resultid="2598" heatid="2806" lane="5" entrytime="00:01:55.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="164" swimtime="00:00:38.12" resultid="2599" heatid="2890" lane="4" entrytime="00:00:52.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Wenceslau Bitencourt" birthdate="2012-02-11" gender="M" nation="BRA" license="377318" swrid="5602591" athleteid="2555" externalid="377318">
              <RESULTS>
                <RESULT eventid="1089" points="194" swimtime="00:01:29.08" resultid="2556" heatid="2767" lane="4" entrytime="00:01:39.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="208" swimtime="00:00:37.54" resultid="2557" heatid="2844" lane="2" />
                <RESULT eventid="1119" points="175" swimtime="00:00:42.03" resultid="2558" heatid="2794" lane="5" entrytime="00:00:46.32" entrycourse="LCM" />
                <RESULT eventid="1211" points="207" swimtime="00:00:35.30" resultid="2559" heatid="2903" lane="3" entrytime="00:00:36.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose" lastname="Vinicius Batistella" birthdate="2012-05-15" gender="M" nation="BRA" license="403785" swrid="5684613" athleteid="2692" externalid="403785">
              <RESULTS>
                <RESULT eventid="1149" points="147" swimtime="00:03:13.16" resultid="2693" heatid="2831" lane="4" entrytime="00:03:32.46" entrycourse="LCM" />
                <RESULT eventid="1135" points="163" swimtime="00:01:25.75" resultid="2694" heatid="2818" lane="4" entrytime="00:01:36.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="199" swimtime="00:00:35.79" resultid="2695" heatid="2902" lane="4" entrytime="00:00:39.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Prestes Alves Pinto" birthdate="2012-01-19" gender="F" nation="BRA" license="377324" swrid="5588867" athleteid="2560" externalid="377324">
              <RESULTS>
                <RESULT eventid="1086" points="298" swimtime="00:01:25.74" resultid="2561" heatid="2765" lane="2" entrytime="00:01:28.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="360" swimtime="00:01:12.65" resultid="2562" heatid="2815" lane="3" entrytime="00:01:13.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="306" swimtime="00:00:39.84" resultid="2563" heatid="2791" lane="2" entrytime="00:00:40.39" entrycourse="LCM" />
                <RESULT eventid="1192" points="305" swimtime="00:03:07.16" resultid="2564" heatid="2874" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.22" />
                    <SPLIT distance="100" swimtime="00:01:33.15" />
                    <SPLIT distance="150" swimtime="00:02:27.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Gabriel Broto" birthdate="2014-09-14" gender="M" nation="BRA" license="402171" swrid="5661345" athleteid="2670" externalid="402171">
              <RESULTS>
                <RESULT eventid="1125" status="DNS" swimtime="00:00:00.00" resultid="2671" heatid="2805" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Andrade Guarido" birthdate="2014-05-17" gender="M" nation="BRA" license="400031" swrid="5652873" athleteid="2655" externalid="400031">
              <RESULTS>
                <RESULT eventid="1071" points="139" swimtime="00:03:16.74" resultid="2656" heatid="2743" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                    <SPLIT distance="100" swimtime="00:01:31.98" />
                    <SPLIT distance="150" swimtime="00:02:25.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="110" swimtime="00:00:54.04" resultid="2657" heatid="2761" lane="4" entrytime="00:00:58.84" entrycourse="LCM" />
                <RESULT eventid="1125" points="129" swimtime="00:01:32.52" resultid="2658" heatid="2807" lane="5" entrytime="00:01:42.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="142" swimtime="00:00:40.07" resultid="2659" heatid="2892" lane="2" entrytime="00:00:43.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Victoria De Medeiros" birthdate="2014-08-14" gender="F" nation="BRA" license="403782" swrid="5684611" athleteid="2687" externalid="403782">
              <RESULTS>
                <RESULT eventid="1080" points="105" swimtime="00:01:01.71" resultid="2688" heatid="2754" lane="3" />
                <RESULT eventid="1106" points="86" swimtime="00:00:55.20" resultid="2689" heatid="2781" lane="5" />
                <RESULT eventid="1164" points="99" reactiontime="+31" swimtime="00:00:57.93" resultid="2690" heatid="2850" lane="4" entrytime="00:01:10.50" entrycourse="LCM" />
                <RESULT eventid="1202" points="121" swimtime="00:00:47.73" resultid="2691" heatid="2884" lane="3" entrytime="00:01:11.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Ryan Rosa" birthdate="2014-01-14" gender="M" nation="BRA" license="400032" swrid="5652898" athleteid="2660" externalid="400032">
              <RESULTS>
                <RESULT eventid="1083" points="104" swimtime="00:00:55.09" resultid="2661" heatid="2761" lane="8" entrytime="00:01:06.50" entrycourse="LCM" />
                <RESULT eventid="1167" points="102" swimtime="00:00:50.32" resultid="2662" heatid="2856" lane="4" entrytime="00:00:58.79" entrycourse="LCM" />
                <RESULT eventid="1125" points="79" swimtime="00:01:49.16" resultid="2663" heatid="2806" lane="6" entrytime="00:02:05.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="96" swimtime="00:00:45.60" resultid="2664" heatid="2891" lane="1" entrytime="00:00:51.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Aparecida Lourenço Alves" birthdate="2013-11-06" gender="F" nation="BRA" license="387374" swrid="5588530" athleteid="2585" externalid="387374">
              <RESULTS>
                <RESULT eventid="1086" status="DNS" swimtime="00:00:00.00" resultid="2586" heatid="2763" lane="7" />
                <RESULT eventid="1132" status="DNS" swimtime="00:00:00.00" resultid="2587" heatid="2813" lane="1" entrytime="00:01:39.44" entrycourse="LCM" />
                <RESULT eventid="1116" status="DNS" swimtime="00:00:00.00" resultid="2588" heatid="2790" lane="6" entrytime="00:00:48.90" entrycourse="LCM" />
                <RESULT eventid="1208" status="DNS" swimtime="00:00:00.00" resultid="2589" heatid="2896" lane="5" entrytime="00:00:43.03" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Luiza Rocha Batista" birthdate="2013-11-24" gender="F" nation="BRA" license="387379" swrid="5588784" athleteid="2605" externalid="387379">
              <RESULTS>
                <RESULT eventid="1158" points="123" swimtime="00:00:49.00" resultid="2606" heatid="2842" lane="8" entrytime="00:00:56.10" entrycourse="LCM" />
                <RESULT eventid="1132" points="220" swimtime="00:01:25.62" resultid="2607" heatid="2813" lane="8" entrytime="00:01:40.19" entrycourse="LCM" />
                <RESULT eventid="1100" points="132" swimtime="00:01:48.88" resultid="2608" heatid="2776" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="233" swimtime="00:00:38.32" resultid="2609" heatid="2896" lane="3" entrytime="00:00:43.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lais" lastname="Manika Broto" birthdate="2013-03-27" gender="F" nation="BRA" license="378054" swrid="5588795" athleteid="2565" externalid="378054">
              <RESULTS>
                <RESULT eventid="1062" points="346" swimtime="00:05:34.99" resultid="2566" heatid="2733" lane="7" />
                <RESULT eventid="1158" points="298" swimtime="00:00:36.56" resultid="2567" heatid="2842" lane="3" entrytime="00:00:49.40" entrycourse="LCM" />
                <RESULT eventid="1132" points="378" swimtime="00:01:11.50" resultid="2568" heatid="2815" lane="7" entrytime="00:01:20.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="319" swimtime="00:03:04.45" resultid="2569" heatid="2875" lane="3" entrytime="00:03:42.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="100" swimtime="00:01:28.18" />
                    <SPLIT distance="150" swimtime="00:02:24.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mathias" lastname="Lopes Batista" birthdate="2012-08-22" gender="M" nation="BRA" license="399740" swrid="5652889" athleteid="2650" externalid="399740">
              <RESULTS>
                <RESULT eventid="1089" points="181" swimtime="00:01:31.14" resultid="2651" heatid="2768" lane="8" entrytime="00:01:38.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="180" swimtime="00:01:22.97" resultid="2652" heatid="2819" lane="1" entrytime="00:01:35.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="177" swimtime="00:00:41.88" resultid="2653" heatid="2795" lane="7" entrytime="00:00:44.29" entrycourse="LCM" />
                <RESULT eventid="1211" points="176" swimtime="00:00:37.30" resultid="2654" heatid="2903" lane="8" entrytime="00:00:39.22" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Zanotto De Souza" birthdate="2013-08-24" gender="M" nation="BRA" license="388361" swrid="5588974" athleteid="2615" externalid="388361">
              <RESULTS>
                <RESULT eventid="1065" points="260" swimtime="00:05:44.41" resultid="2616" heatid="2736" lane="7" />
                <RESULT eventid="1149" points="226" swimtime="00:02:47.23" resultid="2617" heatid="2833" lane="1" entrytime="00:02:51.35" entrycourse="LCM" />
                <RESULT eventid="1135" points="235" swimtime="00:01:15.91" resultid="2618" heatid="2820" lane="7" entrytime="00:01:20.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="206" swimtime="00:03:12.87" resultid="2619" heatid="2878" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lis" lastname="Cristini Harmatiuk" birthdate="2014-07-19" gender="F" nation="BRA" license="396830" swrid="5641759" athleteid="2696" externalid="396830">
              <RESULTS>
                <RESULT eventid="1068" points="167" swimtime="00:03:24.68" resultid="2697" heatid="2738" lane="2" />
                <RESULT eventid="1080" points="162" swimtime="00:00:53.47" resultid="2698" heatid="2756" lane="6" entrytime="00:00:54.41" entrycourse="LCM" />
                <RESULT eventid="1164" points="175" swimtime="00:00:48.00" resultid="2699" heatid="2852" lane="3" entrytime="00:00:50.46" entrycourse="LCM" />
                <RESULT eventid="1202" points="188" swimtime="00:00:41.18" resultid="2700" heatid="2886" lane="8" entrytime="00:00:44.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="De Siqueira Machado" birthdate="2012-05-25" gender="F" nation="BRA" license="377312" swrid="5588649" athleteid="2535" externalid="377312">
              <RESULTS>
                <RESULT eventid="1074" points="272" swimtime="00:00:44.97" resultid="2536" heatid="2745" lane="6" />
                <RESULT eventid="1158" points="191" swimtime="00:00:42.37" resultid="2537" heatid="2843" lane="1" entrytime="00:00:45.99" entrycourse="LCM" />
                <RESULT eventid="1116" points="284" swimtime="00:00:40.85" resultid="2538" heatid="2791" lane="7" entrytime="00:00:42.21" entrycourse="LCM" />
                <RESULT eventid="1208" points="390" swimtime="00:00:32.29" resultid="2539" heatid="2899" lane="2" entrytime="00:00:34.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Fachini Kovalski" birthdate="2012-05-15" gender="M" nation="BRA" license="403404" swrid="5676297" athleteid="2682" externalid="403404">
              <RESULTS>
                <RESULT eventid="1089" points="116" swimtime="00:01:45.70" resultid="2683" heatid="2766" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="91" swimtime="00:01:44.00" resultid="2684" heatid="2818" lane="3" entrytime="00:01:38.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="103" swimtime="00:00:50.08" resultid="2685" heatid="2794" lane="2" entrytime="00:00:50.71" entrycourse="LCM" />
                <RESULT eventid="1211" points="124" swimtime="00:00:41.87" resultid="2686" heatid="2902" lane="2" entrytime="00:00:43.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helenna" lastname="Banzatto Silva" birthdate="2013-07-11" gender="F" nation="BRA" license="393210" swrid="5616439" athleteid="2630" externalid="393210">
              <RESULTS>
                <RESULT eventid="1074" points="144" swimtime="00:00:55.62" resultid="2631" heatid="2745" lane="4" entrytime="00:01:04.76" entrycourse="LCM" />
                <RESULT eventid="1116" points="70" swimtime="00:01:05.14" resultid="2632" heatid="2789" lane="2" entrytime="00:01:15.04" entrycourse="LCM" />
                <RESULT eventid="1170" points="148" swimtime="00:02:01.09" resultid="2633" heatid="2859" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="78" swimtime="00:00:55.25" resultid="2634" heatid="2895" lane="3" entrytime="00:01:19.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Camily Moraes" birthdate="2014-07-13" gender="F" nation="BRA" license="397159" swrid="5641755" athleteid="2640" externalid="397159">
              <RESULTS>
                <RESULT eventid="1068" points="153" swimtime="00:03:30.55" resultid="2641" heatid="2740" lane="1" entrytime="00:04:07.93" entrycourse="LCM" />
                <RESULT eventid="1164" points="169" reactiontime="+59" swimtime="00:00:48.54" resultid="2642" heatid="2852" lane="7" entrytime="00:00:52.04" entrycourse="LCM" />
                <RESULT eventid="1122" points="147" swimtime="00:01:37.93" resultid="2643" heatid="2800" lane="6" entrytime="00:01:56.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="179" swimtime="00:00:41.86" resultid="2644" heatid="2885" lane="6" entrytime="00:00:47.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauren" lastname="Kurecki" birthdate="2014-03-06" gender="F" nation="BRA" license="377314" swrid="5602549" athleteid="2540" externalid="377314">
              <RESULTS>
                <RESULT eventid="1068" points="280" swimtime="00:02:52.42" resultid="2541" heatid="2740" lane="4" entrytime="00:02:58.56" entrycourse="LCM" />
                <RESULT eventid="1080" points="278" swimtime="00:00:44.66" resultid="2542" heatid="2756" lane="4" entrytime="00:00:47.71" entrycourse="LCM" />
                <RESULT eventid="1122" points="289" swimtime="00:01:18.18" resultid="2543" heatid="2801" lane="4" entrytime="00:01:21.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="346" swimtime="00:00:33.61" resultid="2544" heatid="2886" lane="4" entrytime="00:00:35.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Borges Piekarzievicz" birthdate="2013-09-10" gender="M" nation="BRA" license="403142" swrid="5676294" athleteid="2672" externalid="403142">
              <RESULTS>
                <RESULT eventid="1077" points="113" swimtime="00:00:53.58" resultid="2673" heatid="2749" lane="2" entrytime="00:01:02.75" entrycourse="LCM" />
                <RESULT eventid="1135" points="117" swimtime="00:01:35.74" resultid="2674" heatid="2817" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="101" swimtime="00:02:02.11" resultid="2675" heatid="2863" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="135" swimtime="00:00:40.71" resultid="2676" heatid="2901" lane="2" entrytime="00:00:49.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cleverson" lastname="Cardoso" birthdate="2013-07-20" gender="M" nation="BRA" license="387382" swrid="5588577" athleteid="2610" externalid="387382">
              <RESULTS>
                <RESULT eventid="1077" points="139" swimtime="00:00:50.01" resultid="2611" heatid="2749" lane="6" entrytime="00:00:57.67" entrycourse="LCM" />
                <RESULT eventid="1135" points="154" swimtime="00:01:27.27" resultid="2612" heatid="2818" lane="8" entrytime="00:01:48.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="111" swimtime="00:00:48.90" resultid="2613" heatid="2794" lane="8" entrytime="00:00:51.80" entrycourse="LCM" />
                <RESULT eventid="1211" points="142" swimtime="00:00:39.99" resultid="2614" heatid="2901" lane="6" entrytime="00:00:47.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Zattar" birthdate="2012-04-19" gender="F" nation="BRA" license="401736" swrid="5661351" athleteid="2665" externalid="401736">
              <RESULTS>
                <RESULT eventid="1086" points="239" swimtime="00:01:32.30" resultid="2666" heatid="2765" lane="7" entrytime="00:01:32.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="250" swimtime="00:00:46.25" resultid="2667" heatid="2744" lane="2" />
                <RESULT eventid="1116" points="336" swimtime="00:00:38.62" resultid="2668" heatid="2791" lane="3" entrytime="00:00:39.15" entrycourse="LCM" />
                <RESULT eventid="1208" points="370" swimtime="00:00:32.88" resultid="2669" heatid="2898" lane="5" entrytime="00:00:35.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="Cirilo Da Cunha" birthdate="2013-05-26" gender="F" nation="BRA" license="377316" swrid="5588595" athleteid="2545" externalid="377316">
              <RESULTS>
                <RESULT eventid="1146" points="293" swimtime="00:02:49.77" resultid="2546" heatid="2828" lane="1" />
                <RESULT eventid="1132" points="265" swimtime="00:01:20.49" resultid="2547" heatid="2813" lane="3" entrytime="00:01:32.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="218" swimtime="00:03:29.33" resultid="2548" heatid="2875" lane="2" entrytime="00:04:00.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.12" />
                    <SPLIT distance="100" swimtime="00:01:44.53" />
                    <SPLIT distance="150" swimtime="00:02:45.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="252" swimtime="00:00:37.35" resultid="2549" heatid="2896" lane="4" entrytime="00:00:42.96" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Rodrigues Bortoluzzi" birthdate="2013-10-07" gender="M" nation="BRA" license="387375" swrid="5652897" athleteid="2590" externalid="387375">
              <RESULTS>
                <RESULT eventid="1089" points="152" swimtime="00:01:36.63" resultid="2591" heatid="2767" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="158" swimtime="00:01:26.64" resultid="2592" heatid="2818" lane="5" entrytime="00:01:37.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="142" swimtime="00:00:45.11" resultid="2593" heatid="2794" lane="6" entrytime="00:00:47.75" entrycourse="LCM" />
                <RESULT eventid="1211" points="173" swimtime="00:00:37.50" resultid="2594" heatid="2902" lane="6" entrytime="00:00:40.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Lucachinski Villatore" birthdate="2013-10-04" gender="M" nation="BRA" license="382248" swrid="5588778" athleteid="2575" externalid="382248">
              <RESULTS>
                <RESULT eventid="1161" points="68" swimtime="00:00:54.30" resultid="2576" heatid="2845" lane="6" entrytime="00:01:00.58" entrycourse="LCM" />
                <RESULT eventid="1135" points="90" swimtime="00:01:44.39" resultid="2577" heatid="2818" lane="7" entrytime="00:01:46.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="94" swimtime="00:00:51.74" resultid="2578" heatid="2793" lane="5" entrytime="00:00:58.14" entrycourse="LCM" />
                <RESULT eventid="1211" points="115" swimtime="00:00:42.93" resultid="2579" heatid="2901" lane="5" entrytime="00:00:46.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Hugo Dos Santos" birthdate="2014-07-25" gender="M" nation="BRA" license="397420" swrid="5641766" athleteid="2645" externalid="397420">
              <RESULTS>
                <RESULT eventid="1083" points="78" swimtime="00:01:00.69" resultid="2646" heatid="2761" lane="1" entrytime="00:01:06.39" entrycourse="LCM" />
                <RESULT eventid="1155" points="91" swimtime="00:04:13.23" resultid="2647" heatid="2837" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.69" />
                    <SPLIT distance="100" swimtime="00:02:05.83" />
                    <SPLIT distance="150" swimtime="00:03:20.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="115" swimtime="00:01:36.32" resultid="2648" heatid="2807" lane="2" entrytime="00:01:46.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="120" swimtime="00:00:42.38" resultid="2649" heatid="2891" lane="3" entrytime="00:00:46.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Gouvea" birthdate="2013-04-19" gender="M" nation="BRA" license="387378" swrid="5588729" athleteid="2600" externalid="387378">
              <RESULTS>
                <RESULT eventid="1077" points="148" swimtime="00:00:49.02" resultid="2601" heatid="2750" lane="1" entrytime="00:00:52.83" entrycourse="LCM" />
                <RESULT eventid="1135" points="182" swimtime="00:01:22.66" resultid="2602" heatid="2819" lane="8" entrytime="00:01:36.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="171" swimtime="00:01:42.34" resultid="2603" heatid="2863" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="214" swimtime="00:00:34.92" resultid="2604" heatid="2902" lane="3" entrytime="00:00:40.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Julia Rocha" birthdate="2014-02-10" gender="F" nation="BRA" license="397158" swrid="5641767" athleteid="2635" externalid="397158">
              <RESULTS>
                <RESULT eventid="1106" points="177" swimtime="00:00:43.44" resultid="2636" heatid="2782" lane="4" entrytime="00:01:00.85" entrycourse="LCM" />
                <RESULT eventid="1164" points="225" reactiontime="+34" swimtime="00:00:44.14" resultid="2637" heatid="2852" lane="4" entrytime="00:00:47.71" entrycourse="LCM" />
                <RESULT eventid="1122" points="210" swimtime="00:01:26.92" resultid="2638" heatid="2801" lane="6" entrytime="00:01:37.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="251" swimtime="00:00:37.41" resultid="2639" heatid="2886" lane="6" entrytime="00:00:41.36" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Hoffmann Zoschke" birthdate="2015-03-22" gender="M" nation="BRA" license="390917" swrid="5602547" athleteid="2620" externalid="390917">
              <RESULTS>
                <RESULT eventid="1071" points="178" swimtime="00:03:01.26" resultid="2621" heatid="2742" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="100" swimtime="00:01:29.57" />
                    <SPLIT distance="150" swimtime="00:02:18.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="147" swimtime="00:03:35.58" resultid="2622" heatid="2838" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.95" />
                    <SPLIT distance="100" swimtime="00:01:47.49" />
                    <SPLIT distance="150" swimtime="00:02:51.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="166" swimtime="00:01:25.11" resultid="2623" heatid="2804" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="173" swimtime="00:00:37.50" resultid="2624" heatid="2892" lane="6" entrytime="00:00:43.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Strapasson" birthdate="2012-03-01" gender="M" nation="BRA" license="371377" swrid="5602585" athleteid="2530" externalid="371377">
              <RESULTS>
                <RESULT eventid="1077" points="264" swimtime="00:00:40.42" resultid="2531" heatid="2751" lane="5" entrytime="00:00:40.34" entrycourse="LCM" />
                <RESULT eventid="1135" points="330" swimtime="00:01:07.75" resultid="2532" heatid="2821" lane="5" entrytime="00:01:10.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="257" swimtime="00:01:29.35" resultid="2533" heatid="2864" lane="5" entrytime="00:01:30.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="301" swimtime="00:00:31.18" resultid="2534" heatid="2905" lane="7" entrytime="00:00:32.57" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Prestes" birthdate="2014-01-16" gender="M" nation="BRA" license="382249" swrid="5602574" athleteid="2580" externalid="382249">
              <RESULTS>
                <RESULT eventid="1071" points="144" swimtime="00:03:14.39" resultid="2581" heatid="2743" lane="3" entrytime="00:03:16.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                    <SPLIT distance="100" swimtime="00:01:30.23" />
                    <SPLIT distance="150" swimtime="00:02:24.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="138" swimtime="00:00:50.15" resultid="2582" heatid="2762" lane="7" entrytime="00:00:54.94" entrycourse="LCM" />
                <RESULT eventid="1125" points="165" swimtime="00:01:25.37" resultid="2583" heatid="2808" lane="6" entrytime="00:01:29.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="182" swimtime="00:00:36.88" resultid="2584" heatid="2893" lane="3" entrytime="00:00:38.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helloisa" lastname="De Bassani" birthdate="2012-09-23" gender="F" nation="BRA" license="403403" swrid="5676296" athleteid="2677" externalid="403403">
              <RESULTS>
                <RESULT eventid="1074" points="122" swimtime="00:00:58.73" resultid="2678" heatid="2745" lane="5" entrytime="00:01:16.00" entrycourse="LCM" />
                <RESULT eventid="1116" points="126" swimtime="00:00:53.54" resultid="2679" heatid="2789" lane="7" />
                <RESULT eventid="1170" points="111" swimtime="00:02:13.09" resultid="2680" heatid="2859" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="172" swimtime="00:00:42.44" resultid="2681" heatid="2895" lane="5" entrytime="00:00:50.32" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Celli Schneider" birthdate="2013-02-04" gender="M" nation="BRA" license="377317" swrid="5588588" athleteid="2550" externalid="377317">
              <RESULTS>
                <RESULT eventid="1089" points="162" swimtime="00:01:34.62" resultid="2551" heatid="2766" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="177" swimtime="00:01:23.38" resultid="2552" heatid="2820" lane="8" entrytime="00:01:22.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="165" swimtime="00:00:42.89" resultid="2553" heatid="2795" lane="6" entrytime="00:00:44.00" entrycourse="LCM" />
                <RESULT eventid="1211" points="222" swimtime="00:00:34.50" resultid="2554" heatid="2903" lane="4" entrytime="00:00:35.87" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Marini" birthdate="2014-04-09" gender="M" nation="BRA" license="382247" swrid="5684582" athleteid="2570" externalid="382247">
              <RESULTS>
                <RESULT eventid="1083" points="73" swimtime="00:01:01.99" resultid="2571" heatid="2760" lane="5" entrytime="00:01:08.58" entrycourse="LCM" />
                <RESULT eventid="1167" points="114" reactiontime="+66" swimtime="00:00:48.54" resultid="2572" heatid="2858" lane="8" entrytime="00:00:50.80" entrycourse="LCM" />
                <RESULT eventid="1125" points="135" swimtime="00:01:31.13" resultid="2573" heatid="2808" lane="7" entrytime="00:01:33.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="137" swimtime="00:00:40.52" resultid="2574" heatid="2892" lane="1" entrytime="00:00:44.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1182" points="158" swimtime="00:02:36.99" resultid="2712" heatid="2868" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                    <SPLIT distance="100" swimtime="00:01:16.37" />
                    <SPLIT distance="150" swimtime="00:01:56.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2580" number="1" />
                    <RELAYPOSITION athleteid="2595" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2655" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2570" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1224" status="DSQ" swimtime="00:03:08.63" resultid="2716" heatid="2911" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.77" />
                    <SPLIT distance="150" swimtime="00:02:29.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2580" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2655" number="2" reactiontime="+3276" status="DSQ" />
                    <RELAYPOSITION athleteid="2570" number="3" reactiontime="+3276" status="DSQ" />
                    <RELAYPOSITION athleteid="2595" number="4" reactiontime="+3276" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1188" points="213" swimtime="00:02:22.02" resultid="2713" heatid="2871" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2550" number="1" />
                    <RELAYPOSITION athleteid="2600" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2590" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2615" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1230" points="171" reactiontime="+66" swimtime="00:02:47.85" resultid="2717" heatid="2914" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.21" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2550" number="1" reactiontime="+66" />
                    <RELAYPOSITION athleteid="2600" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2615" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2590" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1190" points="221" swimtime="00:02:20.28" resultid="2714" heatid="2872" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                    <SPLIT distance="100" swimtime="00:01:12.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2555" number="1" />
                    <RELAYPOSITION athleteid="2650" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2625" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2530" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1232" points="207" swimtime="00:02:37.58" resultid="2715" heatid="2915" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                    <SPLIT distance="100" swimtime="00:01:22.95" />
                    <SPLIT distance="150" swimtime="00:02:02.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2650" number="1" />
                    <RELAYPOSITION athleteid="2530" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2555" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2625" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1178" points="246" swimtime="00:02:32.14" resultid="2706" heatid="2866" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.17" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2635" number="1" />
                    <RELAYPOSITION athleteid="2640" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2696" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2540" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1220" points="220" reactiontime="+53" swimtime="00:02:54.71" resultid="2710" heatid="2909" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.16" />
                    <SPLIT distance="100" swimtime="00:01:30.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2640" number="1" reactiontime="+53" />
                    <RELAYPOSITION athleteid="2540" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2635" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2696" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1184" points="225" swimtime="00:02:36.60" resultid="2707" heatid="2869" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                    <SPLIT distance="100" swimtime="00:01:11.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2565" number="1" />
                    <RELAYPOSITION athleteid="2605" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2701" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2545" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1226" points="201" reactiontime="+107" swimtime="00:03:00.25" resultid="2709" heatid="2912" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.94" />
                    <SPLIT distance="100" swimtime="00:01:43.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2545" number="1" reactiontime="+107" />
                    <RELAYPOSITION athleteid="2630" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2565" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2605" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1186" points="311" swimtime="00:02:20.60" resultid="2708" heatid="2870" lane="6">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:01:47.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2535" number="1" />
                    <RELAYPOSITION athleteid="2665" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2677" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2560" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1228" points="261" reactiontime="+69" swimtime="00:02:45.23" resultid="2711" heatid="2913" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:23.50" />
                    <SPLIT distance="150" swimtime="00:02:04.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2665" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2535" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2560" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2677" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1096" swimtime="00:02:16.69" resultid="2718" heatid="2772" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.89" />
                    <SPLIT distance="150" swimtime="00:01:42.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2550" number="1" />
                    <RELAYPOSITION athleteid="2565" number="2" />
                    <RELAYPOSITION athleteid="2545" number="3" />
                    <RELAYPOSITION athleteid="2615" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1142" swimtime="00:02:53.35" resultid="2723" heatid="2825" lane="8">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2550" number="1" />
                    <RELAYPOSITION athleteid="2545" number="2" />
                    <RELAYPOSITION athleteid="2565" number="3" />
                    <RELAYPOSITION athleteid="2615" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1098" swimtime="00:02:11.85" resultid="2719" heatid="2773" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:08.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2555" number="1" />
                    <RELAYPOSITION athleteid="2535" number="2" />
                    <RELAYPOSITION athleteid="2560" number="3" />
                    <RELAYPOSITION athleteid="2530" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1144" swimtime="00:02:32.89" resultid="2721" heatid="2826" lane="5">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2665" number="1" />
                    <RELAYPOSITION athleteid="2530" number="2" />
                    <RELAYPOSITION athleteid="2555" number="3" />
                    <RELAYPOSITION athleteid="2560" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1094" swimtime="00:02:26.76" resultid="2720" heatid="2771" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                    <SPLIT distance="150" swimtime="00:01:52.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2580" number="1" />
                    <RELAYPOSITION athleteid="2570" number="2" />
                    <RELAYPOSITION athleteid="2635" number="3" />
                    <RELAYPOSITION athleteid="2540" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1140" status="DSQ" swimtime="00:03:20.51" resultid="2722" heatid="2823" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2640" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2696" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="2655" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="2595" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1096" swimtime="00:02:37.69" resultid="2724" heatid="2772" lane="7" entrytime="00:02:46.79">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2605" number="1" />
                    <RELAYPOSITION athleteid="2600" number="2" />
                    <RELAYPOSITION athleteid="2701" number="3" />
                    <RELAYPOSITION athleteid="2590" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1142" swimtime="00:03:16.53" resultid="2729" heatid="2825" lane="7" entrytime="00:03:24.48">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2701" number="1" />
                    <RELAYPOSITION athleteid="2600" number="2" />
                    <RELAYPOSITION athleteid="2605" number="3" />
                    <RELAYPOSITION athleteid="2590" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1098" swimtime="00:02:31.70" resultid="2725" heatid="2773" lane="4" entrytime="00:02:31.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="100" swimtime="00:01:14.62" />
                    <SPLIT distance="150" swimtime="00:01:47.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2625" number="1" />
                    <RELAYPOSITION athleteid="2650" number="2" />
                    <RELAYPOSITION athleteid="2665" number="3" />
                    <RELAYPOSITION athleteid="2677" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1144" swimtime="00:02:57.42" resultid="2727" heatid="2827" lane="1" entrytime="00:02:53.00">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2650" number="1" />
                    <RELAYPOSITION athleteid="2535" number="2" />
                    <RELAYPOSITION athleteid="2625" number="3" />
                    <RELAYPOSITION athleteid="2677" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1094" swimtime="00:02:45.17" resultid="2726" heatid="2771" lane="7" entrytime="00:02:44.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2696" number="1" />
                    <RELAYPOSITION athleteid="2655" number="2" />
                    <RELAYPOSITION athleteid="2595" number="3" />
                    <RELAYPOSITION athleteid="2640" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1140" swimtime="00:02:57.26" resultid="2728" heatid="2824" lane="7" entrytime="00:02:56.36">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2635" number="1" />
                    <RELAYPOSITION athleteid="2580" number="2" />
                    <RELAYPOSITION athleteid="2540" number="3" />
                    <RELAYPOSITION athleteid="2570" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1096" status="WDR" swimtime="00:00:00.00" resultid="2730" heatid="2772" lane="8" />
                <RESULT eventid="1142" status="WDR" swimtime="00:00:00.00" resultid="2731" heatid="2825" lane="1" />
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="13025" nation="BRA" region="PR" clubid="1498" swrid="93779" name="Instituto Desportos Aquáticos De Foz Do Iguaçu" shortname="Cataratas Natação">
          <ATHLETES>
            <ATHLETE firstname="Vitor" lastname="Riam Nagorski De Lima" birthdate="2014-04-26" gender="M" nation="BRA" license="407802" swrid="5721507" athleteid="1543" externalid="407802">
              <RESULTS>
                <RESULT eventid="1083" points="62" swimtime="00:01:05.44" resultid="1544" heatid="2757" lane="4" />
                <RESULT eventid="1167" points="37" reactiontime="+62" swimtime="00:01:10.48" resultid="1545" heatid="2856" lane="7" />
                <RESULT eventid="1125" points="68" swimtime="00:01:54.31" resultid="1546" heatid="2804" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="65" swimtime="00:00:51.95" resultid="1547" heatid="2889" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paula" lastname="Palma Fornarolli" birthdate="2013-08-07" gender="F" nation="BRA" license="411995" athleteid="1553" externalid="411995">
              <RESULTS>
                <RESULT eventid="1158" points="91" swimtime="00:00:54.26" resultid="1554" heatid="2840" lane="5" />
                <RESULT eventid="1132" points="166" swimtime="00:01:34.02" resultid="1555" heatid="2812" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="204" swimtime="00:00:45.58" resultid="1556" heatid="2788" lane="5" />
                <RESULT eventid="1208" points="250" swimtime="00:00:37.43" resultid="1557" heatid="2894" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="De Souza" birthdate="2014-03-30" gender="M" nation="BRA" license="407800" swrid="5721499" athleteid="1538" externalid="407800">
              <RESULTS>
                <RESULT eventid="1083" points="127" swimtime="00:00:51.59" resultid="1539" heatid="2758" lane="1" />
                <RESULT eventid="1167" points="66" reactiontime="+73" swimtime="00:00:58.23" resultid="1540" heatid="2856" lane="8" />
                <RESULT eventid="1125" points="88" swimtime="00:01:45.13" resultid="1541" heatid="2805" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="98" swimtime="00:00:45.35" resultid="1542" heatid="2887" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alessandro" lastname="Cazzola" birthdate="2014-09-15" gender="M" nation="PRY" license="390713" athleteid="1514" externalid="390713" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1083" points="186" swimtime="00:00:45.38" resultid="1515" heatid="2762" lane="5" entrytime="00:00:50.24" entrycourse="LCM" />
                <RESULT eventid="1155" points="157" swimtime="00:03:31.07" resultid="1516" heatid="2839" lane="6" entrytime="00:03:54.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.97" />
                    <SPLIT distance="100" swimtime="00:01:44.87" />
                    <SPLIT distance="150" swimtime="00:02:46.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="170" swimtime="00:01:24.56" resultid="1517" heatid="2808" lane="3" entrytime="00:01:28.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="208" swimtime="00:00:35.29" resultid="1518" heatid="2893" lane="1" entrytime="00:00:38.87" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaleo" lastname="Bruno Da Luz" birthdate="2014-03-11" gender="M" nation="BRA" license="406658" swrid="4740124" athleteid="1524" externalid="406658" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1167" points="49" reactiontime="+68" swimtime="00:01:03.99" resultid="1525" heatid="2856" lane="1" />
                <RESULT eventid="1125" points="68" swimtime="00:01:54.79" resultid="1526" heatid="2802" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="73" swimtime="00:00:49.82" resultid="1527" heatid="2888" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benjamin" lastname="Perius Goncalves De Lima" birthdate="2016-06-09" gender="M" nation="BRA" license="407798" swrid="5721506" athleteid="1533" externalid="407798">
              <RESULTS>
                <RESULT eventid="1130" points="74" swimtime="00:00:56.03" resultid="1534" heatid="2810" lane="4" />
                <RESULT eventid="1114" points="76" swimtime="00:00:52.48" resultid="1535" heatid="2787" lane="4" />
                <RESULT eventid="1216" points="99" swimtime="00:00:45.16" resultid="1536" heatid="2907" lane="1" />
                <RESULT eventid="1200" points="66" swimtime="00:01:04.07" resultid="1537" heatid="2881" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Roza" birthdate="2013-06-05" gender="M" nation="BRA" license="374412" swrid="5588949" athleteid="1499" externalid="374412" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1161" points="223" swimtime="00:00:36.67" resultid="1500" heatid="2847" lane="7" entrytime="00:00:40.09" entrycourse="LCM" />
                <RESULT eventid="1135" points="253" swimtime="00:01:14.09" resultid="1501" heatid="2820" lane="4" entrytime="00:01:16.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="165" swimtime="00:01:30.10" resultid="1502" heatid="2779" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="264" swimtime="00:00:32.59" resultid="1503" heatid="2905" lane="8" entrytime="00:00:32.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Ioris Souza" birthdate="2015-09-10" gender="F" nation="BRA" license="406693" swrid="5042791" athleteid="1528" externalid="406693" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1080" points="111" swimtime="00:01:00.64" resultid="1529" heatid="2753" lane="1" />
                <RESULT eventid="1164" points="132" reactiontime="+65" swimtime="00:00:52.72" resultid="1530" heatid="2848" lane="3" />
                <RESULT eventid="1122" points="92" swimtime="00:01:54.37" resultid="1531" heatid="2798" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="126" swimtime="00:00:47.06" resultid="1532" heatid="2884" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joshua" lastname="Davalos Gimenez" birthdate="2013-10-22" gender="M" nation="PRY" license="380598" athleteid="1509" externalid="380598" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1065" points="215" swimtime="00:06:06.80" resultid="1510" heatid="2735" lane="2" />
                <RESULT eventid="1077" points="181" swimtime="00:00:45.84" resultid="1511" heatid="2750" lane="4" entrytime="00:00:46.40" entrycourse="LCM" />
                <RESULT eventid="1149" points="206" swimtime="00:02:52.66" resultid="1512" heatid="2831" lane="6" />
                <RESULT eventid="1173" points="176" swimtime="00:01:41.49" resultid="1513" heatid="2862" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrieli" lastname="Brietzke Sbardelatti" birthdate="2014-07-14" gender="F" nation="BRA" license="400456" swrid="4379861" athleteid="1519" externalid="400456" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1068" points="195" swimtime="00:03:14.37" resultid="1520" heatid="2739" lane="3" />
                <RESULT eventid="1080" points="138" swimtime="00:00:56.34" resultid="1521" heatid="2753" lane="7" />
                <RESULT eventid="1122" points="169" swimtime="00:01:33.42" resultid="1522" heatid="2798" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="198" swimtime="00:00:40.44" resultid="1523" heatid="2883" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Marcio Peixoto" birthdate="2012-10-22" gender="M" nation="BRA" license="411994" athleteid="1548" externalid="411994">
              <RESULTS>
                <RESULT eventid="1077" status="DSQ" swimtime="00:01:18.87" resultid="1549" heatid="2749" lane="8" />
                <RESULT eventid="1135" status="DSQ" swimtime="00:01:38.31" resultid="1550" heatid="2817" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="91" swimtime="00:00:52.23" resultid="1551" heatid="2793" lane="2" />
                <RESULT eventid="1211" points="148" swimtime="00:00:39.45" resultid="1552" heatid="2900" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edward" lastname="Mikael De Lima" birthdate="2012-03-11" gender="M" nation="BRA" license="376445" swrid="5588816" athleteid="1504" externalid="376445" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1065" points="313" swimtime="00:05:24.10" resultid="1505" heatid="2736" lane="3" entrytime="00:05:35.04" entrycourse="LCM" />
                <RESULT eventid="1149" points="330" swimtime="00:02:27.60" resultid="1506" heatid="2833" lane="4" entrytime="00:02:26.06" entrycourse="LCM" />
                <RESULT eventid="1135" points="351" swimtime="00:01:06.40" resultid="1507" heatid="2817" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="241" swimtime="00:01:19.44" resultid="1508" heatid="2779" lane="3" entrytime="00:01:28.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="M" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1182" points="104" swimtime="00:03:00.48" resultid="1558" heatid="2868" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1514" number="1" />
                    <RELAYPOSITION athleteid="1524" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1538" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1543" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1224" points="82" reactiontime="+65" swimtime="00:03:34.09" resultid="1561" heatid="2911" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1543" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="1538" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1514" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1524" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="M" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1190" points="237" swimtime="00:02:17.10" resultid="1559" heatid="2872" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.85" />
                    <SPLIT distance="150" swimtime="00:01:39.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1504" number="1" />
                    <RELAYPOSITION athleteid="1509" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1499" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1548" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1232" points="200" reactiontime="+77" swimtime="00:02:39.26" resultid="1560" heatid="2915" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:20.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1504" number="1" reactiontime="+77" />
                    <RELAYPOSITION athleteid="1509" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1499" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1548" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="X" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1094" swimtime="00:02:45.63" resultid="1562" heatid="2770" lane="5">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:04.11" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1519" number="1" />
                    <RELAYPOSITION athleteid="1528" number="2" />
                    <RELAYPOSITION athleteid="1514" number="3" />
                    <RELAYPOSITION athleteid="1538" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1140" swimtime="00:03:19.76" resultid="1563" heatid="2823" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1514" number="1" />
                    <RELAYPOSITION athleteid="1528" number="2" />
                    <RELAYPOSITION athleteid="1519" number="3" />
                    <RELAYPOSITION athleteid="1538" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="263" nation="BRA" region="PR" clubid="1661" swrid="75436" name="Clube Curitibano" shortname="Curitibano">
          <ATHLETES>
            <ATHLETE firstname="Alice" lastname="Karam Barbosa Lima" birthdate="2012-12-11" gender="F" nation="BRA" license="376956" swrid="5588758" athleteid="1762" externalid="376956">
              <RESULTS>
                <RESULT eventid="1062" points="313" swimtime="00:05:46.58" resultid="1763" heatid="2734" lane="6" entrytime="00:05:51.90" entrycourse="LCM" />
                <RESULT eventid="1086" points="306" swimtime="00:01:25.05" resultid="1764" heatid="2765" lane="3" entrytime="00:01:25.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="329" swimtime="00:01:14.88" resultid="1765" heatid="2815" lane="2" entrytime="00:01:17.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="333" swimtime="00:00:38.73" resultid="1766" heatid="2791" lane="6" entrytime="00:00:39.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Albuquerque" birthdate="2012-08-17" gender="F" nation="BRA" license="369275" swrid="5602507" athleteid="1712" externalid="369275">
              <RESULTS>
                <RESULT eventid="1074" points="416" swimtime="00:00:39.04" resultid="1713" heatid="2747" lane="4" entrytime="00:00:40.03" entrycourse="LCM" />
                <RESULT eventid="1170" points="417" swimtime="00:01:25.83" resultid="1714" heatid="2861" lane="4" entrytime="00:01:26.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="307" swimtime="00:03:06.89" resultid="1715" heatid="2876" lane="6" entrytime="00:03:10.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                    <SPLIT distance="100" swimtime="00:01:36.15" />
                    <SPLIT distance="150" swimtime="00:02:23.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="359" swimtime="00:00:33.21" resultid="1716" heatid="2899" lane="6" entrytime="00:00:34.51" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Lazzarotti Matias" birthdate="2012-03-19" gender="F" nation="BRA" license="391026" swrid="5602552" athleteid="1981" externalid="391026">
              <RESULTS>
                <RESULT eventid="1086" points="369" swimtime="00:01:19.89" resultid="1982" heatid="2765" lane="6" entrytime="00:01:26.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="428" swimtime="00:00:35.63" resultid="1983" heatid="2791" lane="5" entrytime="00:00:38.94" entrycourse="LCM" />
                <RESULT eventid="1170" points="296" swimtime="00:01:36.16" resultid="1984" heatid="2861" lane="7" entrytime="00:01:43.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="404" swimtime="00:00:31.93" resultid="1985" heatid="2899" lane="3" entrytime="00:00:33.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Francia Soares" birthdate="2014-06-01" gender="F" nation="BRA" license="391011" swrid="5602540" athleteid="1931" externalid="391011">
              <RESULTS>
                <RESULT eventid="1068" points="140" swimtime="00:03:37.28" resultid="1932" heatid="2739" lane="1" />
                <RESULT eventid="1106" points="76" swimtime="00:00:57.44" resultid="1933" heatid="2781" lane="6" />
                <RESULT eventid="1122" points="136" swimtime="00:01:40.41" resultid="1934" heatid="2800" lane="5" entrytime="00:01:48.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="166" swimtime="00:00:42.89" resultid="1935" heatid="2885" lane="5" entrytime="00:00:46.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Trevisan De Paula" birthdate="2014-01-27" gender="M" nation="BRA" license="377152" swrid="5602568" athleteid="1881" externalid="377152">
              <RESULTS>
                <RESULT eventid="1071" points="204" swimtime="00:02:53.22" resultid="1882" heatid="2743" lane="4" entrytime="00:02:54.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                    <SPLIT distance="100" swimtime="00:01:22.10" />
                    <SPLIT distance="150" swimtime="00:02:08.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="180" swimtime="00:00:39.38" resultid="1883" heatid="2786" lane="4" entrytime="00:00:39.86" entrycourse="LCM" />
                <RESULT eventid="1125" points="204" swimtime="00:01:19.50" resultid="1884" heatid="2808" lane="4" entrytime="00:01:19.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="241" swimtime="00:00:33.59" resultid="1885" heatid="2893" lane="5" entrytime="00:00:36.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="De Macedo Martynychen" birthdate="2015-06-12" gender="F" nation="BRA" license="399681" swrid="5652885" athleteid="2076" externalid="399681">
              <RESULTS>
                <RESULT eventid="1068" points="87" swimtime="00:04:13.92" resultid="2077" heatid="2739" lane="2" />
                <RESULT eventid="1106" points="69" swimtime="00:00:59.53" resultid="2078" heatid="2781" lane="1" />
                <RESULT eventid="1164" points="80" reactiontime="+68" swimtime="00:01:02.12" resultid="2079" heatid="2851" lane="8" entrytime="00:01:08.76" entrycourse="LCM" />
                <RESULT eventid="1122" points="69" swimtime="00:02:05.97" resultid="2080" heatid="2797" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Jacob Brunetti" birthdate="2015-11-10" gender="M" nation="BRA" license="406837" swrid="5717274" athleteid="2151" externalid="406837">
              <RESULTS>
                <RESULT eventid="1083" points="32" swimtime="00:01:21.56" resultid="2152" heatid="2757" lane="2" />
                <RESULT eventid="1167" points="36" swimtime="00:01:10.95" resultid="2153" heatid="2854" lane="7" />
                <RESULT eventid="1125" points="29" swimtime="00:02:32.30" resultid="2154" heatid="2803" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="29" swimtime="00:01:07.43" resultid="2155" heatid="2889" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joana" lastname="Asinelli Casagrande" birthdate="2013-10-26" gender="F" nation="BRA" license="376970" swrid="5588536" athleteid="1796" externalid="376970">
              <RESULTS>
                <RESULT eventid="1086" points="269" swimtime="00:01:28.72" resultid="1797" heatid="2763" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="228" swimtime="00:00:39.97" resultid="1798" heatid="2843" lane="2" entrytime="00:00:43.83" entrycourse="LCM" />
                <RESULT eventid="1100" points="210" swimtime="00:01:33.30" resultid="1799" heatid="2777" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="272" swimtime="00:03:14.43" resultid="1800" heatid="2875" lane="5" entrytime="00:03:38.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:34.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Bittencourt Ribas" birthdate="2013-02-01" gender="F" nation="BRA" license="372682" swrid="5588555" athleteid="1752" externalid="372682">
              <RESULTS>
                <RESULT eventid="1086" points="296" swimtime="00:01:25.97" resultid="1753" heatid="2763" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="235" swimtime="00:00:39.54" resultid="1754" heatid="2843" lane="3" entrytime="00:00:43.19" entrycourse="LCM" />
                <RESULT eventid="1116" points="294" swimtime="00:00:40.35" resultid="1755" heatid="2791" lane="1" entrytime="00:00:42.55" entrycourse="LCM" />
                <RESULT eventid="1208" points="315" swimtime="00:00:34.68" resultid="1756" heatid="2898" lane="6" entrytime="00:00:36.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Vanzo Assumpcao" birthdate="2012-05-15" gender="M" nation="BRA" license="369258" swrid="5588942" athleteid="1662" externalid="369258">
              <RESULTS>
                <RESULT eventid="1089" points="275" swimtime="00:01:19.28" resultid="1663" heatid="2768" lane="4" entrytime="00:01:23.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="318" swimtime="00:00:32.62" resultid="1664" heatid="2847" lane="4" entrytime="00:00:34.77" entrycourse="LCM" />
                <RESULT eventid="1103" points="248" swimtime="00:01:18.67" resultid="1665" heatid="2779" lane="5" entrytime="00:01:22.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="262" swimtime="00:00:36.80" resultid="1666" heatid="2796" lane="4" entrytime="00:00:38.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Sieczkowski Pacheco" birthdate="2015-11-20" gender="F" nation="BRA" license="393261" swrid="5616450" athleteid="2021" externalid="393261">
              <RESULTS>
                <RESULT eventid="1068" points="111" swimtime="00:03:54.72" resultid="2022" heatid="2739" lane="6" />
                <RESULT eventid="1080" points="120" swimtime="00:00:58.97" resultid="2023" heatid="2755" lane="3" entrytime="00:01:03.04" entrycourse="LCM" />
                <RESULT eventid="1152" points="122" swimtime="00:04:13.61" resultid="2024" heatid="2834" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.04" />
                    <SPLIT distance="100" swimtime="00:02:03.25" />
                    <SPLIT distance="150" swimtime="00:03:15.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1106" points="75" swimtime="00:00:57.77" resultid="2025" heatid="2782" lane="3" entrytime="00:01:11.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Della Villa Yang" birthdate="2012-10-08" gender="F" nation="BRA" license="369276" swrid="5588653" athleteid="1717" externalid="369276">
              <RESULTS>
                <RESULT eventid="1062" points="431" swimtime="00:05:11.46" resultid="1718" heatid="2734" lane="4" entrytime="00:05:15.29" entrycourse="LCM" />
                <RESULT eventid="1158" points="288" swimtime="00:00:36.96" resultid="1719" heatid="2840" lane="3" />
                <RESULT eventid="1132" points="421" swimtime="00:01:08.95" resultid="1720" heatid="2815" lane="5" entrytime="00:01:09.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="356" swimtime="00:02:57.91" resultid="1721" heatid="2876" lane="5" entrytime="00:03:04.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                    <SPLIT distance="100" swimtime="00:01:26.98" />
                    <SPLIT distance="150" swimtime="00:02:21.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alan" lastname="Batista Grise" birthdate="2014-03-27" gender="M" nation="BRA" license="391007" swrid="5602513" athleteid="1921" externalid="391007">
              <RESULTS>
                <RESULT eventid="1083" points="79" swimtime="00:01:00.33" resultid="1922" heatid="2761" lane="7" entrytime="00:01:04.85" entrycourse="LCM" />
                <RESULT eventid="1167" points="73" swimtime="00:00:56.30" resultid="1923" heatid="2857" lane="8" entrytime="00:00:57.38" entrycourse="LCM" />
                <RESULT eventid="1125" points="84" swimtime="00:01:46.79" resultid="1924" heatid="2806" lane="3" entrytime="00:01:55.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="78" swimtime="00:00:48.74" resultid="1925" heatid="2891" lane="7" entrytime="00:00:51.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Xavier Jardim" birthdate="2012-01-23" gender="M" nation="BRA" license="369259" swrid="5641781" athleteid="1667" externalid="369259">
              <RESULTS>
                <RESULT eventid="1089" points="226" swimtime="00:01:24.67" resultid="1668" heatid="2768" lane="7" entrytime="00:01:32.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1149" points="266" swimtime="00:02:38.44" resultid="1669" heatid="2833" lane="7" entrytime="00:02:46.75" entrycourse="LCM" />
                <RESULT eventid="1135" points="291" swimtime="00:01:10.67" resultid="1670" heatid="2821" lane="8" entrytime="00:01:14.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="282" swimtime="00:00:31.86" resultid="1671" heatid="2905" lane="1" entrytime="00:00:32.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Garcia" birthdate="2015-10-26" gender="M" nation="BRA" license="406967" swrid="5717271" athleteid="2176" externalid="406967">
              <RESULTS>
                <RESULT eventid="1083" points="26" swimtime="00:01:27.24" resultid="2177" heatid="2757" lane="3" />
                <RESULT eventid="1167" points="51" swimtime="00:01:03.30" resultid="2178" heatid="2853" lane="3" />
                <RESULT eventid="1125" points="22" swimtime="00:02:47.23" resultid="2179" heatid="2805" lane="5" />
                <RESULT eventid="1205" points="28" swimtime="00:01:08.06" resultid="2180" heatid="2887" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luigi" lastname="Antoniuk Paganini" birthdate="2014-11-13" gender="M" nation="BRA" license="382127" swrid="5602509" athleteid="1906" externalid="382127">
              <RESULTS>
                <RESULT eventid="1083" points="105" swimtime="00:00:54.96" resultid="1907" heatid="2759" lane="3" />
                <RESULT eventid="1167" status="DNS" swimtime="00:00:00.00" resultid="1908" heatid="2858" lane="7" entrytime="00:00:50.05" entrycourse="LCM" />
                <RESULT eventid="1125" points="145" swimtime="00:01:29.15" resultid="1909" heatid="2808" lane="8" entrytime="00:01:39.60" entrycourse="LCM" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="1910" heatid="2892" lane="8" entrytime="00:00:44.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Szpak De Vasconcelos" birthdate="2012-06-29" gender="M" nation="BRA" license="369271" swrid="5588928" athleteid="1702" externalid="369271">
              <RESULTS>
                <RESULT eventid="1077" points="297" swimtime="00:00:38.88" resultid="1703" heatid="2751" lane="4" entrytime="00:00:38.61" entrycourse="LCM" />
                <RESULT eventid="1149" points="309" swimtime="00:02:30.80" resultid="1704" heatid="2833" lane="5" entrytime="00:02:32.39" entrycourse="LCM" />
                <RESULT eventid="1135" points="343" swimtime="00:01:06.90" resultid="1705" heatid="2821" lane="4" entrytime="00:01:09.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="283" swimtime="00:01:26.59" resultid="1706" heatid="2864" lane="4" entrytime="00:01:27.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Toscani Kim" birthdate="2013-02-15" gender="F" nation="BRA" license="372683" swrid="5588939" athleteid="1757" externalid="372683">
              <RESULTS>
                <RESULT eventid="1074" points="307" swimtime="00:00:43.19" resultid="1758" heatid="2747" lane="6" entrytime="00:00:45.87" entrycourse="LCM" />
                <RESULT eventid="1100" points="196" swimtime="00:01:35.36" resultid="1759" heatid="2776" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="296" swimtime="00:01:36.12" resultid="1760" heatid="2860" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="291" swimtime="00:03:10.19" resultid="1761" heatid="2876" lane="1" entrytime="00:03:21.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.40" />
                    <SPLIT distance="100" swimtime="00:01:36.36" />
                    <SPLIT distance="150" swimtime="00:02:26.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Poletto Abrahao" birthdate="2014-10-20" gender="M" nation="BRA" license="382128" swrid="5602571" athleteid="1911" externalid="382128">
              <RESULTS>
                <RESULT eventid="1083" points="165" swimtime="00:00:47.23" resultid="1912" heatid="2762" lane="4" entrytime="00:00:44.75" entrycourse="LCM" />
                <RESULT eventid="1155" points="157" swimtime="00:03:30.92" resultid="1913" heatid="2839" lane="4" entrytime="00:03:23.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.17" />
                    <SPLIT distance="100" swimtime="00:01:41.87" />
                    <SPLIT distance="150" swimtime="00:02:44.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="118" swimtime="00:00:45.29" resultid="1914" heatid="2786" lane="3" entrytime="00:00:45.17" entrycourse="LCM" />
                <RESULT eventid="1125" points="142" swimtime="00:01:29.71" resultid="1915" heatid="2804" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Vian" birthdate="2014-03-25" gender="F" nation="BRA" license="393919" swrid="5641779" athleteid="2046" externalid="393919">
              <RESULTS>
                <RESULT eventid="1106" points="113" swimtime="00:00:50.48" resultid="2047" heatid="2781" lane="3" />
                <RESULT eventid="1164" points="171" reactiontime="+76" swimtime="00:00:48.38" resultid="2048" heatid="2849" lane="7" />
                <RESULT eventid="1122" points="139" swimtime="00:01:39.69" resultid="2049" heatid="2798" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="187" swimtime="00:00:41.27" resultid="2050" heatid="2883" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Lauand Lorenci" birthdate="2013-03-06" gender="M" nation="BRA" license="376982" swrid="5588764" athleteid="1821" externalid="376982">
              <RESULTS>
                <RESULT eventid="1077" status="DSQ" swimtime="00:00:42.34" resultid="1822" heatid="2751" lane="2" entrytime="00:00:43.83" entrycourse="LCM" />
                <RESULT eventid="1161" points="175" swimtime="00:00:39.74" resultid="1823" heatid="2846" lane="4" entrytime="00:00:41.66" entrycourse="LCM" />
                <RESULT eventid="1173" status="DSQ" swimtime="00:01:34.88" resultid="1824" heatid="2863" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="214" swimtime="00:03:10.35" resultid="1825" heatid="2879" lane="2" entrytime="00:03:16.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.47" />
                    <SPLIT distance="100" swimtime="00:01:36.62" />
                    <SPLIT distance="150" swimtime="00:02:27.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Morais Shibata" birthdate="2014-02-09" gender="M" nation="BRA" license="391018" swrid="5602561" athleteid="1946" externalid="391018">
              <RESULTS>
                <RESULT eventid="1083" points="116" swimtime="00:00:53.07" resultid="1947" heatid="2761" lane="3" entrytime="00:01:01.41" entrycourse="LCM" />
                <RESULT eventid="1167" points="127" swimtime="00:00:46.77" resultid="1948" heatid="2857" lane="3" entrytime="00:00:54.42" entrycourse="LCM" />
                <RESULT eventid="1125" points="116" swimtime="00:01:35.96" resultid="1949" heatid="2807" lane="7" entrytime="00:01:46.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="127" swimtime="00:00:41.57" resultid="1950" heatid="2891" lane="2" entrytime="00:00:47.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Dolberth Alcantara" birthdate="2014-09-26" gender="F" nation="BRA" license="382124" swrid="5602532" athleteid="1896" externalid="382124">
              <RESULTS>
                <RESULT eventid="1080" points="108" swimtime="00:01:01.13" resultid="1897" heatid="2755" lane="2" entrytime="00:01:03.67" entrycourse="LCM" />
                <RESULT eventid="1152" points="149" swimtime="00:03:57.81" resultid="1898" heatid="2836" lane="7" entrytime="00:04:17.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.75" />
                    <SPLIT distance="100" swimtime="00:01:58.71" />
                    <SPLIT distance="150" swimtime="00:03:05.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1106" points="107" swimtime="00:00:51.41" resultid="1899" heatid="2783" lane="8" entrytime="00:01:00.18" entrycourse="LCM" />
                <RESULT eventid="1164" points="138" reactiontime="+75" swimtime="00:00:51.88" resultid="1900" heatid="2852" lane="8" entrytime="00:00:55.47" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="De Lima Cavalcanti" birthdate="2014-10-07" gender="M" nation="BRA" license="385884" swrid="5684550" athleteid="2091" externalid="385884">
              <RESULTS>
                <RESULT eventid="1071" points="174" swimtime="00:03:02.42" resultid="2092" heatid="2743" lane="5" entrytime="00:03:12.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.46" />
                    <SPLIT distance="100" swimtime="00:01:28.95" />
                    <SPLIT distance="150" swimtime="00:02:18.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="94" swimtime="00:00:48.94" resultid="2093" heatid="2784" lane="3" />
                <RESULT eventid="1167" points="160" reactiontime="+49" swimtime="00:00:43.37" resultid="2094" heatid="2858" lane="4" entrytime="00:00:43.07" entrycourse="LCM" />
                <RESULT eventid="1125" points="173" swimtime="00:01:24.01" resultid="2095" heatid="2808" lane="5" entrytime="00:01:26.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Petraglia" birthdate="2012-03-28" gender="M" nation="BRA" license="369282" swrid="5602569" athleteid="1742" externalid="369282">
              <RESULTS>
                <RESULT eventid="1065" points="260" swimtime="00:05:44.72" resultid="1743" heatid="2736" lane="6" entrytime="00:05:35.54" entrycourse="LCM" />
                <RESULT eventid="1077" points="187" swimtime="00:00:45.37" resultid="1744" heatid="2751" lane="7" entrytime="00:00:45.51" entrycourse="LCM" />
                <RESULT eventid="1119" points="222" swimtime="00:00:38.88" resultid="1745" heatid="2795" lane="4" entrytime="00:00:41.26" entrycourse="LCM" />
                <RESULT eventid="1173" points="187" swimtime="00:01:39.37" resultid="1746" heatid="2864" lane="2" entrytime="00:01:42.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Viera Correa" birthdate="2012-03-07" gender="M" nation="BRA" license="369269" swrid="5602590" athleteid="1692" externalid="369269">
              <RESULTS>
                <RESULT eventid="1065" points="291" swimtime="00:05:31.86" resultid="1693" heatid="2735" lane="5" />
                <RESULT eventid="1149" points="298" swimtime="00:02:32.63" resultid="1694" heatid="2833" lane="3" entrytime="00:02:37.92" entrycourse="LCM" />
                <RESULT eventid="1135" points="307" swimtime="00:01:09.41" resultid="1695" heatid="2821" lane="6" entrytime="00:01:10.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="293" swimtime="00:00:31.46" resultid="1696" heatid="2905" lane="5" entrytime="00:00:31.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enrico" lastname="Hallage Bianchini" birthdate="2014-02-27" gender="M" nation="BRA" license="397164" swrid="5661348" athleteid="2051" externalid="397164">
              <RESULTS>
                <RESULT eventid="1155" points="123" swimtime="00:03:49.10" resultid="2052" heatid="2837" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.68" />
                    <SPLIT distance="150" swimtime="00:02:58.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="102" swimtime="00:00:47.54" resultid="2053" heatid="2786" lane="8" entrytime="00:00:54.28" entrycourse="LCM" />
                <RESULT eventid="1167" points="127" reactiontime="+67" swimtime="00:00:46.80" resultid="2054" heatid="2858" lane="2" entrytime="00:00:49.95" entrycourse="LCM" />
                <RESULT eventid="1125" points="153" swimtime="00:01:27.47" resultid="2055" heatid="2807" lane="8" entrytime="00:01:50.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Antunes Luzzi" birthdate="2014-02-14" gender="M" nation="BRA" license="391019" swrid="5602510" athleteid="1951" externalid="391019">
              <RESULTS>
                <RESULT eventid="1083" points="73" swimtime="00:01:02.04" resultid="1952" heatid="2760" lane="6" entrytime="00:01:10.90" entrycourse="LCM" />
                <RESULT eventid="1167" points="63" swimtime="00:00:58.95" resultid="1953" heatid="2856" lane="3" entrytime="00:01:07.48" entrycourse="LCM" />
                <RESULT eventid="1125" points="67" swimtime="00:01:55.23" resultid="1954" heatid="2806" lane="2" entrytime="00:02:22.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="52" swimtime="00:00:55.78" resultid="1955" heatid="2890" lane="6" entrytime="00:01:08.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Afonso Fowler" birthdate="2014-01-22" gender="M" nation="BRA" license="393264" swrid="5661338" athleteid="2036" externalid="393264">
              <RESULTS>
                <RESULT eventid="1109" points="78" swimtime="00:00:52.07" resultid="2037" heatid="2784" lane="5" />
                <RESULT eventid="1167" points="110" swimtime="00:00:49.09" resultid="2038" heatid="2857" lane="7" entrytime="00:00:55.35" entrycourse="LCM" />
                <RESULT eventid="1125" points="112" swimtime="00:01:36.96" resultid="2039" heatid="2807" lane="6" entrytime="00:01:45.05" entrycourse="LCM" />
                <RESULT eventid="1205" points="169" swimtime="00:00:37.78" resultid="2040" heatid="2891" lane="4" entrytime="00:00:46.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Nishimura Ramina" birthdate="2013-11-25" gender="M" nation="BRA" license="376989" swrid="5588831" athleteid="1861" externalid="376989">
              <RESULTS>
                <RESULT eventid="1065" points="183" swimtime="00:06:27.00" resultid="1862" heatid="2735" lane="7" />
                <RESULT eventid="1149" points="159" swimtime="00:03:07.89" resultid="1863" heatid="2832" lane="8" entrytime="00:03:27.26" entrycourse="LCM" />
                <RESULT eventid="1119" points="125" swimtime="00:00:47.09" resultid="1864" heatid="2793" lane="3" />
                <RESULT eventid="1211" points="161" swimtime="00:00:38.38" resultid="1865" heatid="2902" lane="8" entrytime="00:00:43.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Guimaraes Mesquita" birthdate="2013-12-30" gender="F" nation="BRA" license="391027" swrid="5602544" athleteid="1986" externalid="391027">
              <RESULTS>
                <RESULT eventid="1074" points="156" swimtime="00:00:54.12" resultid="1987" heatid="2746" lane="7" entrytime="00:00:57.59" entrycourse="LCM" />
                <RESULT eventid="1132" points="183" swimtime="00:01:31.04" resultid="1988" heatid="2813" lane="2" entrytime="00:01:36.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="187" swimtime="00:01:51.97" resultid="1989" heatid="2860" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="173" swimtime="00:00:42.34" resultid="1990" heatid="2896" lane="6" entrytime="00:00:44.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Massimo" lastname="Puppi Cardoso" birthdate="2015-03-30" gender="M" nation="BRA" license="406742" swrid="5717290" athleteid="2106" externalid="406742">
              <RESULTS>
                <RESULT eventid="1083" points="87" swimtime="00:00:58.44" resultid="2107" heatid="2759" lane="4" />
                <RESULT eventid="1155" points="62" swimtime="00:04:46.93" resultid="2108" heatid="2838" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.13" />
                    <SPLIT distance="100" swimtime="00:02:24.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="62" reactiontime="+49" swimtime="00:00:59.33" resultid="2109" heatid="2853" lane="5" />
                <RESULT eventid="1125" points="50" swimtime="00:02:06.43" resultid="2110" heatid="2805" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Clara Prado Biscaia" birthdate="2013-10-24" gender="F" nation="BRA" license="391015" swrid="5602526" athleteid="1936" externalid="391015">
              <RESULTS>
                <RESULT eventid="1062" points="181" swimtime="00:06:55.94" resultid="1937" heatid="2733" lane="4" />
                <RESULT eventid="1158" points="171" swimtime="00:00:43.95" resultid="1938" heatid="2842" lane="6" entrytime="00:00:50.62" entrycourse="LCM" />
                <RESULT eventid="1100" points="154" swimtime="00:01:43.45" resultid="1939" heatid="2776" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="187" swimtime="00:03:40.35" resultid="1940" heatid="2875" lane="8" entrytime="00:04:27.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:48.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Hallage Papp" birthdate="2012-07-02" gender="M" nation="BRA" license="377042" swrid="5588736" athleteid="1846" externalid="377042">
              <RESULTS>
                <RESULT eventid="1077" status="DSQ" swimtime="00:00:51.39" resultid="1847" heatid="2749" lane="3" entrytime="00:00:54.37" entrycourse="LCM" />
                <RESULT eventid="1135" points="174" swimtime="00:01:23.78" resultid="1848" heatid="2819" lane="5" entrytime="00:01:28.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" status="DSQ" swimtime="00:01:55.88" resultid="1849" heatid="2863" lane="4" entrytime="00:01:59.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="211" swimtime="00:00:35.08" resultid="1850" heatid="2903" lane="7" entrytime="00:00:37.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gael" lastname="Stramandinoli Zanicotti" birthdate="2015-03-21" gender="M" nation="BRA" license="406954" swrid="5717298" athleteid="2161" externalid="406954">
              <RESULTS>
                <RESULT eventid="1083" points="28" swimtime="00:01:24.58" resultid="2162" heatid="2759" lane="1" />
                <RESULT eventid="1167" points="46" swimtime="00:01:05.59" resultid="2163" heatid="2855" lane="7" />
                <RESULT eventid="1125" points="40" swimtime="00:02:16.58" resultid="2164" heatid="2804" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="41" swimtime="00:01:00.21" resultid="2165" heatid="2887" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Toscani Kim" birthdate="2015-10-02" gender="F" nation="BRA" license="397276" swrid="5641778" athleteid="2066" externalid="397276">
              <RESULTS>
                <RESULT eventid="1068" points="141" swimtime="00:03:36.75" resultid="2067" heatid="2739" lane="8" />
                <RESULT eventid="1080" points="167" swimtime="00:00:52.94" resultid="2068" heatid="2755" lane="6" entrytime="00:01:03.29" entrycourse="LCM" />
                <RESULT eventid="1152" points="155" swimtime="00:03:54.54" resultid="2069" heatid="2835" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.68" />
                    <SPLIT distance="100" swimtime="00:01:55.38" />
                    <SPLIT distance="150" swimtime="00:02:59.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1106" points="89" swimtime="00:00:54.59" resultid="2070" heatid="2781" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Corte Flor" birthdate="2016-12-03" gender="M" nation="BRA" license="412013" athleteid="2207" externalid="412013">
              <RESULTS>
                <RESULT eventid="1130" points="38" swimtime="00:01:09.91" resultid="2208" heatid="2810" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Ruschka Druszcz" birthdate="2016-05-09" gender="F" nation="BRA" license="412025" athleteid="2220" externalid="412025">
              <RESULTS>
                <RESULT eventid="1128" points="85" swimtime="00:01:00.99" resultid="2221" heatid="2809" lane="3" />
                <RESULT eventid="1214" points="93" swimtime="00:00:52.02" resultid="2222" heatid="2906" lane="4" />
                <RESULT eventid="1198" points="85" swimtime="00:01:06.26" resultid="2223" heatid="2880" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elisa" lastname="Osternack Almeida" birthdate="2015-04-14" gender="F" nation="BRA" license="406747" swrid="5717286" athleteid="2121" externalid="406747">
              <RESULTS>
                <RESULT eventid="1080" points="113" swimtime="00:01:00.25" resultid="2122" heatid="2753" lane="6" />
                <RESULT eventid="1106" points="73" swimtime="00:00:58.23" resultid="2123" heatid="2780" lane="5" />
                <RESULT eventid="1164" points="109" reactiontime="+57" swimtime="00:00:56.15" resultid="2124" heatid="2849" lane="1" />
                <RESULT eventid="1122" points="85" swimtime="00:01:57.52" resultid="2125" heatid="2798" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Fernandes  Dos Reis" birthdate="2012-09-18" gender="M" nation="BRA" license="369279" swrid="5588696" athleteid="1732" externalid="369279">
              <RESULTS>
                <RESULT eventid="1161" points="251" swimtime="00:00:35.26" resultid="1733" heatid="2847" lane="5" entrytime="00:00:34.87" entrycourse="LCM" />
                <RESULT eventid="1103" points="228" swimtime="00:01:20.85" resultid="1734" heatid="2779" lane="4" entrytime="00:01:19.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="261" swimtime="00:00:32.68" resultid="1735" heatid="2905" lane="2" entrytime="00:00:32.50" entrycourse="LCM" />
                <RESULT eventid="1195" points="238" swimtime="00:03:03.93" resultid="1736" heatid="2879" lane="4" entrytime="00:03:05.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.01" />
                    <SPLIT distance="100" swimtime="00:01:25.54" />
                    <SPLIT distance="150" swimtime="00:02:24.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Betina" lastname="Vieira Pellanda" birthdate="2014-02-16" gender="F" nation="BRA" license="391041" swrid="5602589" athleteid="1991" externalid="391041">
              <RESULTS>
                <RESULT eventid="1068" points="179" swimtime="00:03:19.95" resultid="1992" heatid="2740" lane="6" entrytime="00:03:25.17" entrycourse="LCM" />
                <RESULT eventid="1080" points="129" swimtime="00:00:57.62" resultid="1993" heatid="2754" lane="6" />
                <RESULT eventid="1152" points="162" swimtime="00:03:51.23" resultid="1994" heatid="2836" lane="3" entrytime="00:03:58.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.91" />
                    <SPLIT distance="100" swimtime="00:01:54.13" />
                    <SPLIT distance="150" swimtime="00:03:03.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="169" swimtime="00:00:42.63" resultid="1995" heatid="2886" lane="2" entrytime="00:00:43.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Cipriani Presiazniuk" birthdate="2012-07-03" gender="M" nation="BRA" license="369267" swrid="5588594" athleteid="1687" externalid="369267">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="1688" heatid="2768" lane="6" entrytime="00:01:30.49" entrycourse="LCM" />
                <RESULT eventid="1149" status="DNS" swimtime="00:00:00.00" resultid="1689" heatid="2832" lane="4" entrytime="00:02:53.37" entrycourse="LCM" />
                <RESULT eventid="1119" status="DNS" swimtime="00:00:00.00" resultid="1690" heatid="2796" lane="7" entrytime="00:00:39.75" entrycourse="LCM" />
                <RESULT eventid="1195" status="DNS" swimtime="00:00:00.00" resultid="1691" heatid="2878" lane="4" entrytime="00:03:23.29" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="De Moraes" birthdate="2014-09-18" gender="M" nation="BRA" license="391024" swrid="5602529" athleteid="1971" externalid="391024">
              <RESULTS>
                <RESULT eventid="1071" points="189" swimtime="00:02:57.69" resultid="1972" heatid="2743" lane="6" entrytime="00:03:17.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                    <SPLIT distance="100" swimtime="00:01:23.77" />
                    <SPLIT distance="150" swimtime="00:02:11.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="161" swimtime="00:03:29.31" resultid="1973" heatid="2839" lane="3" entrytime="00:03:35.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.92" />
                    <SPLIT distance="100" swimtime="00:01:39.29" />
                    <SPLIT distance="150" swimtime="00:02:43.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="165" swimtime="00:00:40.53" resultid="1974" heatid="2786" lane="6" entrytime="00:00:47.15" entrycourse="LCM" />
                <RESULT eventid="1205" points="207" swimtime="00:00:35.31" resultid="1975" heatid="2893" lane="7" entrytime="00:00:38.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia" lastname="Ziliotto Mehl" birthdate="2015-10-09" gender="F" nation="BRA" license="400122" swrid="5652905" athleteid="2086" externalid="400122">
              <RESULTS>
                <RESULT eventid="1068" points="119" swimtime="00:03:48.96" resultid="2087" heatid="2738" lane="4" />
                <RESULT eventid="1080" points="116" swimtime="00:00:59.69" resultid="2088" heatid="2754" lane="4" entrytime="00:01:10.32" entrycourse="LCM" />
                <RESULT eventid="1106" points="69" swimtime="00:00:59.52" resultid="2089" heatid="2782" lane="2" entrytime="00:01:15.49" entrycourse="LCM" />
                <RESULT eventid="1202" points="172" swimtime="00:00:42.40" resultid="2090" heatid="2885" lane="8" entrytime="00:00:52.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Spadari Soso" birthdate="2012-12-28" gender="F" nation="BRA" license="377313" swrid="5588921" athleteid="2141" externalid="377313">
              <RESULTS>
                <RESULT eventid="1074" points="273" swimtime="00:00:44.90" resultid="2142" heatid="2744" lane="7" />
                <RESULT eventid="1146" points="405" swimtime="00:02:32.48" resultid="2143" heatid="2829" lane="6" entrytime="00:02:58.08" entrycourse="LCM" />
                <RESULT eventid="1170" points="286" swimtime="00:01:37.26" resultid="2144" heatid="2861" lane="1" entrytime="00:01:50.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="419" swimtime="00:00:31.53" resultid="2145" heatid="2898" lane="4" entrytime="00:00:35.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Artigas Pinheiro" birthdate="2013-07-31" gender="F" nation="BRA" license="377153" swrid="5588534" athleteid="1886" externalid="377153">
              <RESULTS>
                <RESULT eventid="1086" points="221" swimtime="00:01:34.78" resultid="1887" heatid="2763" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1158" points="115" swimtime="00:00:50.21" resultid="1888" heatid="2842" lane="2" entrytime="00:00:51.30" entrycourse="LCM" />
                <RESULT eventid="1132" points="233" swimtime="00:01:23.99" resultid="1889" heatid="2813" lane="5" entrytime="00:01:31.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="195" swimtime="00:03:37.40" resultid="1890" heatid="2875" lane="6" entrytime="00:03:45.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.25" />
                    <SPLIT distance="100" swimtime="00:01:44.86" />
                    <SPLIT distance="150" swimtime="00:02:55.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Saporiti Salvi" birthdate="2013-06-28" gender="M" nation="BRA" license="377032" swrid="5588896" athleteid="1836" externalid="377032">
              <RESULTS>
                <RESULT eventid="1077" points="125" swimtime="00:00:51.77" resultid="1837" heatid="2750" lane="8" entrytime="00:00:53.40" entrycourse="LCM" />
                <RESULT eventid="1149" points="235" swimtime="00:02:45.16" resultid="1838" heatid="2832" lane="3" entrytime="00:02:56.42" entrycourse="LCM" />
                <RESULT eventid="1103" points="167" swimtime="00:01:29.67" resultid="1839" heatid="2778" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="215" swimtime="00:03:10.25" resultid="1840" heatid="2878" lane="5" entrytime="00:03:23.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.20" />
                    <SPLIT distance="100" swimtime="00:01:31.38" />
                    <SPLIT distance="150" swimtime="00:02:32.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Fernandes Tramujas" birthdate="2015-01-15" gender="F" nation="BRA" license="406750" swrid="5717263" athleteid="2136" externalid="406750">
              <RESULTS>
                <RESULT eventid="1068" points="90" swimtime="00:04:11.15" resultid="2137" heatid="2738" lane="3" />
                <RESULT eventid="1080" points="70" swimtime="00:01:10.52" resultid="2138" heatid="2754" lane="7" />
                <RESULT eventid="1164" points="66" reactiontime="+84" swimtime="00:01:06.35" resultid="2139" heatid="2848" lane="4" />
                <RESULT eventid="1122" points="81" swimtime="00:01:59.16" resultid="2140" heatid="2800" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Szpak Zraik" birthdate="2015-04-10" gender="M" nation="BRA" license="393259" swrid="5616451" athleteid="2011" externalid="393259">
              <RESULTS>
                <RESULT eventid="1071" points="99" swimtime="00:03:40.19" resultid="2012" heatid="2742" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.67" />
                    <SPLIT distance="150" swimtime="00:02:43.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="132" swimtime="00:00:50.96" resultid="2013" heatid="2762" lane="2" entrytime="00:00:54.54" entrycourse="LCM" />
                <RESULT eventid="1155" points="105" swimtime="00:04:01.60" resultid="2014" heatid="2838" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:05.04" />
                    <SPLIT distance="150" swimtime="00:03:06.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="98" swimtime="00:01:41.34" resultid="2015" heatid="2804" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cecilia Carvalho" birthdate="2014-10-30" gender="F" nation="BRA" license="391021" swrid="5602525" athleteid="1961" externalid="391021">
              <RESULTS>
                <RESULT eventid="1068" status="DNS" swimtime="00:00:00.00" resultid="1962" heatid="2740" lane="8" entrytime="00:04:17.55" entrycourse="LCM" />
                <RESULT eventid="1106" status="DNS" swimtime="00:00:00.00" resultid="1963" heatid="2782" lane="8" />
                <RESULT eventid="1164" status="DNS" swimtime="00:00:00.00" resultid="1964" heatid="2851" lane="2" entrytime="00:01:00.22" entrycourse="LCM" />
                <RESULT eventid="1122" status="DNS" swimtime="00:00:00.00" resultid="1965" heatid="2800" lane="2" entrytime="00:02:05.11" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Alice Silva Gomes Xavier" birthdate="2013-02-25" gender="F" nation="BRA" license="371040" swrid="5717241" athleteid="2156" externalid="371040">
              <RESULTS>
                <RESULT eventid="1074" points="300" swimtime="00:00:43.54" resultid="2157" heatid="2747" lane="2" entrytime="00:00:46.04" entrycourse="LCM" />
                <RESULT eventid="1132" points="361" swimtime="00:01:12.56" resultid="2158" heatid="2815" lane="6" entrytime="00:01:16.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="293" swimtime="00:01:36.52" resultid="2159" heatid="2861" lane="2" entrytime="00:01:41.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="374" swimtime="00:00:32.75" resultid="2160" heatid="2899" lane="7" entrytime="00:00:34.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Prosdocimo" birthdate="2012-11-30" gender="M" nation="BRA" license="369272" swrid="5602575" athleteid="1707" externalid="369272">
              <RESULTS>
                <RESULT eventid="1065" points="300" swimtime="00:05:28.53" resultid="1708" heatid="2736" lane="4" entrytime="00:05:32.70" entrycourse="LCM" />
                <RESULT eventid="1149" points="278" swimtime="00:02:36.19" resultid="1709" heatid="2833" lane="2" entrytime="00:02:39.68" entrycourse="LCM" />
                <RESULT eventid="1119" points="231" swimtime="00:00:38.33" resultid="1710" heatid="2796" lane="1" entrytime="00:00:40.24" entrycourse="LCM" />
                <RESULT eventid="1211" points="265" swimtime="00:00:32.53" resultid="1711" heatid="2904" lane="7" entrytime="00:00:34.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Miranda Carvalho" birthdate="2015-07-07" gender="F" nation="BRA" license="410200" athleteid="2186" externalid="410200">
              <RESULTS>
                <RESULT eventid="1080" points="75" swimtime="00:01:09.01" resultid="2187" heatid="2753" lane="3" />
                <RESULT eventid="1164" points="73" reactiontime="+44" swimtime="00:01:04.00" resultid="2188" heatid="2850" lane="7" />
                <RESULT eventid="1122" points="57" swimtime="00:02:14.19" resultid="2189" heatid="2799" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="72" swimtime="00:00:56.54" resultid="2190" heatid="2882" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Wolff Contin" birthdate="2015-10-10" gender="M" nation="BRA" license="406745" swrid="5717303" athleteid="2116" externalid="406745">
              <RESULTS>
                <RESULT eventid="1071" points="68" swimtime="00:04:09.84" resultid="2117" heatid="2742" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.59" />
                    <SPLIT distance="100" swimtime="00:01:58.65" />
                    <SPLIT distance="150" swimtime="00:03:07.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="48" swimtime="00:01:04.76" resultid="2118" heatid="2853" lane="4" />
                <RESULT eventid="1125" points="58" swimtime="00:02:00.58" resultid="2119" heatid="2803" lane="3" />
                <RESULT eventid="1205" points="70" swimtime="00:00:50.69" resultid="2120" heatid="2889" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Liam" lastname="Batista Grise" birthdate="2014-03-27" gender="M" nation="BRA" license="391008" swrid="5602514" athleteid="1926" externalid="391008">
              <RESULTS>
                <RESULT eventid="1083" points="105" swimtime="00:00:54.92" resultid="1927" heatid="2760" lane="4" entrytime="00:01:07.81" entrycourse="LCM" />
                <RESULT eventid="1167" points="72" reactiontime="+58" swimtime="00:00:56.44" resultid="1928" heatid="2857" lane="1" entrytime="00:00:56.56" entrycourse="LCM" />
                <RESULT eventid="1125" points="91" swimtime="00:01:43.84" resultid="1929" heatid="2807" lane="1" entrytime="00:01:49.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="107" swimtime="00:00:43.92" resultid="1930" heatid="2891" lane="6" entrytime="00:00:47.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Pisani Ferreira" birthdate="2012-08-06" gender="F" nation="BRA" license="376985" swrid="5588862" athleteid="1876" externalid="376985">
              <RESULTS>
                <RESULT eventid="1074" points="226" swimtime="00:00:47.85" resultid="1877" heatid="2746" lane="5" entrytime="00:00:50.39" entrycourse="LCM" />
                <RESULT eventid="1132" points="183" swimtime="00:01:30.94" resultid="1878" heatid="2811" lane="2" />
                <RESULT eventid="1170" points="218" swimtime="00:01:46.43" resultid="1879" heatid="2861" lane="8" entrytime="00:01:54.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="202" swimtime="00:00:40.19" resultid="1880" heatid="2897" lane="1" entrytime="00:00:41.51" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Saber" birthdate="2014-06-04" gender="F" nation="BRA" license="392141" swrid="5602554" athleteid="2001" externalid="392141">
              <RESULTS>
                <RESULT eventid="1080" points="177" swimtime="00:00:51.88" resultid="2002" heatid="2756" lane="1" entrytime="00:00:59.19" entrycourse="LCM" />
                <RESULT eventid="1152" points="156" swimtime="00:03:53.93" resultid="2003" heatid="2835" lane="4" entrytime="00:04:51.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.81" />
                    <SPLIT distance="100" swimtime="00:02:00.42" />
                    <SPLIT distance="150" swimtime="00:03:04.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="131" swimtime="00:00:52.79" resultid="2004" heatid="2851" lane="3" entrytime="00:00:58.98" entrycourse="LCM" />
                <RESULT eventid="1122" points="155" swimtime="00:01:36.24" resultid="2005" heatid="2800" lane="3" entrytime="00:01:51.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ravi" lastname="Osternack Erbe" birthdate="2013-08-10" gender="M" nation="BRA" license="372681" swrid="5588841" athleteid="1747" externalid="372681">
              <RESULTS>
                <RESULT eventid="1089" points="204" swimtime="00:01:27.59" resultid="1748" heatid="2767" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1149" status="DSQ" swimtime="00:02:45.13" resultid="1749" heatid="2832" lane="5" entrytime="00:02:56.16" entrycourse="LCM" />
                <RESULT eventid="1103" status="DSQ" swimtime="00:01:35.08" resultid="1750" heatid="2779" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="197" swimtime="00:00:35.91" resultid="1751" heatid="2904" lane="8" entrytime="00:00:35.36" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olavo" lastname="Valduga Artigas" birthdate="2012-06-26" gender="M" nation="BRA" license="369270" swrid="5588941" athleteid="1697" externalid="369270">
              <RESULTS>
                <RESULT eventid="1077" points="153" swimtime="00:00:48.49" resultid="1698" heatid="2751" lane="8" entrytime="00:00:45.83" entrycourse="LCM" />
                <RESULT eventid="1119" points="139" swimtime="00:00:45.41" resultid="1699" heatid="2792" lane="6" />
                <RESULT eventid="1173" points="148" swimtime="00:01:47.44" resultid="1700" heatid="2864" lane="1" entrytime="00:01:44.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="165" swimtime="00:03:27.72" resultid="1701" heatid="2879" lane="8" entrytime="00:03:21.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Henrique Tiboni Araujo" birthdate="2013-06-11" gender="M" nation="BRA" license="376968" swrid="5588747" athleteid="1791" externalid="376968">
              <RESULTS>
                <RESULT eventid="1089" points="130" swimtime="00:01:41.79" resultid="1792" heatid="2766" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="149" swimtime="00:01:28.29" resultid="1793" heatid="2819" lane="7" entrytime="00:01:32.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="133" swimtime="00:00:46.11" resultid="1794" heatid="2795" lane="8" entrytime="00:00:45.70" entrycourse="LCM" />
                <RESULT eventid="1195" points="128" swimtime="00:03:45.94" resultid="1795" heatid="2877" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.20" />
                    <SPLIT distance="100" swimtime="00:01:45.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Bernardi Pedrosa" birthdate="2013-03-09" gender="F" nation="BRA" license="376977" swrid="5588551" athleteid="1811" externalid="376977">
              <RESULTS>
                <RESULT eventid="1086" points="244" swimtime="00:01:31.64" resultid="1812" heatid="2764" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="260" swimtime="00:01:21.00" resultid="1813" heatid="2813" lane="6" entrytime="00:01:36.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="257" swimtime="00:00:42.24" resultid="1814" heatid="2790" lane="7" entrytime="00:00:49.07" entrycourse="LCM" />
                <RESULT eventid="1208" points="263" swimtime="00:00:36.84" resultid="1815" heatid="2897" lane="2" entrytime="00:00:40.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Schmidt Wozniaki" birthdate="2012-07-07" gender="M" nation="BRA" license="376963" swrid="5588905" athleteid="1782" externalid="376963">
              <RESULTS>
                <RESULT eventid="1077" points="124" swimtime="00:00:52.03" resultid="1783" heatid="2750" lane="7" entrytime="00:00:52.30" entrycourse="LCM" />
                <RESULT eventid="1119" points="115" swimtime="00:00:48.38" resultid="1784" heatid="2794" lane="7" entrytime="00:00:51.19" entrycourse="LCM" />
                <RESULT eventid="1173" points="104" swimtime="00:02:00.95" resultid="1785" heatid="2863" lane="5" entrytime="00:02:08.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Mayer Paludetto" birthdate="2012-10-30" gender="F" nation="BRA" license="369264" swrid="5588811" athleteid="1682" externalid="369264">
              <RESULTS>
                <RESULT eventid="1062" points="412" swimtime="00:05:16.15" resultid="1683" heatid="2733" lane="2" />
                <RESULT eventid="1146" points="409" swimtime="00:02:32.01" resultid="1684" heatid="2829" lane="5" entrytime="00:02:41.43" entrycourse="LCM" />
                <RESULT eventid="1100" points="274" swimtime="00:01:25.33" resultid="1685" heatid="2776" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="383" swimtime="00:02:53.55" resultid="1686" heatid="2876" lane="4" entrytime="00:03:00.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                    <SPLIT distance="100" swimtime="00:01:23.69" />
                    <SPLIT distance="150" swimtime="00:02:15.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Moreira Pasqual" birthdate="2014-07-09" gender="M" nation="BRA" license="382125" swrid="5602562" athleteid="1901" externalid="382125">
              <RESULTS>
                <RESULT eventid="1071" status="DNS" swimtime="00:00:00.00" resultid="1902" heatid="2743" lane="7" entrytime="00:03:42.12" entrycourse="LCM" />
                <RESULT eventid="1155" status="DNS" swimtime="00:00:00.00" resultid="1903" heatid="2839" lane="2" entrytime="00:04:12.28" entrycourse="LCM" />
                <RESULT eventid="1125" status="DNS" swimtime="00:00:00.00" resultid="1904" heatid="2807" lane="4" entrytime="00:01:41.44" entrycourse="LCM" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="1905" heatid="2892" lane="5" entrytime="00:00:42.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Albuquerque" birthdate="2012-11-16" gender="F" nation="BRA" license="369281" swrid="5602506" athleteid="1737" externalid="369281">
              <RESULTS>
                <RESULT eventid="1062" points="333" swimtime="00:05:39.27" resultid="1738" heatid="2734" lane="2" entrytime="00:05:55.07" entrycourse="LCM" />
                <RESULT eventid="1100" points="274" swimtime="00:01:25.35" resultid="1739" heatid="2777" lane="3" entrytime="00:01:33.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="305" swimtime="00:01:35.21" resultid="1740" heatid="2861" lane="6" entrytime="00:01:40.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="344" swimtime="00:02:59.96" resultid="1741" heatid="2876" lane="2" entrytime="00:03:12.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.59" />
                    <SPLIT distance="100" swimtime="00:01:27.83" />
                    <SPLIT distance="150" swimtime="00:02:20.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Pens Correa" birthdate="2015-11-27" gender="M" nation="BRA" license="393262" swrid="5616449" athleteid="2026" externalid="393262">
              <RESULTS>
                <RESULT eventid="1071" points="178" swimtime="00:03:01.08" resultid="2027" heatid="2742" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                    <SPLIT distance="100" swimtime="00:01:26.86" />
                    <SPLIT distance="150" swimtime="00:02:15.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="165" swimtime="00:03:27.48" resultid="2028" heatid="2838" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                    <SPLIT distance="100" swimtime="00:01:30.23" />
                    <SPLIT distance="150" swimtime="00:02:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="167" swimtime="00:00:40.39" resultid="2029" heatid="2786" lane="2" entrytime="00:00:47.84" entrycourse="LCM" />
                <RESULT eventid="1167" points="185" swimtime="00:00:41.28" resultid="2030" heatid="2858" lane="5" entrytime="00:00:45.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Marie Silva" birthdate="2014-08-24" gender="F" nation="BRA" license="391025" swrid="5602556" athleteid="1976" externalid="391025">
              <RESULTS>
                <RESULT eventid="1068" points="174" swimtime="00:03:22.07" resultid="1977" heatid="2740" lane="7" entrytime="00:03:50.55" entrycourse="LCM" />
                <RESULT eventid="1152" points="145" swimtime="00:03:59.93" resultid="1978" heatid="2836" lane="2" entrytime="00:04:12.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.37" />
                    <SPLIT distance="100" swimtime="00:02:04.96" />
                    <SPLIT distance="150" swimtime="00:03:11.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1106" points="118" swimtime="00:00:49.69" resultid="1979" heatid="2780" lane="4" />
                <RESULT eventid="1122" points="180" swimtime="00:01:31.58" resultid="1980" heatid="2801" lane="1" entrytime="00:01:42.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Cury Abreu" birthdate="2013-05-17" gender="F" nation="BRA" license="376974" swrid="5588614" athleteid="1801" externalid="376974">
              <RESULTS>
                <RESULT eventid="1086" points="270" swimtime="00:01:28.64" resultid="1802" heatid="2764" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1132" points="295" swimtime="00:01:17.65" resultid="1803" heatid="2814" lane="3" entrytime="00:01:23.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="316" swimtime="00:00:39.41" resultid="1804" heatid="2790" lane="8" entrytime="00:00:50.14" entrycourse="LCM" />
                <RESULT eventid="1208" points="347" swimtime="00:00:33.59" resultid="1805" heatid="2898" lane="7" entrytime="00:00:36.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Ribas Luz" birthdate="2015-02-05" gender="F" nation="BRA" license="406743" swrid="5717291" athleteid="2111" externalid="406743">
              <RESULTS>
                <RESULT eventid="1080" points="43" swimtime="00:01:22.80" resultid="2112" heatid="2754" lane="1" />
                <RESULT eventid="1164" points="101" swimtime="00:00:57.53" resultid="2113" heatid="2849" lane="5" />
                <RESULT eventid="1122" points="68" swimtime="00:02:06.25" resultid="2114" heatid="2798" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="101" swimtime="00:00:50.61" resultid="2115" heatid="2883" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Shwetz Clivatti" birthdate="2015-03-05" gender="M" nation="BRA" license="406963" swrid="5717297" athleteid="2171" externalid="406963">
              <RESULTS>
                <RESULT eventid="1083" points="38" swimtime="00:01:16.70" resultid="2172" heatid="2757" lane="5" />
                <RESULT eventid="1167" points="46" reactiontime="+59" swimtime="00:01:05.36" resultid="2173" heatid="2855" lane="8" />
                <RESULT eventid="1125" points="43" swimtime="00:02:13.20" resultid="2174" heatid="2802" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="30" swimtime="00:01:06.93" resultid="2175" heatid="2888" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Puppi Cardoso" birthdate="2015-03-30" gender="F" nation="BRA" license="406741" swrid="5717289" athleteid="2101" externalid="406741">
              <RESULTS>
                <RESULT eventid="1080" points="81" swimtime="00:01:07.31" resultid="2102" heatid="2753" lane="5" />
                <RESULT eventid="1152" points="80" swimtime="00:04:51.52" resultid="2103" heatid="2834" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.67" />
                    <SPLIT distance="100" swimtime="00:02:19.58" />
                    <SPLIT distance="150" swimtime="00:03:46.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1106" points="47" swimtime="00:01:07.31" resultid="2104" heatid="2781" lane="8" />
                <RESULT eventid="1164" points="106" swimtime="00:00:56.75" resultid="2105" heatid="2850" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="De Fortes" birthdate="2015-06-01" gender="M" nation="BRA" license="399680" swrid="5652884" athleteid="2071" externalid="399680">
              <RESULTS>
                <RESULT eventid="1071" points="87" swimtime="00:03:49.34" resultid="2072" heatid="2742" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.98" />
                    <SPLIT distance="100" swimtime="00:01:50.71" />
                    <SPLIT distance="150" swimtime="00:02:51.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="85" swimtime="00:04:19.14" resultid="2073" heatid="2838" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.07" />
                    <SPLIT distance="100" swimtime="00:02:00.34" />
                    <SPLIT distance="150" swimtime="00:03:24.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="84" swimtime="00:00:50.80" resultid="2074" heatid="2785" lane="3" entrytime="00:01:08.79" entrycourse="LCM" />
                <RESULT eventid="1167" points="87" reactiontime="+69" swimtime="00:00:52.95" resultid="2075" heatid="2856" lane="5" entrytime="00:01:00.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivia" lastname="Mayer Paludetto" birthdate="2016-04-01" gender="F" nation="BRA" license="412014" athleteid="2209" externalid="412014">
              <RESULTS>
                <RESULT eventid="1128" points="109" swimtime="00:00:56.13" resultid="2210" heatid="2809" lane="6" />
                <RESULT eventid="1214" points="104" swimtime="00:00:50.17" resultid="2211" heatid="2906" lane="3" />
                <RESULT eventid="1198" points="101" swimtime="00:01:02.43" resultid="2212" heatid="2880" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Felipe Canalli" birthdate="2015-12-23" gender="M" nation="BRA" license="406749" swrid="5717261" athleteid="2131" externalid="406749">
              <RESULTS>
                <RESULT eventid="1083" points="100" swimtime="00:00:55.85" resultid="2132" heatid="2759" lane="7" />
                <RESULT eventid="1155" points="60" swimtime="00:04:49.80" resultid="2133" heatid="2839" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:32.62" />
                    <SPLIT distance="150" swimtime="00:03:42.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="56" swimtime="00:00:58.16" resultid="2134" heatid="2785" lane="7" />
                <RESULT eventid="1125" points="49" swimtime="00:02:07.81" resultid="2135" heatid="2803" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Cabrini Vieira" birthdate="2012-02-11" gender="F" nation="BRA" license="376961" swrid="5588571" athleteid="1772" externalid="376961">
              <RESULTS>
                <RESULT eventid="1062" points="437" swimtime="00:05:09.97" resultid="1773" heatid="2734" lane="3" entrytime="00:05:30.09" entrycourse="LCM" />
                <RESULT eventid="1086" points="403" swimtime="00:01:17.59" resultid="1774" heatid="2765" lane="5" entrytime="00:01:23.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="443" swimtime="00:00:35.22" resultid="1775" heatid="2791" lane="4" entrytime="00:00:38.27" entrycourse="LCM" />
                <RESULT eventid="1208" points="502" swimtime="00:00:29.69" resultid="1776" heatid="2899" lane="4" entrytime="00:00:32.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Guimaraes Mesquita" birthdate="2015-10-05" gender="F" nation="BRA" license="393263" swrid="5616444" athleteid="2031" externalid="393263">
              <RESULTS>
                <RESULT eventid="1080" points="71" swimtime="00:01:10.17" resultid="2032" heatid="2753" lane="2" />
                <RESULT eventid="1164" points="77" swimtime="00:01:03.07" resultid="2033" heatid="2849" lane="6" />
                <RESULT eventid="1122" points="56" swimtime="00:02:14.99" resultid="2034" heatid="2799" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="71" swimtime="00:00:56.88" resultid="2035" heatid="2884" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Antunes Saboia" birthdate="2012-06-28" gender="M" nation="BRA" license="369278" swrid="5602511" athleteid="1727" externalid="369278">
              <RESULTS>
                <RESULT eventid="1077" points="249" swimtime="00:00:41.24" resultid="1728" heatid="2751" lane="6" entrytime="00:00:42.02" entrycourse="LCM" />
                <RESULT eventid="1135" points="291" swimtime="00:01:10.67" resultid="1729" heatid="2821" lane="1" entrytime="00:01:14.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="248" swimtime="00:01:30.44" resultid="1730" heatid="2864" lane="3" entrytime="00:01:32.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="265" swimtime="00:02:57.39" resultid="1731" heatid="2879" lane="5" entrytime="00:03:07.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.37" />
                    <SPLIT distance="100" swimtime="00:01:27.88" />
                    <SPLIT distance="150" swimtime="00:02:20.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Salomao" birthdate="2012-05-07" gender="M" nation="BRA" license="369261" swrid="5602581" athleteid="1672" externalid="369261">
              <RESULTS>
                <RESULT eventid="1065" points="299" swimtime="00:05:28.77" resultid="1673" heatid="2736" lane="5" entrytime="00:05:33.00" entrycourse="LCM" />
                <RESULT eventid="1149" points="273" swimtime="00:02:37.17" resultid="1674" heatid="2833" lane="6" entrytime="00:02:39.09" entrycourse="LCM" />
                <RESULT eventid="1135" points="273" swimtime="00:01:12.22" resultid="1675" heatid="2821" lane="2" entrytime="00:01:12.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="265" swimtime="00:00:32.53" resultid="1676" heatid="2904" lane="4" entrytime="00:00:32.89" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Pisani Ferreira" birthdate="2014-01-26" gender="M" nation="BRA" license="391017" swrid="5602570" athleteid="1941" externalid="391017">
              <RESULTS>
                <RESULT eventid="1083" status="DNS" swimtime="00:00:00.00" resultid="1942" heatid="2762" lane="8" entrytime="00:00:57.70" entrycourse="LCM" />
                <RESULT eventid="1155" status="DNS" swimtime="00:00:00.00" resultid="1943" heatid="2839" lane="1" entrytime="00:04:27.43" entrycourse="LCM" />
                <RESULT eventid="1125" status="DNS" swimtime="00:00:00.00" resultid="1944" heatid="2802" lane="4" />
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="1945" heatid="2889" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Livia Bittencourt" birthdate="2015-11-23" gender="F" nation="BRA" license="393260" swrid="5616446" athleteid="2016" externalid="393260">
              <RESULTS>
                <RESULT eventid="1068" status="DNS" swimtime="00:00:00.00" resultid="2017" heatid="2737" lane="4" />
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="2018" heatid="2754" lane="5" entrytime="00:01:22.77" entrycourse="LCM" />
                <RESULT eventid="1106" status="DNS" swimtime="00:00:00.00" resultid="2019" heatid="2782" lane="7" entrytime="00:01:30.10" entrycourse="LCM" />
                <RESULT eventid="1122" status="DNS" swimtime="00:00:00.00" resultid="2020" heatid="2799" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Almeida Jorge" birthdate="2015-05-27" gender="M" nation="BRA" license="406836" swrid="5717242" athleteid="2146" externalid="406836">
              <RESULTS>
                <RESULT eventid="1083" points="63" swimtime="00:01:04.95" resultid="2147" heatid="2760" lane="7" />
                <RESULT eventid="1167" points="66" reactiontime="+79" swimtime="00:00:58.23" resultid="2148" heatid="2855" lane="5" />
                <RESULT eventid="1125" points="36" swimtime="00:02:21.31" resultid="2149" heatid="2803" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="36" swimtime="00:01:03.14" resultid="2150" heatid="2889" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Paulo Celles" birthdate="2016-09-07" gender="M" nation="BRA" license="411996" athleteid="2201" externalid="411996">
              <RESULTS>
                <RESULT eventid="1216" points="28" swimtime="00:01:08.21" resultid="2202" heatid="2907" lane="4" />
                <RESULT eventid="1200" points="31" swimtime="00:01:21.96" resultid="2203" heatid="2881" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Portes Fabiane" birthdate="2012-12-28" gender="M" nation="BRA" license="376983" swrid="5588864" athleteid="1826" externalid="376983">
              <RESULTS>
                <RESULT eventid="1089" points="80" swimtime="00:01:59.49" resultid="1827" heatid="2767" lane="5" entrytime="00:02:07.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="77" swimtime="00:01:49.98" resultid="1828" heatid="2818" lane="1" entrytime="00:01:48.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="75" swimtime="00:00:55.83" resultid="1829" heatid="2793" lane="4" entrytime="00:00:57.26" entrycourse="LCM" />
                <RESULT eventid="1211" points="105" swimtime="00:00:44.30" resultid="1830" heatid="2901" lane="3" entrytime="00:00:46.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Alzamora Calado" birthdate="2013-04-26" gender="F" nation="BRA" license="376960" swrid="5588522" athleteid="1767" externalid="376960">
              <RESULTS>
                <RESULT eventid="1074" points="253" swimtime="00:00:46.06" resultid="1768" heatid="2747" lane="1" entrytime="00:00:47.83" entrycourse="LCM" />
                <RESULT eventid="1132" points="313" swimtime="00:01:16.15" resultid="1769" heatid="2815" lane="1" entrytime="00:01:21.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="236" swimtime="00:01:43.65" resultid="1770" heatid="2860" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="301" swimtime="00:00:35.20" resultid="1771" heatid="2899" lane="8" entrytime="00:00:35.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="De Almeida Dias" birthdate="2012-02-18" gender="F" nation="BRA" license="369262" swrid="5588638" athleteid="1677" externalid="369262">
              <RESULTS>
                <RESULT eventid="1062" points="421" swimtime="00:05:14.02" resultid="1678" heatid="2734" lane="8" />
                <RESULT eventid="1146" points="443" swimtime="00:02:27.93" resultid="1679" heatid="2829" lane="4" entrytime="00:02:30.70" entrycourse="LCM" />
                <RESULT eventid="1132" points="452" swimtime="00:01:07.35" resultid="1680" heatid="2815" lane="4" entrytime="00:01:08.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="448" swimtime="00:00:30.85" resultid="1681" heatid="2899" lane="5" entrytime="00:00:32.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Tallao Benke" birthdate="2012-01-02" gender="F" nation="BRA" license="376984" swrid="5588931" athleteid="1831" externalid="376984">
              <RESULTS>
                <RESULT eventid="1062" points="454" swimtime="00:05:06.18" resultid="1832" heatid="2734" lane="5" entrytime="00:05:18.33" entrycourse="LCM" />
                <RESULT eventid="1086" points="426" swimtime="00:01:16.17" resultid="1833" heatid="2765" lane="4" entrytime="00:01:16.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="467" swimtime="00:02:25.43" resultid="1834" heatid="2828" lane="7" />
                <RESULT eventid="1100" points="407" swimtime="00:01:14.85" resultid="1835" heatid="2777" lane="4" entrytime="00:01:17.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Zagonel Krempel" birthdate="2015-07-27" gender="F" nation="BRA" license="406962" swrid="5717305" athleteid="2166" externalid="406962">
              <RESULTS>
                <RESULT eventid="1080" points="82" swimtime="00:01:06.98" resultid="2167" heatid="2752" lane="3" />
                <RESULT eventid="1164" points="91" reactiontime="+65" swimtime="00:00:59.60" resultid="2168" heatid="2849" lane="2" />
                <RESULT eventid="1122" points="56" swimtime="00:02:15.15" resultid="2169" heatid="2797" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="72" swimtime="00:00:56.63" resultid="2170" heatid="2883" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Emilia Abrahao" birthdate="2016-06-14" gender="F" nation="BRA" license="412012" athleteid="2204" externalid="412012">
              <RESULTS>
                <RESULT eventid="1214" points="55" swimtime="00:01:01.96" resultid="2205" heatid="2906" lane="2" />
                <RESULT eventid="1198" points="81" swimtime="00:01:07.35" resultid="2206" heatid="2880" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Magalhaes Dabul" birthdate="2014-01-05" gender="M" nation="BRA" license="391023" swrid="5602555" athleteid="1966" externalid="391023">
              <RESULTS>
                <RESULT eventid="1083" points="131" swimtime="00:00:51.05" resultid="1967" heatid="2761" lane="5" entrytime="00:01:00.60" entrycourse="LCM" />
                <RESULT eventid="1155" points="130" swimtime="00:03:44.58" resultid="1968" heatid="2839" lane="7" entrytime="00:04:15.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.51" />
                    <SPLIT distance="100" swimtime="00:01:46.98" />
                    <SPLIT distance="150" swimtime="00:02:53.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="134" swimtime="00:00:43.50" resultid="1969" heatid="2785" lane="4" entrytime="00:01:00.58" entrycourse="LCM" />
                <RESULT eventid="1125" points="110" swimtime="00:01:37.53" resultid="1970" heatid="2806" lane="4" entrytime="00:01:55.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Taborda Ribas" birthdate="2015-12-30" gender="M" nation="BRA" license="406748" swrid="5717299" athleteid="2126" externalid="406748">
              <RESULTS>
                <RESULT eventid="1071" points="68" swimtime="00:04:09.76" resultid="2127" heatid="2741" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:56.21" />
                    <SPLIT distance="150" swimtime="00:03:03.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1155" points="55" swimtime="00:04:58.75" resultid="2128" heatid="2838" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.00" />
                    <SPLIT distance="100" swimtime="00:02:31.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1125" points="67" swimtime="00:01:55.17" resultid="2129" heatid="2803" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="76" swimtime="00:00:49.17" resultid="2130" heatid="2888" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Schiavo Vianna" birthdate="2013-04-27" gender="F" nation="BRA" license="391005" swrid="5602582" athleteid="1916" externalid="391005">
              <RESULTS>
                <RESULT eventid="1074" points="203" swimtime="00:00:49.54" resultid="1917" heatid="2746" lane="3" entrytime="00:00:51.96" entrycourse="LCM" />
                <RESULT eventid="1132" points="188" swimtime="00:01:30.23" resultid="1918" heatid="2812" lane="6" entrytime="00:01:48.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="174" swimtime="00:01:54.87" resultid="1919" heatid="2859" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="247" swimtime="00:00:37.58" resultid="1920" heatid="2895" lane="4" entrytime="00:00:49.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Coelho Ghignone" birthdate="2015-01-05" gender="M" nation="BRA" license="410201" athleteid="2191" externalid="410201">
              <RESULTS>
                <RESULT eventid="1083" points="56" swimtime="00:01:07.51" resultid="2192" heatid="2758" lane="7" />
                <RESULT eventid="1167" points="116" reactiontime="+49" swimtime="00:00:48.24" resultid="2193" heatid="2854" lane="5" />
                <RESULT eventid="1125" points="89" swimtime="00:01:44.70" resultid="2194" heatid="2806" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="100" swimtime="00:00:44.92" resultid="2195" heatid="2889" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Jarenko Gomes" birthdate="2014-05-17" gender="F" nation="BRA" license="407692" swrid="5725992" athleteid="2181" externalid="407692">
              <RESULTS>
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="2182" heatid="2754" lane="8" />
                <RESULT eventid="1106" status="DNS" swimtime="00:00:00.00" resultid="2183" heatid="2781" lane="4" />
                <RESULT eventid="1164" status="DNS" swimtime="00:00:00.00" resultid="2184" heatid="2849" lane="3" />
                <RESULT eventid="1202" points="84" swimtime="00:00:53.75" resultid="2185" heatid="2882" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Stramandinoli Zanicotti" birthdate="2013-06-18" gender="F" nation="BRA" license="376967" swrid="5588924" athleteid="1786" externalid="376967">
              <RESULTS>
                <RESULT eventid="1074" points="133" swimtime="00:00:57.12" resultid="1787" heatid="2746" lane="8" entrytime="00:01:00.32" entrycourse="LCM" />
                <RESULT eventid="1116" points="151" swimtime="00:00:50.37" resultid="1788" heatid="2789" lane="5" entrytime="00:00:50.80" entrycourse="LCM" />
                <RESULT eventid="1170" points="130" swimtime="00:02:06.36" resultid="1789" heatid="2860" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="164" swimtime="00:00:43.05" resultid="1790" heatid="2896" lane="1" entrytime="00:00:46.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Fonseca Ribeiro" birthdate="2016-02-25" gender="F" nation="BRA" license="412016" athleteid="2216" externalid="412016">
              <RESULTS>
                <RESULT eventid="1128" points="65" swimtime="00:01:06.47" resultid="2217" heatid="2809" lane="4" />
                <RESULT eventid="1214" points="76" swimtime="00:00:55.56" resultid="2218" heatid="2906" lane="5" />
                <RESULT eventid="1198" points="72" swimtime="00:01:09.84" resultid="2219" heatid="2880" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Rossi Mattioli" birthdate="2013-05-08" gender="F" nation="BRA" license="376988" swrid="5588892" athleteid="1866" externalid="376988">
              <RESULTS>
                <RESULT eventid="1062" points="245" swimtime="00:06:16.06" resultid="1867" heatid="2733" lane="3" />
                <RESULT eventid="1146" points="267" swimtime="00:02:55.24" resultid="1868" heatid="2829" lane="8" entrytime="00:03:13.02" entrycourse="LCM" />
                <RESULT eventid="1116" points="269" swimtime="00:00:41.58" resultid="1869" heatid="2791" lane="8" entrytime="00:00:43.15" entrycourse="LCM" />
                <RESULT eventid="1208" points="335" swimtime="00:00:33.97" resultid="1870" heatid="2898" lane="3" entrytime="00:00:36.03" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Gonçalves Sperandio" birthdate="2013-05-22" gender="M" nation="BRA" license="376980" swrid="5588851" athleteid="1816" externalid="376980">
              <RESULTS>
                <RESULT eventid="1065" points="248" swimtime="00:05:49.82" resultid="1817" heatid="2735" lane="3" />
                <RESULT eventid="1149" points="223" swimtime="00:02:48.01" resultid="1818" heatid="2833" lane="8" entrytime="00:02:51.95" entrycourse="LCM" />
                <RESULT eventid="1135" points="211" swimtime="00:01:18.62" resultid="1819" heatid="2820" lane="2" entrytime="00:01:19.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="194" swimtime="00:03:16.70" resultid="1820" heatid="2877" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.18" />
                    <SPLIT distance="100" swimtime="00:01:37.35" />
                    <SPLIT distance="150" swimtime="00:02:35.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Della Villa Yang" birthdate="2015-02-27" gender="F" nation="BRA" license="393283" swrid="5616442" athleteid="2041" externalid="393283">
              <RESULTS>
                <RESULT eventid="1068" points="146" swimtime="00:03:33.84" resultid="2042" heatid="2739" lane="4" />
                <RESULT eventid="1152" points="158" swimtime="00:03:52.98" resultid="2043" heatid="2834" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.58" />
                    <SPLIT distance="100" swimtime="00:01:53.00" />
                    <SPLIT distance="150" swimtime="00:03:00.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1106" points="108" swimtime="00:00:51.17" resultid="2044" heatid="2783" lane="6" entrytime="00:00:56.15" entrycourse="LCM" />
                <RESULT eventid="1202" points="155" swimtime="00:00:43.91" resultid="2045" heatid="2885" lane="1" entrytime="00:00:51.44" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Steven" lastname="Matheussi Viana E Silva" birthdate="2012-05-03" gender="M" nation="BRA" license="376986" swrid="5588810" athleteid="1871" externalid="376986">
              <RESULTS>
                <RESULT eventid="1077" points="239" swimtime="00:00:41.79" resultid="1872" heatid="2750" lane="5" entrytime="00:00:47.85" entrycourse="LCM" />
                <RESULT eventid="1161" points="212" swimtime="00:00:37.30" resultid="1873" heatid="2844" lane="6" />
                <RESULT eventid="1103" points="195" swimtime="00:01:25.23" resultid="1874" heatid="2779" lane="6" entrytime="00:01:30.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="226" swimtime="00:01:33.25" resultid="1875" heatid="2864" lane="7" entrytime="00:01:43.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Alice Palhano" birthdate="2016-04-06" gender="F" nation="BRA" license="412015" athleteid="2213" externalid="412015">
              <RESULTS>
                <RESULT eventid="1214" points="36" swimtime="00:01:10.88" resultid="2214" heatid="2906" lane="7" />
                <RESULT eventid="1198" points="50" swimtime="00:01:19.14" resultid="2215" heatid="2880" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Gois Nogueira" birthdate="2014-03-11" gender="F" nation="BRA" license="393258" swrid="5616443" athleteid="2006" externalid="393258">
              <RESULTS>
                <RESULT eventid="1080" points="139" swimtime="00:00:56.26" resultid="2007" heatid="2755" lane="7" entrytime="00:01:04.54" entrycourse="LCM" />
                <RESULT eventid="1106" points="77" swimtime="00:00:57.36" resultid="2008" heatid="2782" lane="6" entrytime="00:01:11.37" entrycourse="LCM" />
                <RESULT eventid="1164" points="139" reactiontime="+81" swimtime="00:00:51.82" resultid="2009" heatid="2851" lane="1" entrytime="00:01:03.15" entrycourse="LCM" />
                <RESULT eventid="1202" points="174" swimtime="00:00:42.23" resultid="2010" heatid="2884" lane="4" entrytime="00:00:54.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Vianna Almeida" birthdate="2014-12-16" gender="M" nation="BRA" license="410292" athleteid="2196" externalid="410292">
              <RESULTS>
                <RESULT eventid="1071" points="69" swimtime="00:04:07.62" resultid="2197" heatid="2743" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.35" />
                    <SPLIT distance="100" swimtime="00:01:55.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="74" swimtime="00:01:01.80" resultid="2198" heatid="2757" lane="6" />
                <RESULT eventid="1125" points="67" swimtime="00:01:55.12" resultid="2199" heatid="2806" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="69" swimtime="00:00:50.79" resultid="2200" heatid="2888" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maya" lastname="Assahida Moreria" birthdate="2014-02-24" gender="F" nation="BRA" license="391020" swrid="5602512" athleteid="1956" externalid="391020">
              <RESULTS>
                <RESULT eventid="1068" points="192" swimtime="00:03:15.45" resultid="1957" heatid="2740" lane="2" entrytime="00:03:27.08" entrycourse="LCM" />
                <RESULT eventid="1152" points="177" swimtime="00:03:44.41" resultid="1958" heatid="2836" lane="8" entrytime="00:04:24.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.32" />
                    <SPLIT distance="100" swimtime="00:01:50.40" />
                    <SPLIT distance="150" swimtime="00:02:55.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1106" points="145" swimtime="00:00:46.48" resultid="1959" heatid="2783" lane="1" entrytime="00:00:59.29" entrycourse="LCM" />
                <RESULT eventid="1122" points="189" swimtime="00:01:30.05" resultid="1960" heatid="2801" lane="2" entrytime="00:01:37.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Azevedo Alanis" birthdate="2013-12-07" gender="M" nation="BRA" license="376991" swrid="5588540" athleteid="1851" externalid="376991">
              <RESULTS>
                <RESULT eventid="1077" points="139" swimtime="00:00:50.09" resultid="1852" heatid="2749" lane="4" entrytime="00:00:54.02" entrycourse="LCM" />
                <RESULT eventid="1135" points="137" swimtime="00:01:30.72" resultid="1853" heatid="2818" lane="6" entrytime="00:01:40.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="141" swimtime="00:01:49.20" resultid="1854" heatid="2863" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1195" points="148" swimtime="00:03:35.20" resultid="1855" heatid="2878" lane="1" entrytime="00:03:51.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.62" />
                    <SPLIT distance="100" swimtime="00:01:43.65" />
                    <SPLIT distance="150" swimtime="00:02:47.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Cabrera Cirino Dos Santos" birthdate="2013-03-30" gender="M" nation="BRA" license="376990" swrid="5588570" athleteid="1856" externalid="376990">
              <RESULTS>
                <RESULT eventid="1065" points="227" swimtime="00:06:00.28" resultid="1857" heatid="2736" lane="2" />
                <RESULT eventid="1161" points="128" swimtime="00:00:44.10" resultid="1858" heatid="2846" lane="7" entrytime="00:00:43.87" entrycourse="LCM" />
                <RESULT eventid="1103" points="100" swimtime="00:01:46.33" resultid="1859" heatid="2778" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="136" swimtime="00:00:45.78" resultid="1860" heatid="2795" lane="1" entrytime="00:00:45.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Da Cunha Souza" birthdate="2015-05-30" gender="F" nation="BRA" license="400016" swrid="5652883" athleteid="2081" externalid="400016">
              <RESULTS>
                <RESULT eventid="1068" points="126" swimtime="00:03:44.58" resultid="2082" heatid="2737" lane="3" />
                <RESULT eventid="1164" points="150" reactiontime="+86" swimtime="00:00:50.51" resultid="2083" heatid="2851" lane="4" entrytime="00:00:55.78" entrycourse="LCM" />
                <RESULT eventid="1122" points="122" swimtime="00:01:44.00" resultid="2084" heatid="2798" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="152" swimtime="00:00:44.15" resultid="2085" heatid="2884" lane="5" entrytime="00:00:57.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Carcereri Navarro" birthdate="2013-12-19" gender="M" nation="BRA" license="376962" swrid="5588576" athleteid="3374" externalid="376962">
              <RESULTS>
                <RESULT eventid="1077" points="188" swimtime="00:00:45.24" resultid="3375" heatid="2750" lane="3" />
                <RESULT eventid="1103" points="148" swimtime="00:01:33.45" resultid="3376" heatid="2778" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="164" swimtime="00:00:40.67" resultid="3377" heatid="2846" lane="5" />
                <RESULT eventid="1211" points="193" swimtime="00:00:36.15" resultid="3378" heatid="2904" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Wolf Macedo" birthdate="2012-01-27" gender="F" nation="BRA" license="369277" swrid="5602592" athleteid="1722" externalid="369277">
              <RESULTS>
                <RESULT eventid="1074" points="303" swimtime="00:00:43.41" resultid="1723" heatid="2744" lane="1" />
                <RESULT eventid="1158" points="378" swimtime="00:00:33.76" resultid="1724" heatid="2843" lane="4" entrytime="00:00:35.45" entrycourse="LCM" />
                <RESULT eventid="1100" points="291" swimtime="00:01:23.68" resultid="1725" heatid="2777" lane="5" entrytime="00:01:24.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="365" swimtime="00:02:56.38" resultid="1726" heatid="2876" lane="3" entrytime="00:03:05.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                    <SPLIT distance="150" swimtime="00:02:18.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Baptistella" birthdate="2013-01-23" gender="M" nation="BRA" license="391152" swrid="5602545" athleteid="1996" externalid="391152">
              <RESULTS>
                <RESULT eventid="1089" points="184" swimtime="00:01:30.64" resultid="1997" heatid="2766" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1161" points="144" swimtime="00:00:42.48" resultid="1998" heatid="2845" lane="8" />
                <RESULT eventid="1119" points="189" swimtime="00:00:40.98" resultid="1999" heatid="2795" lane="5" entrytime="00:00:42.83" entrycourse="LCM" />
                <RESULT eventid="1195" status="DSQ" swimtime="00:03:19.14" resultid="2000" heatid="2877" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                    <SPLIT distance="100" swimtime="00:01:33.28" />
                    <SPLIT distance="150" swimtime="00:02:35.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcela" lastname="Tallao Benke" birthdate="2014-10-07" gender="F" nation="BRA" license="382075" swrid="5602586" athleteid="1891" externalid="382075">
              <RESULTS>
                <RESULT eventid="1068" points="265" swimtime="00:02:55.60" resultid="1892" heatid="2740" lane="3" entrytime="00:03:11.74" entrycourse="LCM" />
                <RESULT eventid="1080" points="218" swimtime="00:00:48.43" resultid="1893" heatid="2756" lane="3" entrytime="00:00:53.37" entrycourse="LCM" />
                <RESULT eventid="1152" points="268" swimtime="00:03:15.60" resultid="1894" heatid="2836" lane="4" entrytime="00:03:42.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                    <SPLIT distance="100" swimtime="00:01:32.85" />
                    <SPLIT distance="150" swimtime="00:02:33.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1106" points="206" swimtime="00:00:41.31" resultid="1895" heatid="2783" lane="5" entrytime="00:00:50.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Kraemer Geremia" birthdate="2013-08-16" gender="M" nation="BRA" license="377041" swrid="5588762" athleteid="1841" externalid="377041">
              <RESULTS>
                <RESULT eventid="1161" points="184" swimtime="00:00:39.11" resultid="1842" heatid="2847" lane="1" entrytime="00:00:40.35" entrycourse="LCM" />
                <RESULT eventid="1135" points="248" swimtime="00:01:14.54" resultid="1843" heatid="2820" lane="6" entrytime="00:01:18.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="218" swimtime="00:00:39.11" resultid="1844" heatid="2796" lane="8" entrytime="00:00:40.35" entrycourse="LCM" />
                <RESULT eventid="1211" points="256" swimtime="00:00:32.90" resultid="1845" heatid="2904" lane="5" entrytime="00:00:33.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Hadad" birthdate="2015-09-09" gender="M" nation="BRA" license="406740" swrid="5717272" athleteid="2096" externalid="406740">
              <RESULTS>
                <RESULT eventid="1071" points="73" swimtime="00:04:04.02" resultid="2097" heatid="2742" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.14" />
                    <SPLIT distance="150" swimtime="00:03:00.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="61" swimtime="00:01:05.79" resultid="2098" heatid="2759" lane="6" />
                <RESULT eventid="1167" points="50" reactiontime="+59" swimtime="00:01:03.66" resultid="2099" heatid="2855" lane="6" />
                <RESULT eventid="1125" points="67" swimtime="00:01:55.31" resultid="2100" heatid="2805" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Cavalca Petraglia" birthdate="2015-08-06" gender="M" nation="BRA" license="397275" swrid="5641757" athleteid="2061" externalid="397275">
              <RESULTS>
                <RESULT eventid="1083" points="74" swimtime="00:01:01.63" resultid="2062" heatid="2759" lane="2" />
                <RESULT eventid="1155" points="84" swimtime="00:04:19.44" resultid="2063" heatid="2838" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.46" />
                    <SPLIT distance="100" swimtime="00:02:06.87" />
                    <SPLIT distance="150" swimtime="00:03:24.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="43" swimtime="00:01:03.40" resultid="2064" heatid="2785" lane="1" />
                <RESULT eventid="1167" points="84" swimtime="00:00:53.65" resultid="2065" heatid="2855" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Da Cunha Souza" birthdate="2013-09-17" gender="M" nation="BRA" license="376975" swrid="5588618" athleteid="1806" externalid="376975">
              <RESULTS>
                <RESULT eventid="1065" points="173" swimtime="00:06:34.71" resultid="1807" heatid="2736" lane="8" />
                <RESULT eventid="1149" points="177" swimtime="00:03:01.63" resultid="1808" heatid="2832" lane="1" entrytime="00:03:16.75" entrycourse="LCM" />
                <RESULT eventid="1161" points="124" swimtime="00:00:44.64" resultid="1809" heatid="2846" lane="1" entrytime="00:00:46.90" entrycourse="LCM" />
                <RESULT eventid="1135" points="184" swimtime="00:01:22.34" resultid="1810" heatid="2819" lane="2" entrytime="00:01:32.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giuliana" lastname="Sovierzoski Ferreira" birthdate="2015-01-20" gender="F" nation="BRA" license="397168" swrid="5641776" athleteid="2056" externalid="397168">
              <RESULTS>
                <RESULT eventid="1080" points="165" swimtime="00:00:53.15" resultid="2057" heatid="2755" lane="4" entrytime="00:01:02.39" entrycourse="LCM" />
                <RESULT eventid="1152" points="85" swimtime="00:04:45.93" resultid="2058" heatid="2835" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:16.42" />
                    <SPLIT distance="100" swimtime="00:02:33.16" />
                    <SPLIT distance="150" swimtime="00:03:37.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="76" reactiontime="+76" swimtime="00:01:03.14" resultid="2059" heatid="2850" lane="5" />
                <RESULT eventid="1122" points="98" swimtime="00:01:52.05" resultid="2060" heatid="2799" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1182" points="204" swimtime="00:02:24.10" resultid="2232" heatid="2868" lane="4" entrytime="00:02:17.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:11.99" />
                    <SPLIT distance="150" swimtime="00:01:49.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1881" number="1" />
                    <RELAYPOSITION athleteid="1911" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2051" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1971" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1224" points="176" reactiontime="+70" swimtime="00:02:46.39" resultid="2238" heatid="2911" lane="4" entrytime="00:02:40.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.17" />
                    <SPLIT distance="100" swimtime="00:01:33.01" />
                    <SPLIT distance="150" swimtime="00:02:12.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2091" number="1" reactiontime="+70" />
                    <RELAYPOSITION athleteid="1911" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1881" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1971" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1188" points="249" swimtime="00:02:14.83" resultid="2233" heatid="2871" lane="4" entrytime="00:02:04.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                    <SPLIT distance="100" swimtime="00:01:08.20" />
                    <SPLIT distance="150" swimtime="00:01:41.62" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1821" number="1" />
                    <RELAYPOSITION athleteid="1841" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1747" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1856" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1230" points="206" reactiontime="+67" swimtime="00:02:37.71" resultid="2239" heatid="2914" lane="4" entrytime="00:02:24.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:01:23.33" />
                    <SPLIT distance="150" swimtime="00:02:04.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1996" number="1" reactiontime="+67" />
                    <RELAYPOSITION athleteid="1821" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1747" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1841" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="9" agemin="9" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1180" points="122" swimtime="00:02:50.73" resultid="2234" heatid="2867" lane="4" entrytime="00:02:33.64">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2026" number="1" />
                    <RELAYPOSITION athleteid="2011" number="2" />
                    <RELAYPOSITION athleteid="2071" number="3" />
                    <RELAYPOSITION athleteid="2061" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1222" points="131" swimtime="00:03:03.41" resultid="2237" heatid="2910" lane="4" entrytime="00:02:53.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.06" />
                    <SPLIT distance="150" swimtime="00:02:18.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2191" number="1" />
                    <RELAYPOSITION athleteid="2011" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2026" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2071" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1190" points="315" swimtime="00:02:04.65" resultid="2235" heatid="2873" lane="5" entrytime="00:02:00.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                    <SPLIT distance="100" swimtime="00:01:03.16" />
                    <SPLIT distance="150" swimtime="00:01:34.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1702" number="1" />
                    <RELAYPOSITION athleteid="1732" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1692" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1662" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1232" points="277" swimtime="00:02:23.05" resultid="2236" heatid="2916" lane="5" entrytime="00:02:17.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.26" />
                    <SPLIT distance="100" swimtime="00:01:17.70" />
                    <SPLIT distance="150" swimtime="00:01:53.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1662" number="1" />
                    <RELAYPOSITION athleteid="1727" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1732" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1702" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1182" points="150" swimtime="00:02:39.74" resultid="2256" heatid="2868" lane="5" entrytime="00:02:22.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.72" />
                    <SPLIT distance="100" swimtime="00:01:20.75" />
                    <SPLIT distance="150" swimtime="00:02:01.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2091" number="1" />
                    <RELAYPOSITION athleteid="1946" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1966" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2036" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1224" points="130" swimtime="00:03:03.95" resultid="2262" heatid="2911" lane="5" entrytime="00:02:49.65">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.83" />
                    <SPLIT distance="100" swimtime="00:01:42.06" />
                    <SPLIT distance="150" swimtime="00:02:26.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1946" number="1" />
                    <RELAYPOSITION athleteid="1926" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1966" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2051" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1188" points="224" swimtime="00:02:19.72" resultid="2257" heatid="2871" lane="5" entrytime="00:02:10.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                    <SPLIT distance="100" swimtime="00:01:07.58" />
                    <SPLIT distance="150" swimtime="00:01:43.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1816" number="1" />
                    <RELAYPOSITION athleteid="1836" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1791" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="3374" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1230" points="178" swimtime="00:02:45.50" resultid="2263" heatid="2914" lane="5" entrytime="00:02:31.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.03" />
                    <SPLIT distance="100" swimtime="00:01:30.82" />
                    <SPLIT distance="150" swimtime="00:02:09.82" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1856" number="1" />
                    <RELAYPOSITION athleteid="3374" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1836" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1816" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="9" agemin="9" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1180" points="77" swimtime="00:03:19.46" resultid="2258" heatid="2867" lane="5" entrytime="00:02:53.32">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2191" number="1" />
                    <RELAYPOSITION athleteid="2106" number="2" />
                    <RELAYPOSITION athleteid="2126" number="3" />
                    <RELAYPOSITION athleteid="2131" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1222" points="65" swimtime="00:03:51.05" resultid="2261" heatid="2910" lane="5" entrytime="00:03:20.00">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.55" />
                    <SPLIT distance="100" swimtime="00:02:01.03" />
                    <SPLIT distance="150" swimtime="00:02:59.48" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2106" number="1" />
                    <RELAYPOSITION athleteid="2146" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2061" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2116" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1190" points="283" swimtime="00:02:09.30" resultid="2259" heatid="2873" lane="3" entrytime="00:02:06.89">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.10" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1727" number="1" />
                    <RELAYPOSITION athleteid="1667" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1742" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1672" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1232" points="243" reactiontime="+72" swimtime="00:02:29.37" resultid="2260" heatid="2916" lane="3" entrytime="00:02:26.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1707" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="1871" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1692" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1667" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1182" points="86" swimtime="00:03:12.01" resultid="2280" heatid="2868" lane="6" entrytime="00:02:51.52">
                  <SPLITS>
                    <SPLIT distance="150" swimtime="00:02:20.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1921" number="1" />
                    <RELAYPOSITION athleteid="2196" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1926" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1951" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1224" points="66" swimtime="00:03:49.94" resultid="2286" heatid="2911" lane="6" entrytime="00:03:13.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.78" />
                    <SPLIT distance="100" swimtime="00:01:49.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2036" number="1" />
                    <RELAYPOSITION athleteid="2196" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1921" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1951" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1188" points="190" swimtime="00:02:27.62" resultid="2281" heatid="2871" lane="3" entrytime="00:02:21.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:15.12" />
                    <SPLIT distance="150" swimtime="00:01:54.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1806" number="1" />
                    <RELAYPOSITION athleteid="1861" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1851" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1996" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1230" points="129" reactiontime="+72" swimtime="00:03:04.51" resultid="2287" heatid="2914" lane="3" entrytime="00:02:39.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.73" />
                    <SPLIT distance="100" swimtime="00:01:39.29" />
                    <SPLIT distance="150" swimtime="00:02:26.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1791" number="1" reactiontime="+72" />
                    <RELAYPOSITION athleteid="1851" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1806" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1861" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="9" agemin="9" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1180" points="57" swimtime="00:03:40.60" resultid="2282" heatid="2867" lane="3" entrytime="00:03:03.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.97" />
                    <SPLIT distance="100" swimtime="00:01:50.38" />
                    <SPLIT distance="150" swimtime="00:02:48.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2171" number="1" />
                    <RELAYPOSITION athleteid="2096" number="2" />
                    <RELAYPOSITION athleteid="2146" number="3" />
                    <RELAYPOSITION athleteid="2116" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1222" points="33" reactiontime="+62" swimtime="00:04:49.34" resultid="2285" heatid="2910" lane="3" entrytime="00:03:35.15">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2096" number="1" reactiontime="+62" />
                    <RELAYPOSITION athleteid="2171" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2126" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2151" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1190" points="241" swimtime="00:02:16.24" resultid="2283" heatid="2873" lane="7" entrytime="00:02:13.06">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                    <SPLIT distance="150" swimtime="00:01:43.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1707" number="1" />
                    <RELAYPOSITION athleteid="1871" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1697" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1846" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1232" points="189" reactiontime="+68" swimtime="00:02:42.39" resultid="2284" heatid="2916" lane="7" entrytime="00:02:38.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                    <SPLIT distance="100" swimtime="00:01:29.50" />
                    <SPLIT distance="150" swimtime="00:02:06.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1742" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="1697" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1672" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1846" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1178" points="206" swimtime="00:02:41.16" resultid="2224" heatid="2866" lane="4" entrytime="00:02:21.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1891" number="1" />
                    <RELAYPOSITION athleteid="2006" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1956" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1976" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1220" points="192" reactiontime="+79" swimtime="00:03:02.98" resultid="2230" heatid="2909" lane="4" entrytime="00:02:46.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.25" />
                    <SPLIT distance="100" swimtime="00:01:36.26" />
                    <SPLIT distance="150" swimtime="00:02:23.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2046" number="1" reactiontime="+79" />
                    <RELAYPOSITION athleteid="1891" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1956" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1976" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1184" points="336" swimtime="00:02:17.08" resultid="2225" heatid="2869" lane="4" entrytime="00:02:07.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                    <SPLIT distance="100" swimtime="00:01:07.63" />
                    <SPLIT distance="150" swimtime="00:01:42.68" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2156" number="1" />
                    <RELAYPOSITION athleteid="1767" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1757" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1752" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1226" points="305" reactiontime="+73" swimtime="00:02:36.74" resultid="2228" heatid="2912" lane="4" entrytime="00:02:24.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                    <SPLIT distance="100" swimtime="00:01:23.15" />
                    <SPLIT distance="150" swimtime="00:02:03.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1801" number="1" reactiontime="+73" />
                    <RELAYPOSITION athleteid="2156" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1757" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1752" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="9" agemin="9" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1176" points="167" swimtime="00:02:52.85" resultid="2226" heatid="2865" lane="4" entrytime="00:02:51.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.64" />
                    <SPLIT distance="100" swimtime="00:01:27.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2066" number="1" />
                    <RELAYPOSITION athleteid="2081" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2041" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2086" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1218" points="137" reactiontime="+69" swimtime="00:03:24.74" resultid="2229" heatid="2908" lane="4" entrytime="00:03:30.32">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.48" />
                    <SPLIT distance="100" swimtime="00:01:44.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2066" number="1" reactiontime="+69" />
                    <RELAYPOSITION athleteid="2056" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2041" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2081" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1186" points="466" swimtime="00:02:02.95" resultid="2227" heatid="2870" lane="4" entrytime="00:02:01.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.48" />
                    <SPLIT distance="150" swimtime="00:01:32.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1831" number="1" />
                    <RELAYPOSITION athleteid="1682" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1762" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1677" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1228" points="448" reactiontime="+68" swimtime="00:02:17.93" resultid="2231" heatid="2913" lane="4" entrytime="00:02:18.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:14.65" />
                    <SPLIT distance="150" swimtime="00:01:47.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1677" number="1" reactiontime="+68" />
                    <RELAYPOSITION athleteid="1712" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1831" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1682" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1178" status="DSQ" swimtime="00:02:52.63" resultid="2248" heatid="2866" lane="3" entrytime="00:02:41.62">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.90" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1991" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="1896" number="2" reactiontime="+3276" status="DSQ" />
                    <RELAYPOSITION athleteid="2046" number="3" reactiontime="+3276" status="DSQ" />
                    <RELAYPOSITION athleteid="2001" number="4" reactiontime="+3276" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1220" points="149" swimtime="00:03:18.84" resultid="2254" heatid="2909" lane="5" entrytime="00:03:00.61">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.58" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2006" number="1" />
                    <RELAYPOSITION athleteid="2001" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1896" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1991" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1184" points="315" swimtime="00:02:20.00" resultid="2249" heatid="2869" lane="5" entrytime="00:02:09.96">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.27" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1811" number="1" />
                    <RELAYPOSITION athleteid="1866" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1796" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1801" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1226" points="258" swimtime="00:02:45.75" resultid="2252" heatid="2912" lane="5" entrytime="00:02:33.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                    <SPLIT distance="100" swimtime="00:01:30.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1866" number="1" />
                    <RELAYPOSITION athleteid="1916" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1796" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1767" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="9" agemin="9" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1176" points="116" swimtime="00:03:15.04" resultid="2250" heatid="2865" lane="3" entrytime="00:03:22.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.37" />
                    <SPLIT distance="100" swimtime="00:01:30.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2121" number="1" />
                    <RELAYPOSITION athleteid="2021" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2136" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2101" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1218" points="116" swimtime="00:03:36.13" resultid="2253" heatid="2908" lane="5" entrytime="00:03:41.43">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:52.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2101" number="1" />
                    <RELAYPOSITION athleteid="2021" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2086" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2121" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1186" points="446" swimtime="00:02:04.69" resultid="2251" heatid="2870" lane="5" entrytime="00:02:19.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                    <SPLIT distance="100" swimtime="00:01:00.78" />
                    <SPLIT distance="150" swimtime="00:01:32.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1772" number="1" />
                    <RELAYPOSITION athleteid="1717" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1981" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1722" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1228" points="389" swimtime="00:02:24.55" resultid="2255" heatid="2913" lane="5" entrytime="00:02:42.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                    <SPLIT distance="100" swimtime="00:01:19.97" />
                    <SPLIT distance="150" swimtime="00:01:54.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1981" number="1" />
                    <RELAYPOSITION athleteid="1737" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1722" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1772" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1178" status="WDR" swimtime="00:00:00.00" resultid="2272" heatid="2866" lane="6" entrytime="00:02:52.13">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="2" reactiontime="0" />
                    <RELAYPOSITION number="3" reactiontime="0" />
                    <RELAYPOSITION number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1220" status="WDR" swimtime="00:00:00.00" resultid="2278" heatid="2909" lane="6" entrytime="00:03:21.59">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION number="2" reactiontime="0" />
                    <RELAYPOSITION number="3" reactiontime="0" />
                    <RELAYPOSITION number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1184" points="210" swimtime="00:02:40.25" resultid="2273" heatid="2869" lane="3" entrytime="00:02:24.37">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1886" number="1" />
                    <RELAYPOSITION athleteid="1986" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1936" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1916" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1226" points="197" reactiontime="+51" swimtime="00:03:01.44" resultid="2276" heatid="2912" lane="6" entrytime="00:02:49.86">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.54" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1811" number="1" reactiontime="+51" />
                    <RELAYPOSITION athleteid="1786" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1936" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1886" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="9" agemin="9" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1176" points="83" swimtime="00:03:37.71" resultid="2274" heatid="2865" lane="5" entrytime="00:03:17.47">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2056" number="1" />
                    <RELAYPOSITION athleteid="2076" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2166" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2111" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1218" points="85" swimtime="00:03:59.43" resultid="2277" heatid="2908" lane="3" entrytime="00:04:06.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.69" />
                    <SPLIT distance="100" swimtime="00:02:07.96" />
                    <SPLIT distance="150" swimtime="00:03:03.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2111" number="1" />
                    <RELAYPOSITION athleteid="2031" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2076" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="2186" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1186" points="335" swimtime="00:02:17.18" resultid="2275" heatid="2870" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:05.99" />
                    <SPLIT distance="150" swimtime="00:01:38.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1737" number="1" />
                    <RELAYPOSITION athleteid="2141" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1712" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1876" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1228" points="286" reactiontime="+65" swimtime="00:02:40.27" resultid="2279" heatid="2913" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                    <SPLIT distance="100" swimtime="00:01:23.29" />
                    <SPLIT distance="150" swimtime="00:02:00.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1762" number="1" reactiontime="+65" />
                    <RELAYPOSITION athleteid="2141" number="2" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1717" number="3" reactiontime="+3276" />
                    <RELAYPOSITION athleteid="1876" number="4" reactiontime="+3276" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1096" swimtime="00:02:14.00" resultid="2240" heatid="2772" lane="4" entrytime="00:02:03.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                    <SPLIT distance="100" swimtime="00:01:07.27" />
                    <SPLIT distance="150" swimtime="00:01:41.06" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1841" number="1" />
                    <RELAYPOSITION athleteid="1747" number="2" />
                    <RELAYPOSITION athleteid="1752" number="3" />
                    <RELAYPOSITION athleteid="2156" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1142" swimtime="00:02:36.27" resultid="2247" heatid="2825" lane="4" entrytime="00:02:23.59">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1801" number="1" />
                    <RELAYPOSITION athleteid="1821" number="2" />
                    <RELAYPOSITION athleteid="1757" number="3" />
                    <RELAYPOSITION athleteid="1841" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1098" swimtime="00:02:01.82" resultid="2241" heatid="2774" lane="4" entrytime="00:02:00.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.35" />
                    <SPLIT distance="100" swimtime="00:01:01.09" />
                    <SPLIT distance="150" swimtime="00:01:31.76" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1831" number="1" />
                    <RELAYPOSITION athleteid="1662" number="2" />
                    <RELAYPOSITION athleteid="1677" number="3" />
                    <RELAYPOSITION athleteid="1702" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1144" swimtime="00:02:17.60" resultid="2244" heatid="2827" lane="4" entrytime="00:02:16.15">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1831" number="1" />
                    <RELAYPOSITION athleteid="1712" number="2" />
                    <RELAYPOSITION athleteid="1662" number="3" />
                    <RELAYPOSITION athleteid="1702" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="9" agemin="9" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1092" swimtime="00:02:45.81" resultid="2242" heatid="2769" lane="4" entrytime="00:03:00.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                    <SPLIT distance="100" swimtime="00:01:19.15" />
                    <SPLIT distance="150" swimtime="00:02:02.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2026" number="1" />
                    <RELAYPOSITION athleteid="2011" number="2" />
                    <RELAYPOSITION athleteid="2066" number="3" />
                    <RELAYPOSITION athleteid="2081" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1138" swimtime="00:03:06.28" resultid="2246" heatid="2822" lane="4" entrytime="00:03:00.99">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2066" number="1" />
                    <RELAYPOSITION athleteid="2011" number="2" />
                    <RELAYPOSITION athleteid="2026" number="3" />
                    <RELAYPOSITION athleteid="2081" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1094" swimtime="00:02:27.03" resultid="2243" heatid="2771" lane="4" entrytime="00:02:19.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                    <SPLIT distance="100" swimtime="00:01:12.10" />
                    <SPLIT distance="150" swimtime="00:01:52.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1881" number="1" />
                    <RELAYPOSITION athleteid="1891" number="2" />
                    <RELAYPOSITION athleteid="1956" number="3" />
                    <RELAYPOSITION athleteid="1971" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1140" swimtime="00:02:50.15" resultid="2245" heatid="2824" lane="4" entrytime="00:02:42.47">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1891" number="1" />
                    <RELAYPOSITION athleteid="1911" number="2" />
                    <RELAYPOSITION athleteid="1881" number="3" />
                    <RELAYPOSITION athleteid="1976" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1096" swimtime="00:02:16.75" resultid="2264" heatid="2772" lane="3" entrytime="00:02:08.55">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.99" />
                    <SPLIT distance="150" swimtime="00:01:43.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1767" number="1" />
                    <RELAYPOSITION athleteid="1757" number="2" />
                    <RELAYPOSITION athleteid="1856" number="3" />
                    <RELAYPOSITION athleteid="1821" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1142" swimtime="00:02:34.63" resultid="2271" heatid="2825" lane="5" entrytime="00:02:25.54">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1752" number="1" />
                    <RELAYPOSITION athleteid="2156" number="2" />
                    <RELAYPOSITION athleteid="1747" number="3" />
                    <RELAYPOSITION athleteid="1856" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1098" swimtime="00:02:05.98" resultid="2265" heatid="2774" lane="5" entrytime="00:02:04.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                    <SPLIT distance="100" swimtime="00:01:01.72" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1682" number="1" />
                    <RELAYPOSITION athleteid="1692" number="2" />
                    <RELAYPOSITION athleteid="1732" number="3" />
                    <RELAYPOSITION athleteid="1762" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1144" swimtime="00:02:23.38" resultid="2268" heatid="2827" lane="5" entrytime="00:02:23.70">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1677" number="1" />
                    <RELAYPOSITION athleteid="1727" number="2" />
                    <RELAYPOSITION athleteid="1732" number="3" />
                    <RELAYPOSITION athleteid="1682" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="9" agemin="9" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1092" swimtime="00:03:00.24" resultid="2266" heatid="2769" lane="5" entrytime="00:03:20.55">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2071" number="1" />
                    <RELAYPOSITION athleteid="2041" number="2" />
                    <RELAYPOSITION athleteid="2086" number="3" />
                    <RELAYPOSITION athleteid="2061" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1138" swimtime="00:03:23.72" resultid="2270" heatid="2822" lane="5" entrytime="00:03:20.55">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2061" number="1" />
                    <RELAYPOSITION athleteid="2056" number="2" />
                    <RELAYPOSITION athleteid="2041" number="3" />
                    <RELAYPOSITION athleteid="2071" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1094" swimtime="00:02:39.12" resultid="2267" heatid="2771" lane="5" entrytime="00:02:19.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                    <SPLIT distance="100" swimtime="00:01:17.38" />
                    <SPLIT distance="150" swimtime="00:01:59.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1911" number="1" />
                    <RELAYPOSITION athleteid="2091" number="2" />
                    <RELAYPOSITION athleteid="1991" number="3" />
                    <RELAYPOSITION athleteid="1976" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1140" swimtime="00:02:58.68" resultid="2269" heatid="2824" lane="6" entrytime="00:02:51.40">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2091" number="1" />
                    <RELAYPOSITION athleteid="2001" number="2" />
                    <RELAYPOSITION athleteid="1971" number="3" />
                    <RELAYPOSITION athleteid="1956" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="11" agemin="11" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1096" swimtime="00:02:15.55" resultid="2288" heatid="2772" lane="5" entrytime="00:02:07.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="100" swimtime="00:01:08.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1801" number="1" />
                    <RELAYPOSITION athleteid="1866" number="2" />
                    <RELAYPOSITION athleteid="1816" number="3" />
                    <RELAYPOSITION athleteid="1836" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1142" swimtime="00:02:39.61" resultid="2295" heatid="2825" lane="3" entrytime="00:02:29.62">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1796" number="1" />
                    <RELAYPOSITION athleteid="3374" number="2" />
                    <RELAYPOSITION athleteid="1836" number="3" />
                    <RELAYPOSITION athleteid="1767" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="12" agemin="12" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1098" swimtime="00:02:06.28" resultid="2289" heatid="2774" lane="6" entrytime="00:02:10.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:04.18" />
                    <SPLIT distance="150" swimtime="00:01:36.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1722" number="1" />
                    <RELAYPOSITION athleteid="1727" number="2" />
                    <RELAYPOSITION athleteid="1667" number="3" />
                    <RELAYPOSITION athleteid="1772" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1144" swimtime="00:02:23.85" resultid="2292" heatid="2827" lane="6" entrytime="00:02:33.25">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1981" number="1" />
                    <RELAYPOSITION athleteid="1871" number="2" />
                    <RELAYPOSITION athleteid="1722" number="3" />
                    <RELAYPOSITION athleteid="1692" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="9" agemin="9" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1092" swimtime="00:03:03.08" resultid="2290" heatid="2769" lane="3" entrytime="00:03:27.10">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.48" />
                    <SPLIT distance="150" swimtime="00:02:15.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2021" number="1" />
                    <RELAYPOSITION athleteid="2121" number="2" />
                    <RELAYPOSITION athleteid="2191" number="3" />
                    <RELAYPOSITION athleteid="2106" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1138" swimtime="00:03:33.65" resultid="2294" heatid="2822" lane="3" entrytime="00:03:27.10">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2021" number="1" />
                    <RELAYPOSITION athleteid="2131" number="2" />
                    <RELAYPOSITION athleteid="2086" number="3" />
                    <RELAYPOSITION athleteid="2191" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;C&quot;" number="3">
              <RESULTS>
                <RESULT eventid="1094" swimtime="00:02:45.19" resultid="2291" heatid="2771" lane="6" entrytime="00:02:28.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.80" />
                    <SPLIT distance="100" swimtime="00:01:17.06" />
                    <SPLIT distance="150" swimtime="00:02:02.70" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1906" number="1" />
                    <RELAYPOSITION athleteid="2051" number="2" />
                    <RELAYPOSITION athleteid="1896" number="3" />
                    <RELAYPOSITION athleteid="2006" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1140" swimtime="00:03:14.19" resultid="2293" heatid="2824" lane="3" entrytime="00:02:45.31">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1906" number="1" />
                    <RELAYPOSITION athleteid="2006" number="2" />
                    <RELAYPOSITION athleteid="1966" number="3" />
                    <RELAYPOSITION athleteid="1991" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="2864" nation="BRA" region="PR" clubid="1234" swrid="93756" name="Associacao De Pais E Amigos Da Natacao De Ponta Gr" shortname="Apan Ponta Grossa">
          <ATHLETES>
            <ATHLETE firstname="Gustavo" lastname="Hilgenberg Lievore" birthdate="2014-04-23" gender="M" nation="BRA" license="391167" swrid="5602546" athleteid="1255" externalid="391167">
              <RESULTS>
                <RESULT eventid="1083" points="135" swimtime="00:00:50.51" resultid="1256" heatid="2762" lane="6" entrytime="00:00:53.35" entrycourse="LCM" />
                <RESULT eventid="1109" points="105" swimtime="00:00:47.20" resultid="1257" heatid="2784" lane="4" />
                <RESULT eventid="1167" points="160" reactiontime="+73" swimtime="00:00:43.29" resultid="1258" heatid="2858" lane="3" entrytime="00:00:46.05" entrycourse="LCM" />
                <RESULT eventid="1205" points="182" swimtime="00:00:36.84" resultid="1259" heatid="2893" lane="2" entrytime="00:00:38.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Bischof Rogoski" birthdate="2014-10-03" gender="M" nation="BRA" license="401860" swrid="5661341" athleteid="1270" externalid="401860">
              <RESULTS>
                <RESULT eventid="1083" points="103" swimtime="00:00:55.28" resultid="1271" heatid="2761" lane="6" entrytime="00:01:02.75" entrycourse="LCM" />
                <RESULT eventid="1167" points="125" reactiontime="+64" swimtime="00:00:47.01" resultid="1272" heatid="2857" lane="5" entrytime="00:00:52.87" entrycourse="LCM" />
                <RESULT eventid="1125" points="147" swimtime="00:01:28.73" resultid="1273" heatid="2807" lane="3" entrytime="00:01:43.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="180" swimtime="00:00:36.97" resultid="1274" heatid="2892" lane="3" entrytime="00:00:42.41" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Victoria Borges" birthdate="2014-01-16" gender="F" nation="BRA" license="376737" swrid="5602587" athleteid="1240" externalid="376737">
              <RESULTS>
                <RESULT eventid="1068" points="143" swimtime="00:03:35.55" resultid="1241" heatid="2738" lane="6" />
                <RESULT eventid="1164" points="166" reactiontime="+74" swimtime="00:00:48.84" resultid="1242" heatid="2852" lane="6" entrytime="00:00:51.16" entrycourse="LCM" />
                <RESULT eventid="1122" points="161" swimtime="00:01:34.92" resultid="1243" heatid="2800" lane="4" entrytime="00:01:46.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="198" swimtime="00:00:40.50" resultid="1244" heatid="2886" lane="7" entrytime="00:00:44.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolly" lastname="Victoria Souza" birthdate="2015-11-15" gender="F" nation="BRA" license="400091" swrid="5652902" athleteid="1265" externalid="400091">
              <RESULTS>
                <RESULT eventid="1080" points="127" swimtime="00:00:57.94" resultid="1266" heatid="2755" lane="1" entrytime="00:01:05.78" entrycourse="LCM" />
                <RESULT eventid="1164" points="112" swimtime="00:00:55.70" resultid="1267" heatid="2851" lane="7" entrytime="00:01:02.94" entrycourse="LCM" />
                <RESULT eventid="1122" points="99" swimtime="00:01:51.62" resultid="1268" heatid="2799" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1202" points="143" swimtime="00:00:45.09" resultid="1269" heatid="2885" lane="7" entrytime="00:00:50.27" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariana" lastname="Brunetti Silva" birthdate="2014-03-24" gender="F" nation="BRA" license="390878" swrid="5602517" athleteid="1250" externalid="390878">
              <RESULTS>
                <RESULT eventid="1080" points="149" swimtime="00:00:54.91" resultid="1251" heatid="2755" lane="5" entrytime="00:01:02.46" entrycourse="LCM" />
                <RESULT eventid="1106" points="96" swimtime="00:00:53.21" resultid="1252" heatid="2782" lane="5" entrytime="00:01:04.40" entrycourse="LCM" />
                <RESULT eventid="1164" points="153" reactiontime="+76" swimtime="00:00:50.19" resultid="1253" heatid="2852" lane="1" entrytime="00:00:52.40" entrycourse="LCM" />
                <RESULT eventid="1202" points="195" swimtime="00:00:40.65" resultid="1254" heatid="2885" lane="3" entrytime="00:00:46.62" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Campagnoli" birthdate="2013-03-13" gender="M" nation="BRA" license="370651" swrid="5602519" athleteid="1235" externalid="370651">
              <RESULTS>
                <RESULT eventid="1089" points="240" swimtime="00:01:22.97" resultid="1236" heatid="2767" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="268" swimtime="00:01:12.68" resultid="1237" heatid="2821" lane="3" entrytime="00:01:10.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="219" swimtime="00:01:21.92" resultid="1238" heatid="2778" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1211" points="280" swimtime="00:00:31.93" resultid="1239" heatid="2905" lane="4" entrytime="00:00:31.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Clara Domingues" birthdate="2012-01-19" gender="F" nation="BRA" license="377291" swrid="5588599" athleteid="1245" externalid="377291">
              <RESULTS>
                <RESULT eventid="1062" status="DSQ" swimtime="00:06:36.77" resultid="1246" heatid="2733" lane="6" />
                <RESULT eventid="1086" points="165" swimtime="00:01:44.52" resultid="1247" heatid="2765" lane="8" entrytime="00:01:48.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1146" points="222" swimtime="00:03:06.23" resultid="1248" heatid="2828" lane="4" entrytime="00:03:19.08" entrycourse="LCM" />
                <RESULT eventid="1132" points="206" swimtime="00:01:27.48" resultid="1249" heatid="2814" lane="1" entrytime="00:01:28.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Clara Rigailo" birthdate="2013-04-06" gender="F" nation="BRA" license="396828" swrid="5641758" athleteid="1260" externalid="396828">
              <RESULTS>
                <RESULT eventid="1074" points="283" swimtime="00:00:44.40" resultid="1261" heatid="2746" lane="4" entrytime="00:00:49.89" entrycourse="LCM" />
                <RESULT eventid="1116" points="187" swimtime="00:00:46.91" resultid="1262" heatid="2790" lane="3" entrytime="00:00:48.89" entrycourse="LCM" />
                <RESULT eventid="1170" points="295" swimtime="00:01:36.33" resultid="1263" heatid="2860" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="236" swimtime="00:00:38.17" resultid="1264" heatid="2897" lane="8" entrytime="00:00:42.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="10" agemin="10" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/PONTA GROSSA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1094" swimtime="00:02:36.36" resultid="1275" heatid="2770" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.32" />
                    <SPLIT distance="100" swimtime="00:01:18.10" />
                    <SPLIT distance="150" swimtime="00:01:59.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1255" number="1" />
                    <RELAYPOSITION athleteid="1240" number="2" />
                    <RELAYPOSITION athleteid="1250" number="3" />
                    <RELAYPOSITION athleteid="1270" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1140" swimtime="00:03:10.99" resultid="1276" heatid="2824" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1240" number="1" />
                    <RELAYPOSITION athleteid="1250" number="2" />
                    <RELAYPOSITION athleteid="1255" number="3" />
                    <RELAYPOSITION athleteid="1270" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="18151" nation="BRA" region="PR" clubid="1585" swrid="95180" name="Clube Uniao Recreativo Palmense" shortname="Clube União">
          <ATHLETES>
            <ATHLETE firstname="Pedro" lastname="Durli Giusti" birthdate="2012-11-06" gender="M" nation="BRA" license="408512" swrid="5725990" athleteid="1592" externalid="408512">
              <RESULTS>
                <RESULT eventid="1161" points="91" swimtime="00:00:49.49" resultid="1593" heatid="2845" lane="1" />
                <RESULT eventid="1135" points="153" swimtime="00:01:27.48" resultid="1594" heatid="2816" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="134" swimtime="00:00:45.98" resultid="1595" heatid="2793" lane="7" />
                <RESULT eventid="1211" points="173" swimtime="00:00:37.46" resultid="1596" heatid="2901" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Durli Giusti" birthdate="2015-07-05" gender="M" nation="BRA" license="408516" swrid="5725989" athleteid="1597" externalid="408516">
              <RESULTS>
                <RESULT eventid="1109" points="59" swimtime="00:00:57.11" resultid="1598" heatid="2785" lane="2" />
                <RESULT eventid="1167" points="117" reactiontime="+62" swimtime="00:00:48.10" resultid="1599" heatid="2854" lane="6" />
                <RESULT eventid="1205" points="140" swimtime="00:00:40.19" resultid="1600" heatid="2890" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Langaro Spaniol" birthdate="2013-06-18" gender="F" nation="BRA" license="406600" swrid="5074027" athleteid="1586" externalid="406600">
              <RESULTS>
                <RESULT eventid="1074" points="294" swimtime="00:00:43.84" resultid="1587" heatid="2744" lane="6" />
                <RESULT eventid="1158" points="213" swimtime="00:00:40.90" resultid="1588" heatid="2841" lane="5" />
                <RESULT eventid="1132" points="291" swimtime="00:01:17.98" resultid="1589" heatid="2811" lane="4" />
                <RESULT eventid="1170" points="257" swimtime="00:01:40.74" resultid="1590" heatid="3396" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="326" swimtime="00:00:34.29" resultid="1591" heatid="2895" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
