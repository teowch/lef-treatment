<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.80168">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Curitiba" name="Torneio Regional da 1ª Região (Infantil/Sênior)" course="LCM" deadline="2024-10-08" entrystartdate="2024-09-30" entrytype="INVITATION" hostclub="Clube Curitibano" hostclub.url="https://clubecuritibano.com.br/" number="38316" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/newInterface/eventos/38316" startmethod="1" timing="AUTOMATIC" touchpad="ONESIDE" masters="F" withdrawuntil="2024-10-09" state="PR" nation="BRA" hytek.courseorder="L">
      <AGEDATE value="2024-01-01" type="YEAR" />
      <POOL name="Parque Aquático do Clube Curitibano" lanemin="1" lanemax="8" />
      <FACILITY city="Curitiba" name="Parque Aquático do Clube Curitibano" nation="BRA" state="PR" street="Avenida Presidente Getúlio Vargas, 2857" street2="Água Verde" zip="80240-040" />
      <POINTTABLE pointtableid="3017" name="AQUA Point Scoring" version="2024" />
      <QUALIFY from="2023-10-12" until="2024-10-11" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-10-12" daytime="09:10" endtime="12:26" number="1" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1060" daytime="09:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1616" />
                    <RANKING order="2" place="2" resultid="1698" />
                    <RANKING order="3" place="3" resultid="1694" />
                    <RANKING order="4" place="4" resultid="1255" />
                    <RANKING order="5" place="5" resultid="1612" />
                    <RANKING order="6" place="6" resultid="1654" />
                    <RANKING order="7" place="7" resultid="1728" />
                    <RANKING order="8" place="8" resultid="1764" />
                    <RANKING order="9" place="9" resultid="1412" />
                    <RANKING order="10" place="10" resultid="1380" />
                    <RANKING order="11" place="11" resultid="1793" />
                    <RANKING order="12" place="12" resultid="1305" />
                    <RANKING order="13" place="13" resultid="2008" />
                    <RANKING order="14" place="14" resultid="1277" />
                    <RANKING order="15" place="15" resultid="1289" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1546" />
                    <RANKING order="2" place="2" resultid="1550" />
                    <RANKING order="3" place="3" resultid="1280" />
                    <RANKING order="4" place="4" resultid="1681" />
                    <RANKING order="5" place="5" resultid="1990" />
                    <RANKING order="6" place="6" resultid="1471" />
                    <RANKING order="7" place="7" resultid="2016" />
                    <RANKING order="8" place="8" resultid="1542" />
                    <RANKING order="9" place="9" resultid="1562" />
                    <RANKING order="10" place="10" resultid="1441" />
                    <RANKING order="11" place="11" resultid="1259" />
                    <RANKING order="12" place="12" resultid="1783" />
                    <RANKING order="13" place="13" resultid="1879" />
                    <RANKING order="14" place="14" resultid="1252" />
                    <RANKING order="15" place="15" resultid="1910" />
                    <RANKING order="16" place="16" resultid="1245" />
                    <RANKING order="17" place="-1" resultid="1298" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1063" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1518" />
                    <RANKING order="2" place="2" resultid="1768" />
                    <RANKING order="3" place="3" resultid="1350" />
                    <RANKING order="4" place="4" resultid="1508" />
                    <RANKING order="5" place="5" resultid="1945" />
                    <RANKING order="6" place="6" resultid="1511" />
                    <RANKING order="7" place="7" resultid="1953" />
                    <RANKING order="8" place="8" resultid="1401" />
                    <RANKING order="9" place="9" resultid="1895" />
                    <RANKING order="10" place="10" resultid="1438" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1891" />
                    <RANKING order="2" place="2" resultid="1272" />
                    <RANKING order="3" place="3" resultid="1658" />
                    <RANKING order="4" place="4" resultid="1859" />
                    <RANKING order="5" place="5" resultid="1374" />
                    <RANKING order="6" place="6" resultid="1805" />
                    <RANKING order="7" place="7" resultid="1284" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1482" />
                    <RANKING order="2" place="2" resultid="1362" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1067" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1823" />
                    <RANKING order="2" place="2" resultid="1827" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2312" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2313" daytime="09:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2314" daytime="09:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2315" daytime="09:18" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2316" daytime="09:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2317" daytime="09:22" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2318" daytime="09:24" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1068" daytime="09:26" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1069" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1646" />
                    <RANKING order="2" place="2" resultid="1620" />
                    <RANKING order="3" place="3" resultid="1249" />
                    <RANKING order="4" place="4" resultid="1590" />
                    <RANKING order="5" place="5" resultid="1294" />
                    <RANKING order="6" place="6" resultid="1417" />
                    <RANKING order="7" place="7" resultid="1960" />
                    <RANKING order="8" place="8" resultid="1582" />
                    <RANKING order="9" place="9" resultid="2003" />
                    <RANKING order="10" place="10" resultid="1586" />
                    <RANKING order="11" place="11" resultid="1633" />
                    <RANKING order="12" place="12" resultid="1675" />
                    <RANKING order="13" place="13" resultid="1870" />
                    <RANKING order="14" place="14" resultid="1358" />
                    <RANKING order="15" place="15" resultid="1301" />
                    <RANKING order="16" place="16" resultid="1261" />
                    <RANKING order="17" place="17" resultid="1428" />
                    <RANKING order="18" place="18" resultid="1600" />
                    <RANKING order="19" place="19" resultid="2005" />
                    <RANKING order="20" place="20" resultid="1788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1445" />
                    <RANKING order="2" place="2" resultid="1689" />
                    <RANKING order="3" place="3" resultid="1555" />
                    <RANKING order="4" place="4" resultid="1575" />
                    <RANKING order="5" place="5" resultid="1567" />
                    <RANKING order="6" place="6" resultid="2024" />
                    <RANKING order="7" place="7" resultid="1535" />
                    <RANKING order="8" place="8" resultid="1571" />
                    <RANKING order="9" place="9" resultid="1907" />
                    <RANKING order="10" place="10" resultid="1353" />
                    <RANKING order="11" place="11" resultid="1391" />
                    <RANKING order="12" place="12" resultid="1761" />
                    <RANKING order="13" place="13" resultid="1368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1223" />
                    <RANKING order="2" place="2" resultid="1478" />
                    <RANKING order="3" place="3" resultid="1344" />
                    <RANKING order="4" place="4" resultid="1938" />
                    <RANKING order="5" place="5" resultid="1811" />
                    <RANKING order="6" place="6" resultid="1947" />
                    <RANKING order="7" place="7" resultid="2013" />
                    <RANKING order="8" place="8" resultid="1856" />
                    <RANKING order="9" place="9" resultid="1733" />
                    <RANKING order="10" place="10" resultid="1384" />
                    <RANKING order="11" place="11" resultid="1522" />
                    <RANKING order="12" place="12" resultid="1422" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1702" />
                    <RANKING order="2" place="2" resultid="1641" />
                    <RANKING order="3" place="3" resultid="1678" />
                    <RANKING order="4" place="4" resultid="1943" />
                    <RANKING order="5" place="5" resultid="1499" />
                    <RANKING order="6" place="6" resultid="1528" />
                    <RANKING order="7" place="7" resultid="1929" />
                    <RANKING order="8" place="8" resultid="1377" />
                    <RANKING order="9" place="9" resultid="1743" />
                    <RANKING order="10" place="10" resultid="1914" />
                    <RANKING order="11" place="11" resultid="1315" />
                    <RANKING order="12" place="12" resultid="1371" />
                    <RANKING order="13" place="13" resultid="1397" />
                    <RANKING order="14" place="14" resultid="1738" />
                    <RANKING order="15" place="15" resultid="1758" />
                    <RANKING order="16" place="16" resultid="1819" />
                    <RANKING order="17" place="17" resultid="1310" />
                    <RANKING order="18" place="-1" resultid="1431" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1923" />
                    <RANKING order="2" place="2" resultid="1887" />
                    <RANKING order="3" place="3" resultid="1798" />
                    <RANKING order="4" place="4" resultid="1774" />
                    <RANKING order="5" place="5" resultid="1748" />
                    <RANKING order="6" place="6" resultid="1829" />
                    <RANKING order="7" place="7" resultid="1779" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1458" />
                    <RANKING order="2" place="2" resultid="1951" />
                    <RANKING order="3" place="3" resultid="1847" />
                    <RANKING order="4" place="4" resultid="1327" />
                    <RANKING order="5" place="5" resultid="1408" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1685" />
                    <RANKING order="2" place="2" resultid="1336" />
                    <RANKING order="3" place="3" resultid="1850" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2319" daytime="09:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2320" daytime="09:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2321" daytime="09:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2322" daytime="09:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2323" daytime="09:36" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2324" daytime="09:38" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2325" daytime="09:40" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="2326" daytime="09:42" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="2327" daytime="09:44" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="2328" daytime="09:46" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1076" daytime="09:48" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1077" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1598" />
                    <RANKING order="2" place="2" resultid="1984" />
                    <RANKING order="3" place="3" resultid="1957" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1472" />
                    <RANKING order="2" place="2" resultid="1995" />
                    <RANKING order="3" place="-1" resultid="1991" />
                    <RANKING order="4" place="-1" resultid="1784" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1347" />
                    <RANKING order="2" place="2" resultid="1512" />
                    <RANKING order="3" place="3" resultid="1239" />
                    <RANKING order="4" place="4" resultid="1403" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1080" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1273" />
                    <RANKING order="2" place="2" resultid="1932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1463" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1708" />
                    <RANKING order="2" place="2" resultid="1233" />
                    <RANKING order="3" place="3" resultid="1801" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1716" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2329" daytime="09:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2330" daytime="09:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2331" daytime="09:56" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1084" daytime="10:02" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1085" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1589" />
                    <RANKING order="2" place="2" resultid="1667" />
                    <RANKING order="3" place="3" resultid="1901" />
                    <RANKING order="4" place="4" resultid="1967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1970" />
                    <RANKING order="2" place="2" resultid="1815" />
                    <RANKING order="3" place="3" resultid="1388" />
                    <RANKING order="4" place="4" resultid="2027" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1228" />
                    <RANKING order="2" place="2" resultid="1338" />
                    <RANKING order="3" place="-1" resultid="1515" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1671" />
                    <RANKING order="2" place="2" resultid="1913" />
                    <RANKING order="3" place="3" resultid="1818" />
                    <RANKING order="4" place="-1" resultid="1664" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1486" />
                    <RANKING order="2" place="2" resultid="1918" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1091" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2332" daytime="10:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2333" daytime="10:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2334" daytime="10:10" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1092" daytime="10:14" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1093" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1629" />
                    <RANKING order="2" place="2" resultid="1597" />
                    <RANKING order="3" place="3" resultid="1617" />
                    <RANKING order="4" place="4" resultid="1613" />
                    <RANKING order="5" place="5" resultid="1604" />
                    <RANKING order="6" place="6" resultid="2009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1975" />
                    <RANKING order="2" place="2" resultid="1843" />
                    <RANKING order="3" place="3" resultid="1563" />
                    <RANKING order="4" place="4" resultid="1268" />
                    <RANKING order="5" place="5" resultid="1756" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1452" />
                    <RANKING order="2" place="2" resultid="1751" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1096" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1483" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1661" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1824" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2335" daytime="10:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2336" daytime="10:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2337" daytime="10:44" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1100" daytime="10:56" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1101" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1645" />
                    <RANKING order="2" place="2" resultid="1900" />
                    <RANKING order="3" place="3" resultid="1869" />
                    <RANKING order="4" place="4" resultid="1594" />
                    <RANKING order="5" place="5" resultid="1987" />
                    <RANKING order="6" place="6" resultid="1980" />
                    <RANKING order="7" place="7" resultid="1722" />
                    <RANKING order="8" place="8" resultid="1435" />
                    <RANKING order="9" place="-1" resultid="1416" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1999" />
                    <RANKING order="2" place="2" resultid="1814" />
                    <RANKING order="3" place="3" resultid="1906" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1524" />
                    <RANKING order="2" place="2" resultid="1505" />
                    <RANKING order="3" place="3" resultid="1502" />
                    <RANKING order="4" place="4" resultid="1719" />
                    <RANKING order="5" place="5" resultid="1855" />
                    <RANKING order="6" place="6" resultid="1421" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1104" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1314" />
                    <RANKING order="2" place="2" resultid="1838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1864" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1107" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1330" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2338" daytime="10:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2339" daytime="11:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2340" daytime="11:22" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1108" daytime="11:34" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1109" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1628" />
                    <RANKING order="2" place="2" resultid="1256" />
                    <RANKING order="3" place="3" resultid="1381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1110" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1543" />
                    <RANKING order="2" place="2" resultid="1547" />
                    <RANKING order="3" place="3" resultid="2395" />
                    <RANKING order="4" place="4" resultid="2021" />
                    <RANKING order="5" place="5" resultid="1842" />
                    <RANKING order="6" place="6" resultid="1875" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1236" />
                    <RANKING order="2" place="2" resultid="1896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1112" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1363" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1114" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1265" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2341" daytime="11:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2342" daytime="11:40" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1116" daytime="11:44" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1117" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1293" />
                    <RANKING order="2" place="2" resultid="1624" />
                    <RANKING order="3" place="3" resultid="1868" />
                    <RANKING order="4" place="-1" resultid="1593" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1688" />
                    <RANKING order="2" place="2" resultid="1538" />
                    <RANKING order="3" place="3" resultid="1558" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1935" />
                    <RANKING order="2" place="2" resultid="1810" />
                    <RANKING order="3" place="3" resultid="1365" />
                    <RANKING order="4" place="4" resultid="1725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1527" />
                    <RANKING order="2" place="2" resultid="1494" />
                    <RANKING order="3" place="3" resultid="1491" />
                    <RANKING order="4" place="-1" resultid="1309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1712" />
                    <RANKING order="2" place="2" resultid="1773" />
                    <RANKING order="3" place="3" resultid="1747" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1123" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1637" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2343" daytime="11:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2344" daytime="11:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2345" daytime="11:54" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1124" daytime="11:58" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1125" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1729" />
                    <RANKING order="2" place="2" resultid="1956" />
                    <RANKING order="3" place="3" resultid="1290" />
                    <RANKING order="4" place="4" resultid="1695" />
                    <RANKING order="5" place="5" resultid="1753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1974" />
                    <RANKING order="2" place="2" resultid="1551" />
                    <RANKING order="3" place="3" resultid="1880" />
                    <RANKING order="4" place="4" resultid="1994" />
                    <RANKING order="5" place="5" resultid="1650" />
                    <RANKING order="6" place="6" resultid="2020" />
                    <RANKING order="7" place="-1" resultid="1874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1769" />
                    <RANKING order="2" place="2" resultid="1475" />
                    <RANKING order="3" place="3" resultid="1451" />
                    <RANKING order="4" place="4" resultid="1750" />
                    <RANKING order="5" place="-1" resultid="1402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1285" />
                    <RANKING order="2" place="-1" resultid="1884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1130" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1925" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2346" daytime="11:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2347" daytime="12:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2348" daytime="12:02" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1132" daytime="12:06" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1133" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2002" />
                    <RANKING order="2" place="2" resultid="1608" />
                    <RANKING order="3" place="3" resultid="1585" />
                    <RANKING order="4" place="4" resultid="1581" />
                    <RANKING order="5" place="5" resultid="1427" />
                    <RANKING order="6" place="6" resultid="1674" />
                    <RANKING order="7" place="7" resultid="1434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1134" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1964" />
                    <RANKING order="2" place="2" resultid="1574" />
                    <RANKING order="3" place="3" resultid="1534" />
                    <RANKING order="4" place="4" resultid="1570" />
                    <RANKING order="5" place="5" resultid="1998" />
                    <RANKING order="6" place="6" resultid="1905" />
                    <RANKING order="7" place="7" resultid="1554" />
                    <RANKING order="8" place="8" resultid="1566" />
                    <RANKING order="9" place="9" resultid="1760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1705" />
                    <RANKING order="2" place="2" resultid="1227" />
                    <RANKING order="3" place="3" resultid="1222" />
                    <RANKING order="4" place="4" resultid="1242" />
                    <RANKING order="5" place="5" resultid="1341" />
                    <RANKING order="6" place="6" resultid="1854" />
                    <RANKING order="7" place="7" resultid="2012" />
                    <RANKING order="8" place="-1" resultid="1521" />
                    <RANKING order="9" place="-1" resultid="1732" />
                    <RANKING order="10" place="-1" resultid="1318" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1497" />
                    <RANKING order="2" place="2" resultid="1692" />
                    <RANKING order="3" place="3" resultid="1640" />
                    <RANKING order="4" place="4" resultid="1376" />
                    <RANKING order="5" place="5" resultid="1928" />
                    <RANKING order="6" place="6" resultid="1313" />
                    <RANKING order="7" place="7" resultid="1912" />
                    <RANKING order="8" place="8" resultid="1396" />
                    <RANKING order="9" place="-1" resultid="1490" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1137" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1467" />
                    <RANKING order="2" place="2" resultid="1797" />
                    <RANKING order="3" place="3" resultid="1778" />
                    <RANKING order="4" place="4" resultid="1424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1457" />
                    <RANKING order="2" place="2" resultid="1578" />
                    <RANKING order="3" place="3" resultid="1950" />
                    <RANKING order="4" place="4" resultid="1978" />
                    <RANKING order="5" place="5" resultid="1846" />
                    <RANKING order="6" place="6" resultid="1326" />
                    <RANKING order="7" place="7" resultid="1407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1139" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1531" />
                    <RANKING order="2" place="2" resultid="1335" />
                    <RANKING order="3" place="3" resultid="1323" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2349" daytime="12:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2350" daytime="12:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2351" daytime="12:12" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2352" daytime="12:14" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2353" daytime="12:16" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2354" daytime="12:18" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2355" daytime="12:20" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-10-12" daytime="15:40" endtime="17:51" number="2" officialmeeting="15:00" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1140" daytime="15:40" gender="F" number="11" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1141" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1754" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1143" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1144" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1145" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1464" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1835" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2356" daytime="15:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1148" daytime="15:48" gender="M" number="12" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1149" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1961" />
                    <RANKING order="2" place="2" resultid="1635" />
                    <RANKING order="3" place="3" resultid="1609" />
                    <RANKING order="4" place="4" resultid="1668" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1560" />
                    <RANKING order="2" place="2" resultid="1971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1151" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1229" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1152" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1915" />
                    <RANKING order="2" place="2" resultid="1839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1889" />
                    <RANKING order="2" place="2" resultid="1865" />
                    <RANKING order="3" place="-1" resultid="1425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1848" />
                    <RANKING order="2" place="-1" resultid="1409" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1851" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2357" daytime="15:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2358" daytime="15:54" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1156" daytime="16:02" gender="F" number="13" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1157" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1630" />
                    <RANKING order="2" place="2" resultid="1618" />
                    <RANKING order="3" place="3" resultid="1765" />
                    <RANKING order="4" place="4" resultid="1699" />
                    <RANKING order="5" place="5" resultid="1614" />
                    <RANKING order="6" place="6" resultid="1696" />
                    <RANKING order="7" place="7" resultid="1655" />
                    <RANKING order="8" place="8" resultid="1605" />
                    <RANKING order="9" place="9" resultid="1730" />
                    <RANKING order="10" place="10" resultid="1794" />
                    <RANKING order="11" place="11" resultid="1306" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1552" />
                    <RANKING order="2" place="2" resultid="1682" />
                    <RANKING order="3" place="3" resultid="1564" />
                    <RANKING order="4" place="4" resultid="2017" />
                    <RANKING order="5" place="5" resultid="1844" />
                    <RANKING order="6" place="6" resultid="1442" />
                    <RANKING order="7" place="7" resultid="1651" />
                    <RANKING order="8" place="8" resultid="1269" />
                    <RANKING order="9" place="9" resultid="1881" />
                    <RANKING order="10" place="10" resultid="1876" />
                    <RANKING order="11" place="-1" resultid="1281" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1453" />
                    <RANKING order="2" place="2" resultid="1770" />
                    <RANKING order="3" place="3" resultid="1941" />
                    <RANKING order="4" place="4" resultid="1404" />
                    <RANKING order="5" place="5" resultid="1954" />
                    <RANKING order="6" place="6" resultid="1351" />
                    <RANKING order="7" place="7" resultid="1897" />
                    <RANKING order="8" place="-1" resultid="1439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1160" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1861" />
                    <RANKING order="2" place="2" resultid="1892" />
                    <RANKING order="3" place="3" resultid="1274" />
                    <RANKING order="4" place="4" resultid="1807" />
                    <RANKING order="5" place="5" resultid="1286" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1161" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1484" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1162" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1662" />
                    <RANKING order="2" place="2" resultid="1926" />
                    <RANKING order="3" place="3" resultid="1709" />
                    <RANKING order="4" place="4" resultid="1836" />
                    <RANKING order="5" place="5" resultid="1740" />
                    <RANKING order="6" place="6" resultid="1802" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1163" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1825" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2359" daytime="16:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2360" daytime="16:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2361" daytime="16:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2362" daytime="16:14" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2363" daytime="16:18" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2364" daytime="16:22" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1164" daytime="16:26" gender="M" number="14" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1165" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1647" />
                    <RANKING order="2" place="2" resultid="1583" />
                    <RANKING order="3" place="3" resultid="1621" />
                    <RANKING order="4" place="4" resultid="1587" />
                    <RANKING order="5" place="5" resultid="1418" />
                    <RANKING order="6" place="6" resultid="1902" />
                    <RANKING order="7" place="7" resultid="1871" />
                    <RANKING order="8" place="8" resultid="1295" />
                    <RANKING order="9" place="9" resultid="1595" />
                    <RANKING order="10" place="10" resultid="1625" />
                    <RANKING order="11" place="11" resultid="1676" />
                    <RANKING order="12" place="12" resultid="1634" />
                    <RANKING order="13" place="13" resultid="1359" />
                    <RANKING order="14" place="14" resultid="1302" />
                    <RANKING order="15" place="15" resultid="1436" />
                    <RANKING order="16" place="-1" resultid="1601" />
                    <RANKING order="17" place="-1" resultid="1981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1559" />
                    <RANKING order="2" place="2" resultid="1576" />
                    <RANKING order="3" place="3" resultid="2025" />
                    <RANKING order="4" place="4" resultid="1536" />
                    <RANKING order="5" place="5" resultid="2000" />
                    <RANKING order="6" place="6" resultid="1539" />
                    <RANKING order="7" place="7" resultid="1572" />
                    <RANKING order="8" place="8" resultid="1354" />
                    <RANKING order="9" place="9" resultid="1392" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1224" />
                    <RANKING order="2" place="2" resultid="1479" />
                    <RANKING order="3" place="3" resultid="1461" />
                    <RANKING order="4" place="4" resultid="1832" />
                    <RANKING order="5" place="5" resultid="1506" />
                    <RANKING order="6" place="6" resultid="1243" />
                    <RANKING order="7" place="7" resultid="1857" />
                    <RANKING order="8" place="8" resultid="2014" />
                    <RANKING order="9" place="9" resultid="1734" />
                    <RANKING order="10" place="10" resultid="1385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1642" />
                    <RANKING order="2" place="2" resultid="1679" />
                    <RANKING order="3" place="3" resultid="1500" />
                    <RANKING order="4" place="4" resultid="1930" />
                    <RANKING order="5" place="5" resultid="1378" />
                    <RANKING order="6" place="6" resultid="1744" />
                    <RANKING order="7" place="7" resultid="1398" />
                    <RANKING order="8" place="8" resultid="1820" />
                    <RANKING order="9" place="-1" resultid="1372" />
                    <RANKING order="10" place="-1" resultid="1432" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1487" />
                    <RANKING order="2" place="2" resultid="1799" />
                    <RANKING order="3" place="3" resultid="1888" />
                    <RANKING order="4" place="4" resultid="1775" />
                    <RANKING order="5" place="5" resultid="1919" />
                    <RANKING order="6" place="6" resultid="1780" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1328" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1686" />
                    <RANKING order="2" place="-1" resultid="1331" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2365" daytime="16:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2366" daytime="16:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2367" daytime="16:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2368" daytime="16:38" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2369" daytime="16:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2370" daytime="16:44" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2371" daytime="16:48" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1172" daytime="16:52" gender="F" number="15" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1173" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1976" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1176" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1177" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1178" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1179" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2372" daytime="16:52" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1180" daytime="16:56" gender="M" number="16" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1181" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1610" />
                    <RANKING order="2" place="2" resultid="1988" />
                    <RANKING order="3" place="3" resultid="1429" />
                    <RANKING order="4" place="-1" resultid="1982" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1908" />
                    <RANKING order="2" place="-1" resultid="1965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1183" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1812" />
                    <RANKING order="2" place="2" resultid="1231" />
                    <RANKING order="3" place="3" resultid="1342" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1184" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1185" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1469" />
                    <RANKING order="2" place="2" resultid="1866" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2373" daytime="16:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2374" daytime="17:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1188" daytime="17:06" gender="F" number="17" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1189" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1257" />
                    <RANKING order="2" place="2" resultid="1766" />
                    <RANKING order="3" place="3" resultid="1795" />
                    <RANKING order="4" place="4" resultid="1382" />
                    <RANKING order="5" place="5" resultid="1414" />
                    <RANKING order="6" place="6" resultid="1606" />
                    <RANKING order="7" place="7" resultid="2010" />
                    <RANKING order="8" place="8" resultid="1307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1548" />
                    <RANKING order="2" place="2" resultid="1282" />
                    <RANKING order="3" place="3" resultid="2018" />
                    <RANKING order="4" place="4" resultid="2022" />
                    <RANKING order="5" place="5" resultid="1786" />
                    <RANKING order="6" place="6" resultid="1247" />
                    <RANKING order="7" place="7" resultid="1877" />
                    <RANKING order="8" place="8" resultid="1882" />
                    <RANKING order="9" place="-1" resultid="1299" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1237" />
                    <RANKING order="2" place="2" resultid="1455" />
                    <RANKING order="3" place="3" resultid="1519" />
                    <RANKING order="4" place="4" resultid="1898" />
                    <RANKING order="5" place="5" resultid="1771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1862" />
                    <RANKING order="2" place="2" resultid="1808" />
                    <RANKING order="3" place="3" resultid="1893" />
                    <RANKING order="4" place="4" resultid="2030" />
                    <RANKING order="5" place="5" resultid="1287" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1194" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1266" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2375" daytime="17:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2376" daytime="17:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2377" daytime="17:12" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2378" daytime="17:16" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1196" daytime="17:18" gender="M" number="18" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1197" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1648" />
                    <RANKING order="2" place="2" resultid="1962" />
                    <RANKING order="3" place="3" resultid="1296" />
                    <RANKING order="4" place="4" resultid="1626" />
                    <RANKING order="5" place="5" resultid="1872" />
                    <RANKING order="6" place="6" resultid="1303" />
                    <RANKING order="7" place="7" resultid="1262" />
                    <RANKING order="8" place="8" resultid="1790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1690" />
                    <RANKING order="2" place="2" resultid="1556" />
                    <RANKING order="3" place="3" resultid="1540" />
                    <RANKING order="4" place="4" resultid="1356" />
                    <RANKING order="5" place="5" resultid="1393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1199" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1936" />
                    <RANKING order="2" place="2" resultid="1225" />
                    <RANKING order="3" place="3" resultid="1525" />
                    <RANKING order="4" place="4" resultid="1345" />
                    <RANKING order="5" place="5" resultid="1706" />
                    <RANKING order="6" place="6" resultid="1480" />
                    <RANKING order="7" place="7" resultid="1939" />
                    <RANKING order="8" place="8" resultid="1720" />
                    <RANKING order="9" place="9" resultid="1366" />
                    <RANKING order="10" place="10" resultid="1503" />
                    <RANKING order="11" place="11" resultid="1735" />
                    <RANKING order="12" place="-1" resultid="1319" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1200" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1529" />
                    <RANKING order="2" place="2" resultid="1703" />
                    <RANKING order="3" place="3" resultid="1492" />
                    <RANKING order="4" place="4" resultid="1495" />
                    <RANKING order="5" place="5" resultid="1745" />
                    <RANKING order="6" place="6" resultid="1399" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1201" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1713" />
                    <RANKING order="2" place="2" resultid="1776" />
                    <RANKING order="3" place="3" resultid="1781" />
                    <RANKING order="4" place="4" resultid="1830" />
                    <RANKING order="5" place="-1" resultid="1468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1203" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1638" />
                    <RANKING order="2" place="2" resultid="1324" />
                    <RANKING order="3" place="3" resultid="1852" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2379" daytime="17:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2380" daytime="17:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2381" daytime="17:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2382" daytime="17:28" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2383" daytime="17:30" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1204" daytime="17:34" gender="F" number="19" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1205" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1447" />
                    <RANKING order="2" place="2" resultid="1700" />
                    <RANKING order="3" place="3" resultid="1985" />
                    <RANKING order="4" place="4" resultid="1631" />
                    <RANKING order="5" place="5" resultid="1656" />
                    <RANKING order="6" place="6" resultid="1958" />
                    <RANKING order="7" place="7" resultid="1278" />
                    <RANKING order="8" place="8" resultid="1413" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1206" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1683" />
                    <RANKING order="2" place="2" resultid="1992" />
                    <RANKING order="3" place="3" resultid="1449" />
                    <RANKING order="4" place="4" resultid="1473" />
                    <RANKING order="5" place="5" resultid="1996" />
                    <RANKING order="6" place="6" resultid="1785" />
                    <RANKING order="7" place="7" resultid="1544" />
                    <RANKING order="8" place="8" resultid="1652" />
                    <RANKING order="9" place="9" resultid="1246" />
                    <RANKING order="10" place="10" resultid="1253" />
                    <RANKING order="11" place="-1" resultid="1270" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1509" />
                    <RANKING order="2" place="2" resultid="1348" />
                    <RANKING order="3" place="3" resultid="1513" />
                    <RANKING order="4" place="4" resultid="1476" />
                    <RANKING order="5" place="5" resultid="1240" />
                    <RANKING order="6" place="6" resultid="1405" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1659" />
                    <RANKING order="2" place="2" resultid="1275" />
                    <RANKING order="3" place="3" resultid="1885" />
                    <RANKING order="4" place="4" resultid="1933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1465" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1210" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1710" />
                    <RANKING order="2" place="2" resultid="1234" />
                    <RANKING order="3" place="3" resultid="1803" />
                    <RANKING order="4" place="4" resultid="1741" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1717" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2384" daytime="17:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2385" daytime="17:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2386" daytime="17:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2387" daytime="17:42" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2388" daytime="17:44" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1212" daytime="17:48" gender="M" number="20" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1213" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1591" />
                    <RANKING order="2" place="2" resultid="1622" />
                    <RANKING order="3" place="3" resultid="1250" />
                    <RANKING order="4" place="4" resultid="1903" />
                    <RANKING order="5" place="5" resultid="1669" />
                    <RANKING order="6" place="6" resultid="1968" />
                    <RANKING order="7" place="7" resultid="1419" />
                    <RANKING order="8" place="8" resultid="1723" />
                    <RANKING order="9" place="9" resultid="1360" />
                    <RANKING order="10" place="10" resultid="1789" />
                    <RANKING order="11" place="11" resultid="2006" />
                    <RANKING order="12" place="-1" resultid="1602" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1816" />
                    <RANKING order="2" place="2" resultid="1972" />
                    <RANKING order="3" place="3" resultid="2028" />
                    <RANKING order="4" place="4" resultid="1389" />
                    <RANKING order="5" place="5" resultid="1369" />
                    <RANKING order="6" place="6" resultid="1355" />
                    <RANKING order="7" place="-1" resultid="1568" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1833" />
                    <RANKING order="2" place="2" resultid="1230" />
                    <RANKING order="3" place="3" resultid="1516" />
                    <RANKING order="4" place="4" resultid="1339" />
                    <RANKING order="5" place="5" resultid="1948" />
                    <RANKING order="6" place="6" resultid="1726" />
                    <RANKING order="7" place="-1" resultid="1386" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1216" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1665" />
                    <RANKING order="2" place="2" resultid="1672" />
                    <RANKING order="3" place="3" resultid="1643" />
                    <RANKING order="4" place="4" resultid="1916" />
                    <RANKING order="5" place="5" resultid="1840" />
                    <RANKING order="6" place="-1" resultid="1821" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1488" />
                    <RANKING order="2" place="2" resultid="1920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1321" />
                    <RANKING order="2" place="-1" resultid="1410" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1532" />
                    <RANKING order="2" place="2" resultid="1333" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2389" daytime="17:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2390" daytime="17:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2391" daytime="17:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2392" daytime="17:56" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2393" daytime="17:58" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="13038" nation="BRA" region="PR" clubid="1263" swrid="93759" name="Associação De Pais E Atletas De Natação Ws/Crb" shortname="Apan/Ws">
          <ATHLETES>
            <ATHLETE firstname="Marjori" lastname="Leticia Oliveira" birthdate="2011-05-23" gender="F" nation="BRA" license="406869" swrid="5717279" athleteid="1304" externalid="406869">
              <RESULTS>
                <RESULT eventid="1060" points="291" swimtime="00:01:18.01" resultid="1305" heatid="2313" lane="3" entrytime="00:01:19.21" entrycourse="LCM" />
                <RESULT eventid="1156" points="266" swimtime="00:02:55.39" resultid="1306" heatid="2360" lane="3" entrytime="00:02:57.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="203" swimtime="00:01:37.44" resultid="1307" heatid="2376" lane="6" entrytime="00:01:30.86" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Fernandes Ferreira" birthdate="2008-07-28" gender="M" nation="BRA" license="414578" swrid="5755373" athleteid="1308" externalid="414578">
              <RESULTS>
                <RESULT eventid="1116" status="DNS" swimtime="00:00:00.00" resultid="1309" heatid="2343" lane="4" />
                <RESULT eventid="1068" points="335" swimtime="00:01:07.44" resultid="1310" heatid="2323" lane="6" entrytime="00:01:03.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Zeclhynski Silva" birthdate="2006-09-14" gender="F" nation="BRA" license="330727" swrid="5600283" athleteid="1264" externalid="330727">
              <RESULTS>
                <RESULT eventid="1108" points="506" swimtime="00:02:34.50" resultid="1265" heatid="2342" lane="4" entrytime="00:02:34.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="583" swimtime="00:01:08.60" resultid="1266" heatid="2378" lane="4" entrytime="00:01:06.10" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Reis" birthdate="2008-04-07" gender="F" nation="BRA" license="378820" swrid="5600243" athleteid="1283" externalid="378820">
              <RESULTS>
                <RESULT eventid="1060" points="272" swimtime="00:01:19.75" resultid="1284" heatid="2313" lane="6" entrytime="00:01:20.14" entrycourse="LCM" />
                <RESULT eventid="1124" points="187" swimtime="00:01:36.99" resultid="1285" heatid="2348" lane="8" entrytime="00:01:36.96" entrycourse="LCM" />
                <RESULT eventid="1156" points="258" swimtime="00:02:57.15" resultid="1286" heatid="2360" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="233" swimtime="00:01:33.11" resultid="1287" heatid="2376" lane="3" entrytime="00:01:30.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Rosa Silva" birthdate="2011-03-25" gender="F" nation="BRA" license="392120" swrid="5602579" athleteid="1276" externalid="392120">
              <RESULTS>
                <RESULT eventid="1060" points="264" swimtime="00:01:20.55" resultid="1277" heatid="2313" lane="1" entrytime="00:01:21.95" entrycourse="LCM" />
                <RESULT eventid="1204" points="210" swimtime="00:01:47.77" resultid="1278" heatid="2384" lane="4" entrytime="00:01:44.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabelly" lastname="Mendonca Bello" birthdate="2008-04-15" gender="F" nation="BRA" license="376996" swrid="5600217" athleteid="1271" externalid="376996">
              <RESULTS>
                <RESULT eventid="1060" points="488" swimtime="00:01:05.65" resultid="1272" heatid="2316" lane="4" entrytime="00:01:07.89" entrycourse="LCM" />
                <RESULT eventid="1076" points="378" swimtime="00:03:10.23" resultid="1273" heatid="2330" lane="3" entrytime="00:03:09.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="457" swimtime="00:02:26.48" resultid="1274" heatid="2360" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="392" swimtime="00:01:27.58" resultid="1275" heatid="2387" lane="7" entrytime="00:01:24.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Sieck" birthdate="2011-01-20" gender="F" nation="BRA" license="382234" swrid="5602584" athleteid="1288" externalid="382234">
              <RESULTS>
                <RESULT eventid="1060" points="233" swimtime="00:01:23.97" resultid="1289" heatid="2313" lane="8" entrytime="00:01:25.84" entrycourse="LCM" />
                <RESULT eventid="1124" points="186" swimtime="00:01:37.09" resultid="1290" heatid="2347" lane="4" entrytime="00:01:37.33" entrycourse="LCM" />
                <RESULT eventid="1172" points="141" swimtime="00:03:53.84" resultid="1291" heatid="2372" lane="5" entrytime="00:03:43.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Zanchetta Silva" birthdate="2010-08-05" gender="F" nation="BRA" license="406865" swrid="5717308" athleteid="1297" externalid="406865">
              <RESULTS>
                <RESULT eventid="1060" status="DNS" swimtime="00:00:00.00" resultid="1298" heatid="2313" lane="7" entrytime="00:01:21.27" entrycourse="LCM" />
                <RESULT eventid="1188" status="DNS" swimtime="00:00:00.00" resultid="1299" heatid="2376" lane="8" entrytime="00:01:41.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="De Reginalda" birthdate="2011-07-22" gender="M" nation="BRA" license="400323" swrid="5717257" athleteid="1292" externalid="400323">
              <RESULTS>
                <RESULT eventid="1116" points="363" swimtime="00:02:36.84" resultid="1293" heatid="2344" lane="5" entrytime="00:02:39.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="416" swimtime="00:01:02.75" resultid="1294" heatid="2324" lane="1" entrytime="00:01:02.15" entrycourse="LCM" />
                <RESULT eventid="1164" points="332" swimtime="00:02:27.21" resultid="1295" heatid="2365" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="364" swimtime="00:01:12.24" resultid="1296" heatid="2381" lane="6" entrytime="00:01:12.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Daniele Silva" birthdate="2010-07-06" gender="F" nation="BRA" license="359593" swrid="5588628" athleteid="1279" externalid="359593">
              <RESULTS>
                <RESULT eventid="1060" points="458" swimtime="00:01:07.05" resultid="1280" heatid="2317" lane="4" entrytime="00:01:06.02" entrycourse="LCM" />
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="1281" heatid="2362" lane="1" entrytime="00:02:34.42" entrycourse="LCM" />
                <RESULT eventid="1188" points="397" swimtime="00:01:17.94" resultid="1282" heatid="2378" lane="1" entrytime="00:01:17.58" entrycourse="LCM" />
                <RESULT eventid="1108" points="372" swimtime="00:02:51.07" resultid="2395" heatid="2341" lane="7" late="yes" entrytime="00:02:54.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonia" lastname="Adam  Fracaro" birthdate="2010-04-27" gender="F" nation="BRA" license="382212" swrid="5588512" athleteid="1267" externalid="382212">
              <RESULTS>
                <RESULT eventid="1092" points="269" swimtime="00:12:30.94" resultid="1268" heatid="2336" lane="6" entrytime="00:12:35.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.59" />
                    <SPLIT distance="200" swimtime="00:02:59.17" />
                    <SPLIT distance="300" swimtime="00:04:34.81" />
                    <SPLIT distance="400" swimtime="00:06:10.85" />
                    <SPLIT distance="500" swimtime="00:07:46.96" />
                    <SPLIT distance="600" swimtime="00:09:23.53" />
                    <SPLIT distance="700" swimtime="00:11:00.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="294" swimtime="00:02:49.53" resultid="1269" heatid="2361" lane="7" entrytime="00:02:43.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" status="DNS" swimtime="00:00:00.00" resultid="1270" heatid="2384" lane="5" entrytime="00:01:58.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Cravcenco Marcondes" birthdate="2011-05-06" gender="M" nation="BRA" license="406867" swrid="5723023" athleteid="1300" externalid="406867">
              <RESULTS>
                <RESULT eventid="1068" points="289" swimtime="00:01:10.87" resultid="1301" heatid="2320" lane="6" entrytime="00:01:10.73" entrycourse="LCM" />
                <RESULT eventid="1164" points="245" swimtime="00:02:42.90" resultid="1302" heatid="2365" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="190" swimtime="00:01:29.70" resultid="1303" heatid="2380" lane="1" entrytime="00:01:35.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2539" nation="BRA" region="PR" clubid="1394" swrid="93771" name="Círculo Militar Do Paraná" shortname="Círculo Militar">
          <ATHLETES>
            <ATHLETE firstname="Gustavo" lastname="De Queiroz" birthdate="2007-08-20" gender="M" nation="BRA" license="406949" swrid="5717256" athleteid="1423" externalid="406949">
              <RESULTS>
                <RESULT eventid="1132" points="214" swimtime="00:01:22.59" resultid="1424" heatid="2351" lane="1" entrytime="00:01:29.84" entrycourse="LCM" />
                <RESULT comment="SW 8.5 - Totalmente submerso durante o nado.  (Tempo: 15:58), Medley Indvidual, Borboleta." eventid="1148" status="DSQ" swimtime="00:06:51.55" resultid="1425" heatid="2357" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.05" />
                    <SPLIT distance="200" swimtime="00:03:21.70" />
                    <SPLIT distance="300" swimtime="00:05:17.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Vieira De Macedo Brasil" birthdate="2009-12-19" gender="F" nation="BRA" license="344143" swrid="5622311" athleteid="1400" externalid="344143">
              <RESULTS>
                <RESULT eventid="1060" points="425" swimtime="00:01:08.77" resultid="1401" heatid="2315" lane="2" entrytime="00:01:10.94" entrycourse="LCM" />
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="1402" heatid="2347" lane="2" />
                <RESULT eventid="1076" points="299" swimtime="00:03:25.56" resultid="1403" heatid="2329" lane="4" entrytime="00:03:34.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="433" swimtime="00:02:29.11" resultid="1404" heatid="2362" lane="8" entrytime="00:02:34.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="320" swimtime="00:01:33.73" resultid="1405" heatid="2386" lane="1" entrytime="00:01:32.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Maria Romanelli" birthdate="2011-04-18" gender="F" nation="BRA" license="378335" swrid="5588803" athleteid="1411" externalid="378335">
              <RESULTS>
                <RESULT eventid="1060" points="411" swimtime="00:01:09.52" resultid="1412" heatid="2315" lane="4" entrytime="00:01:10.02" entrycourse="LCM" />
                <RESULT eventid="1204" points="195" swimtime="00:01:50.50" resultid="1413" heatid="2385" lane="1" entrytime="00:01:44.29" entrycourse="LCM" />
                <RESULT eventid="1188" points="278" swimtime="00:01:27.84" resultid="1414" heatid="2376" lane="5" entrytime="00:01:30.32" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Flavia" lastname="Scheffler Souza" birthdate="2010-09-14" gender="F" nation="BRA" license="417278" swrid="5757095" athleteid="1440" externalid="417278">
              <RESULTS>
                <RESULT eventid="1060" points="371" swimtime="00:01:11.92" resultid="1441" heatid="2314" lane="5" entrytime="00:01:12.71" entrycourse="LCM" />
                <RESULT eventid="1156" points="363" swimtime="00:02:38.16" resultid="1442" heatid="2360" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernando" lastname="Jun Melo Ogima" birthdate="2006-07-05" gender="M" nation="BRA" license="378332" swrid="5622284" athleteid="1406" externalid="378332">
              <RESULTS>
                <RESULT eventid="1132" points="276" swimtime="00:01:15.93" resultid="1407" heatid="2351" lane="7" entrytime="00:01:21.13" entrycourse="LCM" />
                <RESULT eventid="1068" points="410" swimtime="00:01:03.05" resultid="1408" heatid="2324" lane="7" entrytime="00:01:02.12" entrycourse="LCM" />
                <RESULT comment="SW 8.5 - Totalmente submerso durante o nado.  (Tempo: 15:58), Medley Indvidual, Borboleta." eventid="1148" status="DSQ" swimtime="00:06:24.78" resultid="1409" heatid="2357" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.53" />
                    <SPLIT distance="200" swimtime="00:03:06.26" />
                    <SPLIT distance="300" swimtime="00:04:55.32" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.5 - Executou uma pernada de borboleta durante o nado.  (Tempo: 17:46)" eventid="1212" status="DSQ" swimtime="00:01:27.67" resultid="1410" heatid="2391" lane="1" entrytime="00:01:27.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thomas" lastname="Gomes" birthdate="2009-06-15" gender="M" nation="BRA" license="406948" swrid="5717268" athleteid="1420" externalid="406948">
              <RESULTS>
                <RESULT eventid="1100" points="211" swimtime="00:12:39.08" resultid="1421" heatid="2338" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.72" />
                    <SPLIT distance="200" swimtime="00:02:59.26" />
                    <SPLIT distance="300" swimtime="00:04:35.61" />
                    <SPLIT distance="400" swimtime="00:06:13.17" />
                    <SPLIT distance="500" swimtime="00:07:52.24" />
                    <SPLIT distance="600" swimtime="00:09:29.62" />
                    <SPLIT distance="700" swimtime="00:11:07.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="243" swimtime="00:01:15.07" resultid="1422" heatid="2320" lane="2" entrytime="00:01:14.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Karuta" birthdate="2011-10-31" gender="M" nation="BRA" license="414648" swrid="5755375" athleteid="1433" externalid="414648">
              <RESULTS>
                <RESULT eventid="1132" points="104" swimtime="00:01:45.08" resultid="1434" heatid="2350" lane="6" />
                <RESULT eventid="1100" points="249" swimtime="00:11:57.84" resultid="1435" heatid="2339" lane="8" entrytime="00:11:46.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.18" />
                    <SPLIT distance="200" swimtime="00:02:51.61" />
                    <SPLIT distance="300" swimtime="00:04:23.75" />
                    <SPLIT distance="400" swimtime="00:05:57.44" />
                    <SPLIT distance="500" swimtime="00:07:28.65" />
                    <SPLIT distance="600" swimtime="00:08:59.64" />
                    <SPLIT distance="700" swimtime="00:10:29.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="242" swimtime="00:02:43.62" resultid="1436" heatid="2366" lane="1" entrytime="00:02:44.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicole" lastname="Herdy Faria" birthdate="2009-11-10" gender="F" nation="BRA" license="417277" swrid="5757091" athleteid="1437" externalid="417277">
              <RESULTS>
                <RESULT eventid="1060" points="375" swimtime="00:01:11.66" resultid="1438" heatid="2315" lane="7" entrytime="00:01:11.18" entrycourse="LCM" />
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="1439" heatid="2359" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vicente" lastname="Bileski" birthdate="2011-06-29" gender="M" nation="BRA" license="406950" swrid="5717248" athleteid="1426" externalid="406950">
              <RESULTS>
                <RESULT eventid="1132" points="245" swimtime="00:01:19.00" resultid="1427" heatid="2351" lane="8" entrytime="00:01:42.26" entrycourse="LCM" />
                <RESULT eventid="1068" points="263" swimtime="00:01:13.08" resultid="1428" heatid="2320" lane="7" entrytime="00:01:14.97" entrycourse="LCM" />
                <RESULT eventid="1180" points="189" swimtime="00:03:12.25" resultid="1429" heatid="2373" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Oliveira Martini" birthdate="2008-10-31" gender="M" nation="BRA" license="406953" swrid="5717285" athleteid="1430" externalid="406953">
              <RESULTS>
                <RESULT eventid="1068" status="DNS" swimtime="00:00:00.00" resultid="1431" heatid="2322" lane="7" entrytime="00:01:05.12" entrycourse="LCM" />
                <RESULT eventid="1164" status="DNS" swimtime="00:00:00.00" resultid="1432" heatid="2367" lane="8" entrytime="00:02:33.89" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Manocchio" birthdate="2011-07-28" gender="M" nation="BRA" license="384916" swrid="5588573" athleteid="1415" externalid="384916">
              <RESULTS>
                <RESULT eventid="1100" status="DNS" swimtime="00:00:00.00" resultid="1416" heatid="2340" lane="8" entrytime="00:10:35.76" entrycourse="LCM" />
                <RESULT eventid="1068" points="410" swimtime="00:01:03.03" resultid="1417" heatid="2323" lane="4" entrytime="00:01:03.00" entrycourse="LCM" />
                <RESULT eventid="1164" points="386" swimtime="00:02:20.08" resultid="1418" heatid="2368" lane="1" entrytime="00:02:21.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="261" swimtime="00:01:28.95" resultid="1419" heatid="2390" lane="3" entrytime="00:01:29.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Torres Oliveira" birthdate="2008-04-10" gender="M" nation="BRA" license="400274" swrid="5653303" athleteid="1395" externalid="400274">
              <RESULTS>
                <RESULT eventid="1132" points="236" swimtime="00:01:19.97" resultid="1396" heatid="2349" lane="3" />
                <RESULT eventid="1068" points="383" swimtime="00:01:04.50" resultid="1397" heatid="2323" lane="3" entrytime="00:01:03.03" entrycourse="LCM" />
                <RESULT eventid="1164" points="311" swimtime="00:02:30.44" resultid="1398" heatid="2367" lane="6" entrytime="00:02:26.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="236" swimtime="00:01:23.47" resultid="1399" heatid="2379" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="12782" nation="BRA" region="PR" clubid="1714" swrid="93773" name="Clube Duque De Caxias" shortname="Duque De Caxias">
          <ATHLETES>
            <ATHLETE firstname="Lucas" lastname="Bulgarelli Castro" birthdate="2009-04-20" gender="M" nation="BRA" license="401867" swrid="5658058" athleteid="1724" externalid="401867">
              <RESULTS>
                <RESULT eventid="1116" points="224" swimtime="00:03:04.07" resultid="1725" heatid="2343" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="244" swimtime="00:01:30.92" resultid="1726" heatid="2389" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ian" lastname="Berger" birthdate="2011-07-27" gender="M" nation="BRA" license="387966" swrid="5652879" athleteid="1721" externalid="387966">
              <RESULTS>
                <RESULT eventid="1100" points="281" swimtime="00:11:29.87" resultid="1722" heatid="2338" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.65" />
                    <SPLIT distance="200" swimtime="00:02:45.69" />
                    <SPLIT distance="300" swimtime="00:04:14.21" />
                    <SPLIT distance="400" swimtime="00:05:42.59" />
                    <SPLIT distance="500" swimtime="00:07:10.68" />
                    <SPLIT distance="600" swimtime="00:08:39.86" />
                    <SPLIT distance="700" swimtime="00:10:06.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="236" swimtime="00:01:31.99" resultid="1723" heatid="2390" lane="8" entrytime="00:01:42.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tayla" lastname="Kalluf Oliveira" birthdate="2011-12-05" gender="F" nation="BRA" license="414583" swrid="5755374" athleteid="1727" externalid="414583">
              <RESULTS>
                <RESULT eventid="1060" points="425" swimtime="00:01:08.73" resultid="1728" heatid="2316" lane="6" entrytime="00:01:08.39" entrycourse="LCM" />
                <RESULT eventid="1124" points="351" swimtime="00:01:18.62" resultid="1729" heatid="2346" lane="5" />
                <RESULT eventid="1156" points="364" swimtime="00:02:38.04" resultid="1730" heatid="2359" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Vitor Girelli" birthdate="2009-08-01" gender="M" nation="BRA" license="387965" swrid="5622312" athleteid="1718" externalid="387965">
              <RESULTS>
                <RESULT eventid="1100" points="374" swimtime="00:10:27.01" resultid="1719" heatid="2338" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.93" />
                    <SPLIT distance="200" swimtime="00:02:28.33" />
                    <SPLIT distance="300" swimtime="00:03:47.36" />
                    <SPLIT distance="400" swimtime="00:05:05.29" />
                    <SPLIT distance="500" swimtime="00:06:29.04" />
                    <SPLIT distance="600" swimtime="00:07:47.46" />
                    <SPLIT distance="700" swimtime="00:09:09.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="398" swimtime="00:01:10.13" resultid="1720" heatid="2381" lane="1" entrytime="00:01:15.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Flavia Braz" birthdate="2004-10-25" gender="F" nation="BRA" license="280573" swrid="5622281" athleteid="1715" externalid="280573">
              <RESULTS>
                <RESULT eventid="1076" points="447" swimtime="00:02:59.84" resultid="1716" heatid="2331" lane="1" entrytime="00:02:59.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="540" swimtime="00:01:18.75" resultid="1717" heatid="2387" lane="5" entrytime="00:01:22.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Kovalhuk Lima" birthdate="2009-03-16" gender="M" nation="BRA" license="417452" athleteid="1731" externalid="417452">
              <RESULTS>
                <RESULT comment="SW 8.2 - Braços não trazidos para frente simultaneamente sobre (em cima) a água., Nadou crawl." eventid="1132" status="DSQ" swimtime="00:01:24.86" resultid="1732" heatid="2350" lane="3" />
                <RESULT eventid="1068" points="366" swimtime="00:01:05.50" resultid="1733" heatid="2319" lane="6" />
                <RESULT eventid="1164" points="296" swimtime="00:02:33.03" resultid="1734" heatid="2365" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="261" swimtime="00:01:20.69" resultid="1735" heatid="2379" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11303" nation="BRA" region="PR" clubid="1316" swrid="93760" name="Associação De Talentos Da Natação" shortname="Atn/Curitiba">
          <ATHLETES>
            <ATHLETE firstname="Mauricio" lastname="Furtado Niwa" birthdate="1978-05-30" gender="M" nation="BRA" license="398757" swrid="5653291" athleteid="1334" externalid="398757">
              <RESULTS>
                <RESULT eventid="1132" points="501" swimtime="00:01:02.26" resultid="1335" heatid="2354" lane="3" entrytime="00:01:01.95" entrycourse="LCM" />
                <RESULT eventid="1068" points="499" swimtime="00:00:59.04" resultid="1336" heatid="2326" lane="7" entrytime="00:00:58.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Yuji Yamazato" birthdate="2008-10-01" gender="M" nation="BRA" license="392664" swrid="5622313" athleteid="1370" externalid="392664">
              <RESULTS>
                <RESULT eventid="1068" points="399" swimtime="00:01:03.63" resultid="1371" heatid="2323" lane="1" entrytime="00:01:03.80" entrycourse="LCM" />
                <RESULT eventid="1164" status="DNS" swimtime="00:00:00.00" resultid="1372" heatid="2366" lane="4" entrytime="00:02:34.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Garcia De Fraga" birthdate="2009-03-24" gender="M" nation="BRA" license="342147" swrid="5600172" athleteid="1317" externalid="342147">
              <RESULTS>
                <RESULT eventid="1132" status="DNS" swimtime="00:00:00.00" resultid="1318" heatid="2355" lane="8" entrytime="00:01:00.74" entrycourse="LCM" />
                <RESULT eventid="1196" status="DNS" swimtime="00:00:00.00" resultid="1319" heatid="2383" lane="3" entrytime="00:01:00.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Araujo Do Rego Barros" birthdate="2009-04-30" gender="M" nation="BRA" license="376325" swrid="5377739" athleteid="1340" externalid="376325">
              <RESULTS>
                <RESULT eventid="1132" points="363" swimtime="00:01:09.27" resultid="1341" heatid="2353" lane="2" entrytime="00:01:09.00" entrycourse="LCM" />
                <RESULT eventid="1180" points="325" swimtime="00:02:40.46" resultid="1342" heatid="2374" lane="6" entrytime="00:02:36.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Navarro Silva" birthdate="2011-01-10" gender="F" nation="BRA" license="406711" swrid="5717284" athleteid="1379" externalid="406711">
              <RESULTS>
                <RESULT eventid="1060" points="356" swimtime="00:01:12.94" resultid="1380" heatid="2314" lane="7" entrytime="00:01:16.00" entrycourse="LCM" />
                <RESULT eventid="1108" points="255" swimtime="00:03:14.14" resultid="1381" heatid="2341" lane="3" entrytime="00:03:06.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="288" swimtime="00:01:26.72" resultid="1382" heatid="2377" lane="1" entrytime="00:01:25.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcos" lastname="Demchuk" birthdate="2011-06-15" gender="M" nation="BRA" license="388540" swrid="5602530" athleteid="1357" externalid="388540">
              <RESULTS>
                <RESULT eventid="1068" points="332" swimtime="00:01:07.67" resultid="1358" heatid="2320" lane="3" entrytime="00:01:09.05" entrycourse="LCM" />
                <RESULT eventid="1164" points="260" swimtime="00:02:39.70" resultid="1359" heatid="2365" lane="5" entrytime="00:03:09.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="200" swimtime="00:01:37.20" resultid="1360" heatid="2390" lane="7" entrytime="00:01:32.57" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Muller" birthdate="2009-10-10" gender="F" nation="BRA" license="376952" swrid="5600221" athleteid="1346" externalid="376952">
              <RESULTS>
                <RESULT eventid="1076" points="443" swimtime="00:03:00.43" resultid="1347" heatid="2331" lane="7" entrytime="00:02:59.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="485" swimtime="00:01:21.60" resultid="1348" heatid="2388" lane="2" entrytime="00:01:19.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Castellano Purkot" birthdate="2010-01-25" gender="M" nation="BRA" license="392484" swrid="5622268" athleteid="1367" externalid="392484">
              <RESULTS>
                <RESULT eventid="1068" points="286" swimtime="00:01:11.05" resultid="1368" heatid="2320" lane="5" entrytime="00:01:08.39" entrycourse="LCM" />
                <RESULT eventid="1212" points="244" swimtime="00:01:31.00" resultid="1369" heatid="2390" lane="2" entrytime="00:01:31.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Kerppers Kreia" birthdate="2006-12-01" gender="M" nation="BRA" license="366815" swrid="5600195" athleteid="1325" externalid="366815">
              <RESULTS>
                <RESULT eventid="1132" points="372" swimtime="00:01:08.71" resultid="1326" heatid="2352" lane="3" entrytime="00:01:12.73" entrycourse="LCM" />
                <RESULT eventid="1068" points="516" swimtime="00:00:58.42" resultid="1327" heatid="2326" lane="3" entrytime="00:00:58.10" entrycourse="LCM" />
                <RESULT eventid="1164" points="495" swimtime="00:02:08.88" resultid="1328" heatid="2370" lane="3" entrytime="00:02:10.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Riccieri" lastname="Rodrigues Muzolon" birthdate="2010-11-08" gender="M" nation="BRA" license="385439" swrid="5588887" athleteid="1352" externalid="385439">
              <RESULTS>
                <RESULT eventid="1068" points="361" swimtime="00:01:05.81" resultid="1353" heatid="2321" lane="5" entrytime="00:01:06.19" entrycourse="LCM" />
                <RESULT eventid="1164" points="282" swimtime="00:02:35.54" resultid="1354" heatid="2366" lane="3" entrytime="00:02:34.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="237" swimtime="00:01:31.82" resultid="1355" heatid="2390" lane="4" entrytime="00:01:28.01" entrycourse="LCM" />
                <RESULT eventid="1196" points="274" swimtime="00:01:19.40" resultid="1356" heatid="2380" lane="5" entrytime="00:01:17.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Neves Vianna" birthdate="2007-12-30" gender="F" nation="BRA" license="391106" swrid="5600223" athleteid="1361" externalid="391106">
              <RESULTS>
                <RESULT eventid="1060" points="262" swimtime="00:01:20.74" resultid="1362" heatid="2313" lane="2" entrytime="00:01:20.18" entrycourse="LCM" />
                <RESULT eventid="1108" points="206" swimtime="00:03:28.25" resultid="1363" heatid="2341" lane="6" entrytime="00:03:20.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Arthur Ribeiro" birthdate="2010-02-05" gender="M" nation="BRA" license="408025" swrid="5723020" athleteid="1387" externalid="408025">
              <RESULTS>
                <RESULT eventid="1084" points="303" swimtime="00:03:06.66" resultid="1388" heatid="2333" lane="3" entrytime="00:03:11.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="308" swimtime="00:01:24.14" resultid="1389" heatid="2391" lane="6" entrytime="00:01:24.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Iglesias Prado" birthdate="2010-06-15" gender="M" nation="BRA" license="408052" swrid="5723025" athleteid="1390" externalid="408052">
              <RESULTS>
                <RESULT eventid="1068" points="334" swimtime="00:01:07.48" resultid="1391" heatid="2321" lane="7" entrytime="00:01:07.21" entrycourse="LCM" />
                <RESULT eventid="1164" points="268" swimtime="00:02:38.16" resultid="1392" heatid="2366" lane="2" entrytime="00:02:37.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="270" swimtime="00:01:19.74" resultid="1393" heatid="2380" lane="2" entrytime="00:01:24.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Ocanha" birthdate="2005-06-21" gender="M" nation="BRA" license="313769" swrid="5600231" athleteid="1320" externalid="313769">
              <RESULTS>
                <RESULT eventid="1212" points="519" swimtime="00:01:10.77" resultid="1321" heatid="2393" lane="7" entrytime="00:01:10.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Kerniski Demantova" birthdate="1982-05-25" gender="M" nation="BRA" license="398222" swrid="5653293" athleteid="1329" externalid="398222">
              <RESULTS>
                <RESULT eventid="1100" status="DNS" swimtime="00:00:00.00" resultid="1330" heatid="2340" lane="3" entrytime="00:10:20.99" entrycourse="LCM" />
                <RESULT eventid="1164" status="DNS" swimtime="00:00:00.00" resultid="1331" heatid="2368" lane="7" entrytime="00:02:21.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Bortoleto" birthdate="2008-09-05" gender="M" nation="BRA" license="406709" swrid="5717249" athleteid="1375" externalid="406709">
              <RESULTS>
                <RESULT eventid="1132" points="397" swimtime="00:01:07.26" resultid="1376" heatid="2353" lane="6" entrytime="00:01:08.93" entrycourse="LCM" />
                <RESULT eventid="1068" points="506" swimtime="00:00:58.77" resultid="1377" heatid="2325" lane="3" entrytime="00:00:59.45" entrycourse="LCM" />
                <RESULT eventid="1164" points="447" swimtime="00:02:13.37" resultid="1378" heatid="2369" lane="3" entrytime="00:02:15.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Angelo" lastname="De Queiroz Neto" birthdate="2003-10-31" gender="M" nation="BRA" license="342814" swrid="5600149" athleteid="1322" externalid="342814">
              <RESULTS>
                <RESULT eventid="1132" points="423" swimtime="00:01:05.84" resultid="1323" heatid="2353" lane="4" entrytime="00:01:05.71" entrycourse="LCM" />
                <RESULT eventid="1196" points="354" swimtime="00:01:12.90" resultid="1324" heatid="2379" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelo" lastname="Correia Bonfim" birthdate="2009-06-21" gender="M" nation="BRA" license="391663" swrid="5622271" athleteid="1364" externalid="391663">
              <RESULTS>
                <RESULT eventid="1116" points="319" swimtime="00:02:43.72" resultid="1365" heatid="2344" lane="6" entrytime="00:02:44.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="332" swimtime="00:01:14.49" resultid="1366" heatid="2381" lane="2" entrytime="00:01:13.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Fonseca Vendramin" birthdate="2008-09-28" gender="F" nation="BRA" license="393918" swrid="5622282" athleteid="1373" externalid="393918">
              <RESULTS>
                <RESULT eventid="1060" points="412" swimtime="00:01:09.45" resultid="1374" heatid="2315" lane="3" entrytime="00:01:10.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Faria Del Valle" birthdate="2009-08-28" gender="M" nation="BRA" license="376328" swrid="5600155" athleteid="1343" externalid="376328">
              <RESULTS>
                <RESULT eventid="1068" points="546" swimtime="00:00:57.33" resultid="1344" heatid="2326" lane="4" entrytime="00:00:57.69" entrycourse="LCM" />
                <RESULT eventid="1196" points="436" swimtime="00:01:08.02" resultid="1345" heatid="2381" lane="4" entrytime="00:01:10.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Zaleski Dallazem" birthdate="2009-05-16" gender="M" nation="BRA" license="344286" swrid="5600280" athleteid="1337" externalid="344286">
              <RESULTS>
                <RESULT eventid="1084" points="415" swimtime="00:02:48.20" resultid="1338" heatid="2334" lane="7" entrytime="00:02:47.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="419" swimtime="00:01:15.98" resultid="1339" heatid="2392" lane="5" entrytime="00:01:15.53" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Inacio Carneiro" birthdate="2009-09-09" gender="M" nation="BRA" license="408023" swrid="5723026" athleteid="1383" externalid="408023">
              <RESULTS>
                <RESULT eventid="1068" points="336" swimtime="00:01:07.34" resultid="1384" heatid="2321" lane="1" entrytime="00:01:07.27" entrycourse="LCM" />
                <RESULT eventid="1164" points="278" swimtime="00:02:36.23" resultid="1385" heatid="2366" lane="6" entrytime="00:02:35.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.32" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Tempo: 17:40), Na volta dos 50m." eventid="1212" status="DSQ" swimtime="00:01:30.62" resultid="1386" heatid="2389" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="James" lastname="Roberto Zoschke" birthdate="1976-02-08" gender="M" nation="BRA" license="312251" swrid="5688617" athleteid="1332" externalid="312251">
              <RESULTS>
                <RESULT eventid="1212" points="421" swimtime="00:01:15.87" resultid="1333" heatid="2393" lane="8" entrytime="00:01:14.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Camila" lastname="Duarte De Almeida" birthdate="2009-11-26" gender="F" nation="BRA" license="378819" swrid="5600152" athleteid="1349" externalid="378819">
              <RESULTS>
                <RESULT eventid="1060" points="481" swimtime="00:01:05.97" resultid="1350" heatid="2317" lane="2" entrytime="00:01:06.30" entrycourse="LCM" />
                <RESULT eventid="1156" points="410" swimtime="00:02:31.81" resultid="1351" heatid="2362" lane="3" entrytime="00:02:30.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="1762" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Ribeiro Melo" birthdate="2011-07-01" gender="F" nation="BRA" license="390923" swrid="5602577" athleteid="1763" externalid="390923">
              <RESULTS>
                <RESULT eventid="1060" points="411" swimtime="00:01:09.51" resultid="1764" heatid="2316" lane="3" entrytime="00:01:08.22" entrycourse="LCM" />
                <RESULT eventid="1156" points="472" swimtime="00:02:24.92" resultid="1765" heatid="2362" lane="5" entrytime="00:02:29.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="311" swimtime="00:01:24.60" resultid="1766" heatid="2377" lane="2" entrytime="00:01:24.82" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Camillo Sabim" birthdate="2010-08-02" gender="F" nation="BRA" license="406931" swrid="5723021" athleteid="1782" externalid="406931">
              <RESULTS>
                <RESULT eventid="1060" points="311" swimtime="00:01:16.26" resultid="1783" heatid="2314" lane="3" entrytime="00:01:12.79" entrycourse="LCM" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Tempo: 9:51), Na volta dos 150m." eventid="1076" status="DSQ" swimtime="00:03:21.35" resultid="1784" heatid="2329" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="322" swimtime="00:01:33.47" resultid="1785" heatid="2385" lane="4" entrytime="00:01:34.67" entrycourse="LCM" />
                <RESULT eventid="1188" points="261" swimtime="00:01:29.70" resultid="1786" heatid="2376" lane="2" entrytime="00:01:31.53" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Guilherme Ballatka" birthdate="2007-06-24" gender="M" nation="BRA" license="398616" swrid="5697228" athleteid="1772" externalid="398616">
              <RESULTS>
                <RESULT eventid="1116" points="405" swimtime="00:02:31.15" resultid="1773" heatid="2344" lane="3" entrytime="00:02:41.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="468" swimtime="00:01:00.34" resultid="1774" heatid="2324" lane="6" entrytime="00:01:01.48" entrycourse="LCM" />
                <RESULT eventid="1164" points="390" swimtime="00:02:19.56" resultid="1775" heatid="2367" lane="1" entrytime="00:02:32.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="426" swimtime="00:01:08.57" resultid="1776" heatid="2382" lane="3" entrytime="00:01:07.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jennifer" lastname="De Abreu" birthdate="2009-11-07" gender="F" nation="BRA" license="356212" swrid="5600144" athleteid="1767" externalid="356212">
              <RESULTS>
                <RESULT eventid="1060" points="523" swimtime="00:01:04.15" resultid="1768" heatid="2318" lane="3" entrytime="00:01:03.67" entrycourse="LCM" />
                <RESULT eventid="1124" points="445" swimtime="00:01:12.63" resultid="1769" heatid="2348" lane="5" entrytime="00:01:12.89" entrycourse="LCM" />
                <RESULT eventid="1156" points="468" swimtime="00:02:25.31" resultid="1770" heatid="2364" lane="2" entrytime="00:02:19.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="371" swimtime="00:01:19.73" resultid="1771" heatid="2377" lane="5" entrytime="00:01:21.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucca" lastname="Diedrichs Santos" birthdate="2011-10-27" gender="M" nation="BRA" license="414417" swrid="5755372" athleteid="1787" externalid="414417">
              <RESULTS>
                <RESULT eventid="1068" points="144" swimtime="00:01:29.40" resultid="1788" heatid="2319" lane="2" />
                <RESULT eventid="1212" points="163" swimtime="00:01:43.93" resultid="1789" heatid="2389" lane="7" />
                <RESULT eventid="1196" points="167" swimtime="00:01:33.69" resultid="1790" heatid="2379" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Ferreira Rais" birthdate="2007-07-04" gender="M" nation="BRA" license="398656" swrid="5697227" athleteid="1777" externalid="398656">
              <RESULTS>
                <RESULT eventid="1132" points="255" swimtime="00:01:17.88" resultid="1778" heatid="2351" lane="3" entrytime="00:01:18.36" entrycourse="LCM" />
                <RESULT eventid="1068" points="410" swimtime="00:01:03.06" resultid="1779" heatid="2322" lane="2" entrytime="00:01:05.09" entrycourse="LCM" />
                <RESULT eventid="1164" points="324" swimtime="00:02:28.48" resultid="1780" heatid="2366" lane="5" entrytime="00:02:34.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="280" swimtime="00:01:18.87" resultid="1781" heatid="2380" lane="7" entrytime="00:01:25.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13068" nation="BRA" region="PR" clubid="1791" swrid="93787" name="Sociedade Morgenau" shortname="Morgenau">
          <ATHLETES>
            <ATHLETE firstname="Geovana" lastname="Dos Santos" birthdate="2011-01-20" gender="F" nation="BRA" license="367254" swrid="5602533" athleteid="1792" externalid="367254">
              <RESULTS>
                <RESULT eventid="1060" points="302" swimtime="00:01:16.99" resultid="1793" heatid="2314" lane="2" entrytime="00:01:15.96" entrycourse="LCM" />
                <RESULT eventid="1156" points="332" swimtime="00:02:42.86" resultid="1794" heatid="2361" lane="1" entrytime="00:02:45.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="299" swimtime="00:01:25.68" resultid="1795" heatid="2377" lane="7" entrytime="00:01:24.86" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Rodrigues Galvao" birthdate="2007-04-19" gender="M" nation="BRA" license="376586" swrid="5600247" athleteid="1796" externalid="376586">
              <RESULTS>
                <RESULT eventid="1132" points="463" swimtime="00:01:03.90" resultid="1797" heatid="2354" lane="7" entrytime="00:01:03.13" entrycourse="LCM" />
                <RESULT eventid="1068" points="526" swimtime="00:00:58.05" resultid="1798" heatid="2326" lane="6" entrytime="00:00:58.11" entrycourse="LCM" />
                <RESULT eventid="1164" points="468" swimtime="00:02:11.31" resultid="1799" heatid="2370" lane="2" entrytime="00:02:10.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaylane" lastname="Marques Ferreira" birthdate="2010-03-06" gender="F" nation="BRA" license="391146" swrid="5600211" athleteid="1878" externalid="391146">
              <RESULTS>
                <RESULT eventid="1060" points="308" swimtime="00:01:16.56" resultid="1879" heatid="2313" lane="4" entrytime="00:01:17.16" entrycourse="LCM" />
                <RESULT eventid="1124" points="248" swimtime="00:01:28.27" resultid="1880" heatid="2348" lane="6" entrytime="00:01:27.84" entrycourse="LCM" />
                <RESULT eventid="1156" points="266" swimtime="00:02:55.41" resultid="1881" heatid="2360" lane="5" entrytime="00:02:56.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="211" swimtime="00:01:36.19" resultid="1882" heatid="2375" lane="4" entrytime="00:01:47.27" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Andreis Ramos" birthdate="2007-03-26" gender="M" nation="BRA" license="406719" swrid="5717243" athleteid="1828" externalid="406719">
              <RESULTS>
                <RESULT eventid="1068" points="418" swimtime="00:01:02.66" resultid="1829" heatid="2323" lane="5" entrytime="00:01:03.03" entrycourse="LCM" />
                <RESULT eventid="1196" points="275" swimtime="00:01:19.26" resultid="1830" heatid="2380" lane="6" entrytime="00:01:20.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wilson" lastname="Soares Filho" birthdate="2007-12-20" gender="M" nation="BRA" license="414552" swrid="5755379" athleteid="1917" externalid="414552">
              <RESULTS>
                <RESULT eventid="1084" points="251" swimtime="00:03:18.84" resultid="1918" heatid="2332" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="351" swimtime="00:02:24.59" resultid="1919" heatid="2365" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="268" swimtime="00:01:28.16" resultid="1920" heatid="2391" lane="7" entrytime="00:01:26.44" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabryel" lastname="Denk" birthdate="2011-05-09" gender="M" nation="BRA" license="391138" swrid="5602531" athleteid="1867" externalid="391138">
              <RESULTS>
                <RESULT eventid="1116" points="308" swimtime="00:02:45.60" resultid="1868" heatid="2344" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="368" swimtime="00:10:30.80" resultid="1869" heatid="2340" lane="2" entrytime="00:10:26.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.37" />
                    <SPLIT distance="200" swimtime="00:02:32.31" />
                    <SPLIT distance="300" swimtime="00:03:52.55" />
                    <SPLIT distance="400" swimtime="00:05:12.16" />
                    <SPLIT distance="500" swimtime="00:06:32.76" />
                    <SPLIT distance="600" swimtime="00:07:53.30" />
                    <SPLIT distance="700" swimtime="00:09:13.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="333" swimtime="00:01:07.60" resultid="1870" heatid="2321" lane="6" entrytime="00:01:06.23" entrycourse="LCM" />
                <RESULT eventid="1164" points="343" swimtime="00:02:25.70" resultid="1871" heatid="2367" lane="3" entrytime="00:02:25.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="281" swimtime="00:01:18.77" resultid="1872" heatid="2380" lane="4" entrytime="00:01:17.10" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Andrianczik Corcini" birthdate="2008-07-19" gender="M" nation="BRA" license="406685" swrid="5736533" athleteid="1817" externalid="406685">
              <RESULTS>
                <RESULT eventid="1084" points="216" swimtime="00:03:29.06" resultid="1818" heatid="2332" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="338" swimtime="00:01:07.24" resultid="1819" heatid="2321" lane="8" entrytime="00:01:07.60" entrycourse="LCM" />
                <RESULT eventid="1164" points="252" swimtime="00:02:41.43" resultid="1820" heatid="2366" lane="7" entrytime="00:02:38.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.09" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada.  (Tempo: 17:43), Na volta dos 50m." eventid="1212" status="DSQ" swimtime="00:01:35.72" resultid="1821" heatid="2390" lane="6" entrytime="00:01:29.44" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thiago" lastname="Kozera Chiarato" birthdate="2008-01-22" gender="M" nation="BRA" license="406728" swrid="5717276" athleteid="1911" externalid="406728">
              <RESULTS>
                <RESULT eventid="1132" points="352" swimtime="00:01:09.99" resultid="1912" heatid="2353" lane="7" entrytime="00:01:09.31" entrycourse="LCM" />
                <RESULT eventid="1084" points="269" swimtime="00:03:14.27" resultid="1913" heatid="2333" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="475" swimtime="00:01:00.05" resultid="1914" heatid="2325" lane="8" entrytime="00:01:00.29" entrycourse="LCM" />
                <RESULT eventid="1148" points="314" swimtime="00:05:56.60" resultid="1915" heatid="2357" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.54" />
                    <SPLIT distance="200" swimtime="00:02:58.85" />
                    <SPLIT distance="300" swimtime="00:04:38.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="359" swimtime="00:01:19.97" resultid="1916" heatid="2392" lane="6" entrytime="00:01:17.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Henrique Opuchkevich" birthdate="2011-02-22" gender="M" nation="BRA" license="406720" swrid="5717273" athleteid="1899" externalid="406720">
              <RESULTS>
                <RESULT eventid="1100" points="374" swimtime="00:10:27.28" resultid="1900" heatid="2339" lane="6" entrytime="00:10:47.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                    <SPLIT distance="200" swimtime="00:02:32.96" />
                    <SPLIT distance="300" swimtime="00:03:52.21" />
                    <SPLIT distance="400" swimtime="00:05:12.07" />
                    <SPLIT distance="500" swimtime="00:06:31.94" />
                    <SPLIT distance="600" swimtime="00:07:52.54" />
                    <SPLIT distance="700" swimtime="00:09:11.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1084" points="340" swimtime="00:02:59.70" resultid="1901" heatid="2334" lane="8" entrytime="00:03:04.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="352" swimtime="00:02:24.40" resultid="1902" heatid="2366" lane="8" entrytime="00:02:46.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="327" swimtime="00:01:22.53" resultid="1903" heatid="2391" lane="3" entrytime="00:01:23.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kedny" lastname="Correa" birthdate="2004-11-05" gender="M" nation="BRA" license="383858" swrid="5600142" athleteid="1849" externalid="383858">
              <RESULTS>
                <RESULT eventid="1068" points="465" swimtime="00:01:00.46" resultid="1850" heatid="2325" lane="1" entrytime="00:01:00.11" entrycourse="LCM" />
                <RESULT eventid="1148" points="383" swimtime="00:05:33.84" resultid="1851" heatid="2357" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.15" />
                    <SPLIT distance="200" swimtime="00:02:49.13" />
                    <SPLIT distance="300" swimtime="00:04:19.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="287" swimtime="00:01:18.16" resultid="1852" heatid="2379" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauan" lastname="Araujo" birthdate="2009-12-17" gender="M" nation="BRA" license="385119" swrid="5653286" athleteid="1853" externalid="385119">
              <RESULTS>
                <RESULT eventid="1132" points="255" swimtime="00:01:17.91" resultid="1854" heatid="2350" lane="2" />
                <RESULT eventid="1100" points="362" swimtime="00:10:34.11" resultid="1855" heatid="2340" lane="7" entrytime="00:10:32.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.41" />
                    <SPLIT distance="200" swimtime="00:02:28.73" />
                    <SPLIT distance="300" swimtime="00:03:49.49" />
                    <SPLIT distance="400" swimtime="00:05:11.37" />
                    <SPLIT distance="500" swimtime="00:06:33.37" />
                    <SPLIT distance="600" swimtime="00:07:55.99" />
                    <SPLIT distance="700" swimtime="00:09:16.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="401" swimtime="00:01:03.53" resultid="1856" heatid="2323" lane="8" entrytime="00:01:03.96" entrycourse="LCM" />
                <RESULT eventid="1164" points="399" swimtime="00:02:18.45" resultid="1857" heatid="2368" lane="6" entrytime="00:02:20.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Rafaella Dos Santos" birthdate="2005-02-25" gender="F" nation="BRA" license="358849" swrid="5757094" athleteid="1800" externalid="358849">
              <RESULTS>
                <RESULT eventid="1076" points="298" swimtime="00:03:25.76" resultid="1801" heatid="2329" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="253" swimtime="00:02:58.34" resultid="1802" heatid="2360" lane="4" entrytime="00:02:56.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="305" swimtime="00:01:35.19" resultid="1803" heatid="2385" lane="3" entrytime="00:01:36.10" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Liz Skowronski" birthdate="2008-01-24" gender="F" nation="BRA" license="358245" swrid="5600202" athleteid="1804" externalid="358245">
              <RESULTS>
                <RESULT eventid="1060" points="380" swimtime="00:01:11.33" resultid="1805" heatid="2312" lane="3" />
                <RESULT eventid="1108" points="352" swimtime="00:02:54.37" resultid="1806" heatid="2342" lane="7" entrytime="00:02:50.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="369" swimtime="00:02:37.25" resultid="1807" heatid="2362" lane="2" entrytime="00:02:32.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="353" swimtime="00:01:21.11" resultid="1808" heatid="2378" lane="8" entrytime="00:01:19.56" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Mingorance Martins" birthdate="2007-10-13" gender="M" nation="BRA" license="393920" swrid="5622295" athleteid="1886" externalid="393920">
              <RESULTS>
                <RESULT eventid="1068" points="552" swimtime="00:00:57.11" resultid="1887" heatid="2327" lane="7" entrytime="00:00:56.90" entrycourse="LCM" />
                <RESULT eventid="1164" points="433" swimtime="00:02:14.81" resultid="1888" heatid="2371" lane="8" entrytime="00:02:08.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="356" swimtime="00:05:42.08" resultid="1889" heatid="2357" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.83" />
                    <SPLIT distance="200" swimtime="00:02:44.67" />
                    <SPLIT distance="300" swimtime="00:04:25.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Kozera Chiarato" birthdate="2010-05-28" gender="M" nation="BRA" license="406722" swrid="5717275" athleteid="1904" externalid="406722">
              <RESULTS>
                <RESULT eventid="1132" points="269" swimtime="00:01:16.52" resultid="1905" heatid="2352" lane="2" entrytime="00:01:13.56" entrycourse="LCM" />
                <RESULT eventid="1100" points="318" swimtime="00:11:02.21" resultid="1906" heatid="2338" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.38" />
                    <SPLIT distance="200" swimtime="00:02:38.91" />
                    <SPLIT distance="300" swimtime="00:04:04.99" />
                    <SPLIT distance="400" swimtime="00:05:30.63" />
                    <SPLIT distance="500" swimtime="00:06:56.43" />
                    <SPLIT distance="600" swimtime="00:08:21.89" />
                    <SPLIT distance="700" swimtime="00:09:44.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="377" swimtime="00:01:04.84" resultid="1907" heatid="2320" lane="4" entrytime="00:01:08.29" entrycourse="LCM" />
                <RESULT eventid="1180" points="199" swimtime="00:03:08.79" resultid="1908" heatid="2374" lane="1" entrytime="00:03:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karine" lastname="Correa" birthdate="2002-08-01" gender="F" nation="BRA" license="385191" swrid="5600141" athleteid="1822" externalid="385191">
              <RESULTS>
                <RESULT eventid="1060" points="359" swimtime="00:01:12.70" resultid="1823" heatid="2314" lane="4" entrytime="00:01:12.05" entrycourse="LCM" />
                <RESULT eventid="1092" points="281" swimtime="00:12:19.60" resultid="1824" heatid="2336" lane="3" entrytime="00:12:25.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.44" />
                    <SPLIT distance="200" swimtime="00:02:54.31" />
                    <SPLIT distance="300" swimtime="00:04:26.61" />
                    <SPLIT distance="400" swimtime="00:06:01.82" />
                    <SPLIT distance="500" swimtime="00:07:37.69" />
                    <SPLIT distance="600" swimtime="00:09:12.86" />
                    <SPLIT distance="700" swimtime="00:10:47.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="329" swimtime="00:02:43.45" resultid="1825" heatid="2361" lane="2" entrytime="00:02:42.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monike" lastname="Lemos Carvalho" birthdate="2008-03-28" gender="F" nation="BRA" license="307796" swrid="5600199" athleteid="1858" externalid="307796">
              <RESULTS>
                <RESULT eventid="1060" points="444" swimtime="00:01:07.74" resultid="1859" heatid="2317" lane="5" entrytime="00:01:06.06" entrycourse="LCM" />
                <RESULT eventid="1092" points="392" swimtime="00:11:01.88" resultid="1860" heatid="2336" lane="4" entrytime="00:11:05.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="200" swimtime="00:02:38.53" />
                    <SPLIT distance="300" swimtime="00:04:02.99" />
                    <SPLIT distance="400" swimtime="00:05:27.09" />
                    <SPLIT distance="500" swimtime="00:06:51.95" />
                    <SPLIT distance="600" swimtime="00:08:17.26" />
                    <SPLIT distance="700" swimtime="00:09:41.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="504" swimtime="00:02:21.77" resultid="1861" heatid="2363" lane="5" entrytime="00:02:24.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="410" swimtime="00:01:17.16" resultid="1862" heatid="2378" lane="7" entrytime="00:01:16.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Matos Oliveira" birthdate="2007-10-26" gender="M" nation="BRA" license="391136" swrid="5600215" athleteid="1863" externalid="391136">
              <RESULTS>
                <RESULT eventid="1100" points="294" swimtime="00:11:19.60" resultid="1864" heatid="2339" lane="2" entrytime="00:10:55.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.90" />
                    <SPLIT distance="200" swimtime="00:02:41.93" />
                    <SPLIT distance="300" swimtime="00:04:08.40" />
                    <SPLIT distance="400" swimtime="00:05:35.13" />
                    <SPLIT distance="500" swimtime="00:07:02.15" />
                    <SPLIT distance="600" swimtime="00:08:30.69" />
                    <SPLIT distance="700" swimtime="00:09:57.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="224" swimtime="00:06:38.71" resultid="1865" heatid="2358" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.66" />
                    <SPLIT distance="200" swimtime="00:03:14.79" />
                    <SPLIT distance="300" swimtime="00:05:11.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="139" swimtime="00:03:32.94" resultid="1866" heatid="2373" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Luiza Rimbano De Jesus" birthdate="2008-09-02" gender="F" nation="BRA" license="366819" swrid="5653297" athleteid="1890" externalid="366819">
              <RESULTS>
                <RESULT eventid="1060" points="555" swimtime="00:01:02.90" resultid="1891" heatid="2318" lane="5" entrytime="00:01:02.31" entrycourse="LCM" />
                <RESULT eventid="1156" points="473" swimtime="00:02:24.80" resultid="1892" heatid="2363" lane="4" entrytime="00:02:23.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="344" swimtime="00:01:21.82" resultid="1893" heatid="2375" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stella" lastname="Magalhaes Birnbaum" birthdate="2009-05-14" gender="F" nation="BRA" license="399684" swrid="5653298" athleteid="1894" externalid="399684">
              <RESULTS>
                <RESULT eventid="1060" points="391" swimtime="00:01:10.67" resultid="1895" heatid="2316" lane="7" entrytime="00:01:09.13" entrycourse="LCM" />
                <RESULT eventid="1108" points="375" swimtime="00:02:50.62" resultid="1896" heatid="2342" lane="1" entrytime="00:02:54.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="371" swimtime="00:02:37.05" resultid="1897" heatid="2361" lane="5" entrytime="00:02:35.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="389" swimtime="00:01:18.48" resultid="1898" heatid="2377" lane="4" entrytime="00:01:20.33" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mayara" lastname="Fieber" birthdate="2008-08-20" gender="F" nation="BRA" license="391147" swrid="5600161" athleteid="1883" externalid="391147">
              <RESULTS>
                <RESULT comment="SW 10.2 - Não completou a distância total da prova.  (Tempo: 12:07)" eventid="1124" status="DSQ" swimtime="00:00:00.00" resultid="1884" heatid="2348" lane="7" entrytime="00:01:32.14" entrycourse="LCM" />
                <RESULT eventid="1204" points="323" swimtime="00:01:33.44" resultid="1885" heatid="2384" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Vitor Navarro Zanini" birthdate="2008-06-30" gender="M" nation="BRA" license="369415" swrid="5600273" athleteid="1837" externalid="369415">
              <RESULTS>
                <RESULT eventid="1100" points="304" swimtime="00:11:12.16" resultid="1838" heatid="2339" lane="5" entrytime="00:10:36.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.40" />
                    <SPLIT distance="200" swimtime="00:02:42.73" />
                    <SPLIT distance="300" swimtime="00:04:08.01" />
                    <SPLIT distance="400" swimtime="00:05:34.06" />
                    <SPLIT distance="500" swimtime="00:06:58.21" />
                    <SPLIT distance="600" swimtime="00:08:22.51" />
                    <SPLIT distance="700" swimtime="00:09:48.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="280" swimtime="00:06:10.57" resultid="1839" heatid="2358" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.65" />
                    <SPLIT distance="200" swimtime="00:03:09.35" />
                    <SPLIT distance="300" swimtime="00:04:46.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="322" swimtime="00:01:22.92" resultid="1840" heatid="2392" lane="1" entrytime="00:01:18.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Fernanda Pinto" birthdate="2004-09-17" gender="F" nation="BRA" license="391144" swrid="5600157" athleteid="1826" externalid="391144">
              <RESULTS>
                <RESULT eventid="1060" points="350" swimtime="00:01:13.32" resultid="1827" heatid="2315" lane="1" entrytime="00:01:11.53" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduarda" lastname="Azevedo Birsneek" birthdate="2010-03-31" gender="F" nation="BRA" license="391145" swrid="5389427" athleteid="1873" externalid="391145">
              <RESULTS>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Tempo: 12:04), Na volta dos 50m. " eventid="1124" status="DSQ" swimtime="00:01:55.84" resultid="1874" heatid="2347" lane="6" entrytime="00:01:45.89" entrycourse="LCM" />
                <RESULT eventid="1108" points="248" swimtime="00:03:15.99" resultid="1875" heatid="2341" lane="2" entrytime="00:03:23.39" entrycourse="LCM" />
                <RESULT eventid="1156" points="199" swimtime="00:03:13.14" resultid="1876" heatid="2360" lane="6" entrytime="00:03:17.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="226" swimtime="00:01:34.10" resultid="1877" heatid="2376" lane="7" entrytime="00:01:36.29" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcus" lastname="Vinicius De Almeida" birthdate="2009-06-16" gender="M" nation="BRA" license="348099" swrid="5600272" athleteid="1831" externalid="348099">
              <RESULTS>
                <RESULT eventid="1164" points="471" swimtime="00:02:11.03" resultid="1832" heatid="2370" lane="1" entrytime="00:02:12.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="544" swimtime="00:01:09.65" resultid="1833" heatid="2393" lane="2" entrytime="00:01:09.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="De Mello Araujo" birthdate="2010-11-03" gender="F" nation="BRA" license="406723" swrid="5717254" athleteid="1909" externalid="406723">
              <RESULTS>
                <RESULT eventid="1060" points="279" swimtime="00:01:19.09" resultid="1910" heatid="2312" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benito" lastname="Alves Sant&apos;Ana" birthdate="2009-06-01" gender="M" nation="BRA" license="376585" swrid="5351951" athleteid="1809" externalid="376585">
              <RESULTS>
                <RESULT eventid="1116" points="433" swimtime="00:02:27.83" resultid="1810" heatid="2345" lane="1" entrytime="00:02:28.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="480" swimtime="00:00:59.82" resultid="1811" heatid="2319" lane="7" />
                <RESULT eventid="1180" points="411" swimtime="00:02:28.37" resultid="1812" heatid="2373" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Gabriel Sarmento Buski" birthdate="2010-04-05" gender="M" nation="BRA" license="399533" swrid="5717264" athleteid="1813" externalid="399533">
              <RESULTS>
                <RESULT eventid="1100" points="379" swimtime="00:10:24.66" resultid="1814" heatid="2340" lane="6" entrytime="00:10:22.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.54" />
                    <SPLIT distance="200" swimtime="00:02:27.96" />
                    <SPLIT distance="300" swimtime="00:03:46.98" />
                    <SPLIT distance="400" swimtime="00:05:07.53" />
                    <SPLIT distance="500" swimtime="00:06:26.72" />
                    <SPLIT distance="600" swimtime="00:07:46.76" />
                    <SPLIT distance="700" swimtime="00:09:07.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1084" points="340" swimtime="00:02:59.69" resultid="1815" heatid="2332" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="368" swimtime="00:01:19.31" resultid="1816" heatid="2392" lane="7" entrytime="00:01:18.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauren" lastname="Dziura" birthdate="2010-01-11" gender="F" nation="BRA" license="369416" swrid="5588668" athleteid="1841" externalid="369416">
              <RESULTS>
                <RESULT eventid="1108" points="320" swimtime="00:03:00.02" resultid="1842" heatid="2341" lane="5" entrytime="00:03:02.56" entrycourse="LCM" />
                <RESULT eventid="1092" points="389" swimtime="00:11:04.03" resultid="1843" heatid="2337" lane="7" entrytime="00:10:54.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.31" />
                    <SPLIT distance="200" swimtime="00:02:35.40" />
                    <SPLIT distance="300" swimtime="00:03:57.59" />
                    <SPLIT distance="400" swimtime="00:05:22.42" />
                    <SPLIT distance="500" swimtime="00:06:48.40" />
                    <SPLIT distance="600" swimtime="00:08:14.91" />
                    <SPLIT distance="700" swimtime="00:09:40.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="410" swimtime="00:02:31.82" resultid="1844" heatid="2363" lane="1" entrytime="00:02:28.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Lima" birthdate="2006-12-03" gender="M" nation="BRA" license="366749" swrid="5600201" athleteid="1845" externalid="366749">
              <RESULTS>
                <RESULT eventid="1132" points="509" swimtime="00:01:01.91" resultid="1846" heatid="2354" lane="6" entrytime="00:01:02.81" entrycourse="LCM" />
                <RESULT eventid="1068" points="608" swimtime="00:00:55.31" resultid="1847" heatid="2328" lane="8" entrytime="00:00:55.72" entrycourse="LCM" />
                <RESULT eventid="1148" points="423" swimtime="00:05:23.00" resultid="1848" heatid="2357" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.45" />
                    <SPLIT distance="200" swimtime="00:02:32.97" />
                    <SPLIT distance="300" swimtime="00:04:13.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Bora" birthdate="2005-01-06" gender="F" nation="BRA" license="358252" swrid="5600153" athleteid="1834" externalid="358252">
              <RESULTS>
                <RESULT eventid="1140" points="300" swimtime="00:06:36.85" resultid="1835" heatid="2356" lane="4" entrytime="00:06:30.45" entrycourse="LCM" />
                <RESULT eventid="1156" points="364" swimtime="00:02:37.99" resultid="1836" heatid="2361" lane="3" entrytime="00:02:39.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16830" nation="BRA" region="PR" clubid="1311" swrid="94883" name="Arenna Carvalho Ltda" shortname="Arenna Carvalho">
          <ATHLETES>
            <ATHLETE firstname="Pietro" lastname="Lobo Mussoi" birthdate="2008-07-05" gender="M" nation="BRA" license="398573" swrid="5658061" athleteid="1312" externalid="398573">
              <RESULTS>
                <RESULT eventid="1132" points="386" swimtime="00:01:07.91" resultid="1313" heatid="2350" lane="4" />
                <RESULT eventid="1100" points="326" swimtime="00:10:56.39" resultid="1314" heatid="2339" lane="1" entrytime="00:11:03.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.51" />
                    <SPLIT distance="200" swimtime="00:02:38.23" />
                    <SPLIT distance="300" swimtime="00:04:02.20" />
                    <SPLIT distance="500" swimtime="00:06:50.59" />
                    <SPLIT distance="600" swimtime="00:08:14.38" />
                    <SPLIT distance="700" swimtime="00:09:37.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="465" swimtime="00:01:00.47" resultid="1315" heatid="2325" lane="6" entrytime="00:00:59.59" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1007" nation="BRA" region="PR" clubid="1921" swrid="93785" name="Santa Mônica Clube De Campo" shortname="Santa Mônica">
          <ATHLETES>
            <ATHLETE firstname="Carol" lastname="Nalle Bejes" birthdate="2010-04-20" gender="F" nation="BRA" license="377315" swrid="5588824" athleteid="1989" externalid="377315">
              <RESULTS>
                <RESULT eventid="1060" points="434" swimtime="00:01:08.27" resultid="1990" heatid="2317" lane="7" entrytime="00:01:07.35" entrycourse="LCM" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Tempo: 10:06), Na volta dos 150m." eventid="1076" status="DSQ" swimtime="00:02:59.77" resultid="1991" heatid="2331" lane="6" entrytime="00:02:58.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="445" swimtime="00:01:23.96" resultid="1992" heatid="2387" lane="2" entrytime="00:01:23.13" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Leticia Durat" birthdate="2008-02-09" gender="F" nation="BRA" license="331636" swrid="5600200" athleteid="1931" externalid="331636">
              <RESULTS>
                <RESULT eventid="1076" points="287" swimtime="00:03:28.45" resultid="1932" heatid="2330" lane="7" entrytime="00:03:18.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="307" swimtime="00:01:35.05" resultid="1933" heatid="2386" lane="2" entrytime="00:01:31.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucca" lastname="Maceno Araujo" birthdate="2010-09-29" gender="M" nation="BRA" license="367056" swrid="5588788" athleteid="1963" externalid="367056">
              <RESULTS>
                <RESULT eventid="1132" points="426" swimtime="00:01:05.69" resultid="1964" heatid="2353" lane="5" entrytime="00:01:06.66" entrycourse="LCM" />
                <RESULT comment="SW 8.5 - Totalmente submerso durante o nado.  (Tempo: 17:00)" eventid="1180" status="DSQ" swimtime="00:02:42.46" resultid="1965" heatid="2374" lane="2" entrytime="00:02:37.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Araujo Felix" birthdate="2010-05-27" gender="F" nation="BRA" license="393157" swrid="5622260" athleteid="2015" externalid="393157">
              <RESULTS>
                <RESULT eventid="1060" points="413" swimtime="00:01:09.41" resultid="2016" heatid="2316" lane="8" entrytime="00:01:09.23" entrycourse="LCM" />
                <RESULT eventid="1156" points="421" swimtime="00:02:30.47" resultid="2017" heatid="2362" lane="6" entrytime="00:02:30.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="331" swimtime="00:01:22.83" resultid="2018" heatid="2376" lane="4" entrytime="00:01:29.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Breno" lastname="Borges Piekarzievicz" birthdate="2011-11-11" gender="M" nation="BRA" license="403144" swrid="5676295" athleteid="2004" externalid="403144">
              <RESULTS>
                <RESULT eventid="1068" points="206" swimtime="00:01:19.32" resultid="2005" heatid="2320" lane="8" entrytime="00:01:22.64" entrycourse="LCM" />
                <RESULT eventid="1212" points="147" swimtime="00:01:47.69" resultid="2006" heatid="2389" lane="4" entrytime="00:01:45.57" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Ieger" birthdate="2009-02-20" gender="M" nation="BRA" license="356888" swrid="5600180" athleteid="1946" externalid="356888">
              <RESULTS>
                <RESULT eventid="1068" points="479" swimtime="00:00:59.88" resultid="1947" heatid="2325" lane="4" entrytime="00:00:59.21" entrycourse="LCM" />
                <RESULT eventid="1212" points="382" swimtime="00:01:18.39" resultid="1948" heatid="2392" lane="3" entrytime="00:01:17.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Nalle Bejes" birthdate="2010-04-20" gender="F" nation="BRA" license="377323" swrid="5588826" athleteid="1993" externalid="377323">
              <RESULTS>
                <RESULT eventid="1124" points="247" swimtime="00:01:28.41" resultid="1994" heatid="2346" lane="4" />
                <RESULT eventid="1076" points="401" swimtime="00:03:06.46" resultid="1995" heatid="2330" lane="5" entrytime="00:03:08.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="416" swimtime="00:01:25.84" resultid="1996" heatid="2386" lane="4" entrytime="00:01:26.62" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Marques Machado" birthdate="2010-02-17" gender="M" nation="BRA" license="390918" swrid="5600212" athleteid="1997" externalid="390918">
              <RESULTS>
                <RESULT eventid="1132" points="277" swimtime="00:01:15.83" resultid="1998" heatid="2352" lane="6" entrytime="00:01:12.98" entrycourse="LCM" />
                <RESULT eventid="1100" points="385" swimtime="00:10:21.12" resultid="1999" heatid="2340" lane="1" entrytime="00:10:33.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.76" />
                    <SPLIT distance="200" swimtime="00:02:26.80" />
                    <SPLIT distance="300" swimtime="00:03:46.23" />
                    <SPLIT distance="400" swimtime="00:05:06.02" />
                    <SPLIT distance="500" swimtime="00:06:25.37" />
                    <SPLIT distance="600" swimtime="00:07:45.92" />
                    <SPLIT distance="700" swimtime="00:09:06.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="382" swimtime="00:02:20.56" resultid="2000" heatid="2368" lane="4" entrytime="00:02:19.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otto" lastname="Hedeke" birthdate="2011-03-24" gender="M" nation="BRA" license="372643" swrid="5588738" athleteid="1986" externalid="372643">
              <RESULTS>
                <RESULT eventid="1100" points="307" swimtime="00:11:10.20" resultid="1987" heatid="2339" lane="7" entrytime="00:10:55.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.85" />
                    <SPLIT distance="200" swimtime="00:02:42.13" />
                    <SPLIT distance="300" swimtime="00:04:07.14" />
                    <SPLIT distance="400" swimtime="00:05:34.06" />
                    <SPLIT distance="500" swimtime="00:06:58.10" />
                    <SPLIT distance="600" swimtime="00:08:21.63" />
                    <SPLIT distance="700" swimtime="00:09:47.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="196" swimtime="00:03:09.68" resultid="1988" heatid="2374" lane="8" entrytime="00:03:18.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Helena Vieira Jussen" birthdate="2011-12-29" gender="F" nation="BRA" license="372282" swrid="5588740" athleteid="1983" externalid="372282">
              <RESULTS>
                <RESULT eventid="1076" points="364" swimtime="00:03:12.64" resultid="1984" heatid="2330" lane="2" entrytime="00:03:16.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="381" swimtime="00:01:28.40" resultid="1985" heatid="2386" lane="3" entrytime="00:01:29.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Novakoski" birthdate="2009-03-05" gender="F" nation="BRA" license="339136" swrid="5600225" athleteid="1940" externalid="339136">
              <RESULTS>
                <RESULT eventid="1156" points="463" swimtime="00:02:25.84" resultid="1941" heatid="2363" lane="2" entrytime="00:02:27.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Zanardi" birthdate="2008-10-02" gender="F" nation="BRA" license="398572" swrid="5757089" athleteid="2029" externalid="398572">
              <RESULTS>
                <RESULT eventid="1188" points="243" swimtime="00:01:31.80" resultid="2030" heatid="2375" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Dallastra" birthdate="2010-08-21" gender="M" nation="BRA" license="408024" swrid="5723028" athleteid="2023" externalid="408024">
              <RESULTS>
                <RESULT eventid="1068" points="440" swimtime="00:01:01.59" resultid="2024" heatid="2324" lane="2" entrytime="00:01:01.77" entrycourse="LCM" />
                <RESULT eventid="1164" points="428" swimtime="00:02:15.34" resultid="2025" heatid="2369" lane="2" entrytime="00:02:16.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Giuseppe Bulla Lanaro" birthdate="2007-05-22" gender="M" nation="BRA" license="331630" swrid="5600174" athleteid="1922" externalid="331630">
              <RESULTS>
                <RESULT eventid="1068" points="637" swimtime="00:00:54.44" resultid="1923" heatid="2328" lane="3" entrytime="00:00:53.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diego" lastname="Brasil Caropreso" birthdate="2009-10-29" gender="M" nation="BRA" license="399502" swrid="5653287" athleteid="2011" externalid="399502">
              <RESULTS>
                <RESULT eventid="1132" points="227" swimtime="00:01:20.96" resultid="2012" heatid="2351" lane="5" entrytime="00:01:17.20" entrycourse="LCM" />
                <RESULT eventid="1068" points="443" swimtime="00:01:01.47" resultid="2013" heatid="2324" lane="3" entrytime="00:01:01.41" entrycourse="LCM" />
                <RESULT eventid="1164" points="393" swimtime="00:02:19.21" resultid="2014" heatid="2369" lane="7" entrytime="00:02:18.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="De Castro Paiva Maciel" birthdate="2008-04-10" gender="M" nation="BRA" license="378333" swrid="5622275" athleteid="1927" externalid="378333">
              <RESULTS>
                <RESULT eventid="1132" points="389" swimtime="00:01:07.74" resultid="1928" heatid="2354" lane="1" entrytime="00:01:05.10" entrycourse="LCM" />
                <RESULT eventid="1068" points="520" swimtime="00:00:58.27" resultid="1929" heatid="2326" lane="1" entrytime="00:00:58.79" entrycourse="LCM" />
                <RESULT eventid="1164" points="463" swimtime="00:02:11.82" resultid="1930" heatid="2370" lane="7" entrytime="00:02:11.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Augusto Vaz" birthdate="2011-06-25" gender="M" nation="BRA" license="401737" swrid="5661339" athleteid="2001" externalid="401737">
              <RESULTS>
                <RESULT eventid="1132" points="357" swimtime="00:01:09.67" resultid="2002" heatid="2353" lane="1" entrytime="00:01:10.05" entrycourse="LCM" />
                <RESULT eventid="1068" points="376" swimtime="00:01:04.87" resultid="2003" heatid="2322" lane="4" entrytime="00:01:04.03" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Celli Schneider" birthdate="2011-02-21" gender="M" nation="BRA" license="367055" swrid="5588587" athleteid="1959" externalid="367055">
              <RESULTS>
                <RESULT eventid="1068" points="395" swimtime="00:01:03.82" resultid="1960" heatid="2321" lane="4" entrytime="00:01:05.82" entrycourse="LCM" />
                <RESULT eventid="1148" points="382" swimtime="00:05:34.02" resultid="1961" heatid="2358" lane="5" entrytime="00:05:36.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.62" />
                    <SPLIT distance="200" swimtime="00:02:39.88" />
                    <SPLIT distance="300" swimtime="00:04:21.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="385" swimtime="00:01:10.89" resultid="1962" heatid="2381" lane="5" entrytime="00:01:11.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietra" lastname="Vitoria Paczrowski" birthdate="2009-08-12" gender="F" nation="BRA" license="351253" swrid="5600275" athleteid="1944" externalid="351253">
              <RESULTS>
                <RESULT eventid="1060" points="467" swimtime="00:01:06.65" resultid="1945" heatid="2317" lane="3" entrytime="00:01:06.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Marcos Morais" birthdate="2010-01-30" gender="M" nation="BRA" license="416736" swrid="5757093" athleteid="2026" externalid="416736">
              <RESULTS>
                <RESULT eventid="1084" points="286" swimtime="00:03:10.35" resultid="2027" heatid="2333" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="313" swimtime="00:01:23.76" resultid="2028" heatid="2391" lane="8" entrytime="00:01:27.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Vianna" birthdate="2011-01-31" gender="M" nation="BRA" license="371380" swrid="5588947" athleteid="1979" externalid="371380">
              <RESULTS>
                <RESULT eventid="1100" points="289" swimtime="00:11:23.52" resultid="1980" heatid="2339" lane="4" entrytime="00:10:35.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.68" />
                    <SPLIT distance="200" swimtime="00:02:49.15" />
                    <SPLIT distance="300" swimtime="00:04:17.52" />
                    <SPLIT distance="400" swimtime="00:05:44.92" />
                    <SPLIT distance="500" swimtime="00:07:11.70" />
                    <SPLIT distance="600" swimtime="00:08:39.08" />
                    <SPLIT distance="700" swimtime="00:10:03.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" status="DNS" swimtime="00:00:00.00" resultid="1981" heatid="2368" lane="3" entrytime="00:02:20.38" entrycourse="LCM" />
                <RESULT eventid="1180" status="DNS" swimtime="00:00:00.00" resultid="1982" heatid="2373" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Inoue Kuroda" birthdate="2009-04-18" gender="M" nation="BRA" license="324700" swrid="5600190" athleteid="1937" externalid="324700">
              <RESULTS>
                <RESULT eventid="1068" points="525" swimtime="00:00:58.06" resultid="1938" heatid="2327" lane="2" entrytime="00:00:56.78" entrycourse="LCM" />
                <RESULT eventid="1196" points="402" swimtime="00:01:09.90" resultid="1939" heatid="2382" lane="6" entrytime="00:01:07.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cardim Martins" birthdate="2010-09-01" gender="F" nation="BRA" license="390920" swrid="5600130" athleteid="2019" externalid="390920">
              <RESULTS>
                <RESULT eventid="1124" points="182" swimtime="00:01:37.82" resultid="2020" heatid="2346" lane="3" />
                <RESULT eventid="1108" points="335" swimtime="00:02:57.30" resultid="2021" heatid="2342" lane="8" entrytime="00:03:01.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="316" swimtime="00:01:24.11" resultid="2022" heatid="2377" lane="6" entrytime="00:01:24.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Bello Costa Lange" birthdate="2010-09-13" gender="M" nation="BRA" license="367152" swrid="5588547" athleteid="1969" externalid="367152">
              <RESULTS>
                <RESULT eventid="1084" points="365" swimtime="00:02:55.55" resultid="1970" heatid="2333" lane="6" entrytime="00:03:16.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="373" swimtime="00:05:36.87" resultid="1971" heatid="2358" lane="3" entrytime="00:05:43.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.10" />
                    <SPLIT distance="200" swimtime="00:02:46.02" />
                    <SPLIT distance="300" swimtime="00:04:20.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="364" swimtime="00:01:19.66" resultid="1972" heatid="2389" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabrizio" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="M" nation="BRA" license="344303" swrid="5559846" athleteid="1934" externalid="344303">
              <RESULTS>
                <RESULT eventid="1116" points="447" swimtime="00:02:26.31" resultid="1935" heatid="2343" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="474" swimtime="00:01:06.15" resultid="1936" heatid="2382" lane="5" entrytime="00:01:06.59" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emily" lastname="Sayuri Tangueria De Lima" birthdate="2010-06-11" gender="F" nation="BRA" license="367215" swrid="5588901" athleteid="1973" externalid="367215">
              <RESULTS>
                <RESULT eventid="1124" points="360" swimtime="00:01:17.92" resultid="1974" heatid="2348" lane="3" entrytime="00:01:15.89" entrycourse="LCM" />
                <RESULT eventid="1092" points="429" swimtime="00:10:42.53" resultid="1975" heatid="2337" lane="1" entrytime="00:10:54.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.83" />
                    <SPLIT distance="200" swimtime="00:02:35.50" />
                    <SPLIT distance="300" swimtime="00:03:56.06" />
                    <SPLIT distance="400" swimtime="00:05:18.68" />
                    <SPLIT distance="500" swimtime="00:06:39.49" />
                    <SPLIT distance="600" swimtime="00:08:01.61" />
                    <SPLIT distance="700" swimtime="00:09:23.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="334" swimtime="00:02:55.52" resultid="1976" heatid="2372" lane="4" entrytime="00:02:53.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Cavassin Ieger" birthdate="2011-08-31" gender="M" nation="BRA" license="367149" swrid="5588743" athleteid="1966" externalid="367149">
              <RESULTS>
                <RESULT eventid="1084" points="309" swimtime="00:03:05.44" resultid="1967" heatid="2333" lane="5" entrytime="00:03:10.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="302" swimtime="00:01:24.76" resultid="1968" heatid="2390" lane="5" entrytime="00:01:28.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Analyce" lastname="Nunes Porto Luz" birthdate="2006-10-29" gender="F" nation="BRA" license="369322" swrid="5600226" athleteid="1924" externalid="369322">
              <RESULTS>
                <RESULT eventid="1124" points="447" swimtime="00:01:12.52" resultid="1925" heatid="2348" lane="4" entrytime="00:01:11.64" entrycourse="LCM" />
                <RESULT eventid="1156" points="536" swimtime="00:02:18.85" resultid="1926" heatid="2364" lane="6" entrytime="00:02:17.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Garcia Reschetti Rubbo" birthdate="2011-08-06" gender="F" nation="BRA" license="367053" swrid="5588720" athleteid="1955" externalid="367053">
              <RESULTS>
                <RESULT eventid="1124" points="194" swimtime="00:01:35.72" resultid="1956" heatid="2347" lane="8" />
                <RESULT eventid="1076" points="337" swimtime="00:03:17.56" resultid="1957" heatid="2330" lane="6" entrytime="00:03:15.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="318" swimtime="00:01:33.94" resultid="1958" heatid="2386" lane="7" entrytime="00:01:31.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kethelyn" lastname="Ribeiro Rodrigues" birthdate="2009-04-24" gender="F" nation="BRA" license="367052" swrid="5600244" athleteid="1952" externalid="367052">
              <RESULTS>
                <RESULT eventid="1060" points="428" swimtime="00:01:08.57" resultid="1953" heatid="2317" lane="1" entrytime="00:01:07.61" entrycourse="LCM" />
                <RESULT eventid="1156" points="412" swimtime="00:02:31.59" resultid="1954" heatid="2362" lane="4" entrytime="00:02:29.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="Moreira Furtado" birthdate="2011-01-27" gender="F" nation="BRA" license="403783" swrid="5684587" athleteid="2007" externalid="403783">
              <RESULTS>
                <RESULT eventid="1060" points="267" swimtime="00:01:20.28" resultid="2008" heatid="2314" lane="8" entrytime="00:01:16.91" entrycourse="LCM" />
                <RESULT eventid="1092" points="254" swimtime="00:12:45.16" resultid="2009" heatid="2335" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.83" />
                    <SPLIT distance="200" swimtime="00:03:01.24" />
                    <SPLIT distance="300" swimtime="00:04:38.49" />
                    <SPLIT distance="400" swimtime="00:06:16.63" />
                    <SPLIT distance="500" swimtime="00:07:55.06" />
                    <SPLIT distance="600" swimtime="00:09:33.98" />
                    <SPLIT distance="700" swimtime="00:11:11.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="213" swimtime="00:01:35.91" resultid="2010" heatid="2376" lane="1" entrytime="00:01:36.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Pinterich Almeida" birthdate="2005-03-13" gender="M" nation="BRA" license="330749" swrid="5600235" athleteid="1949" externalid="330749">
              <RESULTS>
                <RESULT eventid="1132" points="552" swimtime="00:01:00.27" resultid="1950" heatid="2354" lane="4" entrytime="00:01:01.00" entrycourse="LCM" />
                <RESULT eventid="1068" points="635" swimtime="00:00:54.50" resultid="1951" heatid="2328" lane="5" entrytime="00:00:53.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Gelenski Pelaio" birthdate="2005-10-10" gender="M" nation="BRA" license="281473" swrid="5600173" athleteid="1977" externalid="281473">
              <RESULTS>
                <RESULT eventid="1132" points="534" swimtime="00:01:00.95" resultid="1978" heatid="2355" lane="1" entrytime="00:01:00.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Blansky Hagebock" birthdate="2008-08-15" gender="M" nation="BRA" license="339123" swrid="5455418" athleteid="1942" externalid="339123">
              <RESULTS>
                <RESULT eventid="1068" points="563" swimtime="00:00:56.75" resultid="1943" heatid="2327" lane="5" entrytime="00:00:56.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16131" nation="BRA" region="PR" clubid="1736" swrid="93766" name="Associação Nadar Colombo" shortname="Equipe Nadar">
          <ATHLETES>
            <ATHLETE firstname="Lara" lastname="Carvalho Ezaki" birthdate="2011-10-20" gender="F" nation="BRA" license="399927" swrid="5652882" athleteid="1752" externalid="399927">
              <RESULTS>
                <RESULT eventid="1124" points="145" swimtime="00:01:45.57" resultid="1753" heatid="2347" lane="3" entrytime="00:01:45.68" entrycourse="LCM" />
                <RESULT eventid="1140" points="233" swimtime="00:07:11.72" resultid="1754" heatid="2356" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Guarise" birthdate="2008-11-28" gender="M" nation="BRA" license="408881" swrid="5727650" athleteid="1757" externalid="408881">
              <RESULTS>
                <RESULT eventid="1068" points="349" swimtime="00:01:06.50" resultid="1758" heatid="2322" lane="5" entrytime="00:01:04.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Luiz Sartori" birthdate="2008-04-07" gender="M" nation="BRA" license="384742" swrid="5622287" athleteid="1742" externalid="384742">
              <RESULTS>
                <RESULT eventid="1068" points="494" swimtime="00:00:59.26" resultid="1743" heatid="2325" lane="5" entrytime="00:00:59.28" entrycourse="LCM" />
                <RESULT eventid="1164" points="434" swimtime="00:02:14.63" resultid="1744" heatid="2369" lane="5" entrytime="00:02:15.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="348" swimtime="00:01:13.29" resultid="1745" heatid="2381" lane="7" entrytime="00:01:15.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaylaine" lastname="Sofia Vargas Bueno" birthdate="2006-11-28" gender="F" nation="BRA" license="384739" swrid="5622307" athleteid="1739" externalid="384739">
              <RESULTS>
                <RESULT eventid="1156" points="272" swimtime="00:02:53.97" resultid="1740" heatid="2361" lane="8" entrytime="00:02:48.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="230" swimtime="00:01:44.58" resultid="1741" heatid="2385" lane="2" entrytime="00:01:42.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Marcelo Santos Poli" birthdate="2007-09-01" gender="M" nation="BRA" license="388175" swrid="5622292" athleteid="1746" externalid="388175">
              <RESULTS>
                <RESULT eventid="1116" points="284" swimtime="00:02:50.11" resultid="1747" heatid="2344" lane="1" entrytime="00:02:46.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="425" swimtime="00:01:02.30" resultid="1748" heatid="2319" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Santos Poli" birthdate="2010-02-19" gender="M" nation="BRA" license="414563" swrid="5755378" athleteid="1759" externalid="414563">
              <RESULTS>
                <RESULT eventid="1132" points="227" swimtime="00:01:21.00" resultid="1760" heatid="2351" lane="6" entrytime="00:01:21.07" entrycourse="LCM" />
                <RESULT eventid="1068" points="328" swimtime="00:01:07.88" resultid="1761" heatid="2319" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Rafael D Agostin Batistao" birthdate="2008-05-13" gender="M" nation="BRA" license="384738" swrid="5622300" athleteid="1737" externalid="384738">
              <RESULTS>
                <RESULT eventid="1068" points="350" swimtime="00:01:06.44" resultid="1738" heatid="2322" lane="1" entrytime="00:01:05.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Krik" birthdate="2010-11-24" gender="F" nation="BRA" license="406702" swrid="5717277" athleteid="1755" externalid="406702">
              <RESULTS>
                <RESULT eventid="1092" points="167" swimtime="00:14:38.73" resultid="1756" heatid="2335" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:41.42" />
                    <SPLIT distance="200" swimtime="00:03:31.36" />
                    <SPLIT distance="300" swimtime="00:05:21.14" />
                    <SPLIT distance="400" swimtime="00:07:13.85" />
                    <SPLIT distance="500" swimtime="00:09:06.50" />
                    <SPLIT distance="600" swimtime="00:10:58.80" />
                    <SPLIT distance="700" swimtime="00:12:51.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Rosa De Souza" birthdate="2009-01-01" gender="F" nation="BRA" license="399926" swrid="5653301" athleteid="1749" externalid="399926">
              <RESULTS>
                <RESULT eventid="1124" points="124" swimtime="00:01:51.22" resultid="1750" heatid="2348" lane="1" entrytime="00:01:36.12" entrycourse="LCM" />
                <RESULT eventid="1092" points="198" swimtime="00:13:51.69" resultid="1751" heatid="2336" lane="2" entrytime="00:13:34.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.19" />
                    <SPLIT distance="200" swimtime="00:03:21.95" />
                    <SPLIT distance="300" swimtime="00:05:07.87" />
                    <SPLIT distance="400" swimtime="00:06:54.05" />
                    <SPLIT distance="500" swimtime="00:08:41.75" />
                    <SPLIT distance="600" swimtime="00:10:27.58" />
                    <SPLIT distance="700" swimtime="00:12:14.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="263" nation="BRA" region="PR" clubid="1443" swrid="75436" name="Clube Curitibano" shortname="Curitibano">
          <ATHLETES>
            <ATHLETE firstname="Joao" lastname="Pedro Kirchgassner" birthdate="2007-02-10" gender="M" nation="BRA" license="313535" swrid="5600230" athleteid="1485" externalid="313535">
              <RESULTS>
                <RESULT eventid="1084" points="633" swimtime="00:02:26.11" resultid="1486" heatid="2334" lane="4" entrytime="00:02:21.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="543" swimtime="00:02:05.00" resultid="1487" heatid="2371" lane="7" entrytime="00:02:04.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="562" swimtime="00:01:08.92" resultid="1488" heatid="2393" lane="5" entrytime="00:01:05.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Novak Bredt" birthdate="2009-09-08" gender="F" nation="BRA" license="338909" swrid="5622297" athleteid="1474" externalid="338909">
              <RESULTS>
                <RESULT eventid="1124" points="383" swimtime="00:01:16.38" resultid="1475" heatid="2347" lane="7" />
                <RESULT eventid="1204" points="419" swimtime="00:01:25.70" resultid="1476" heatid="2388" lane="8" entrytime="00:01:21.28" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Araujo Barros" birthdate="2008-12-26" gender="M" nation="BRA" license="331713" swrid="5367497" athleteid="1639" externalid="331713">
              <RESULTS>
                <RESULT eventid="1132" points="461" swimtime="00:01:04.00" resultid="1640" heatid="2349" lane="5" />
                <RESULT eventid="1068" points="585" swimtime="00:00:56.00" resultid="1641" heatid="2328" lane="1" entrytime="00:00:55.32" entrycourse="LCM" />
                <RESULT eventid="1164" points="591" swimtime="00:02:01.48" resultid="1642" heatid="2371" lane="4" entrytime="00:02:00.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="395" swimtime="00:01:17.48" resultid="1643" heatid="2389" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Peret Saboia" birthdate="2009-11-25" gender="F" nation="BRA" license="342238" swrid="5600234" athleteid="1507" externalid="342238">
              <RESULTS>
                <RESULT eventid="1060" points="468" swimtime="00:01:06.59" resultid="1508" heatid="2312" lane="4" />
                <RESULT eventid="1204" points="501" swimtime="00:01:20.70" resultid="1509" heatid="2388" lane="3" entrytime="00:01:18.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Correa Nascimento" birthdate="2009-01-19" gender="M" nation="BRA" license="342235" swrid="5600140" athleteid="1504" externalid="342235">
              <RESULTS>
                <RESULT eventid="1100" points="423" swimtime="00:10:02.05" resultid="1505" heatid="2338" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.44" />
                    <SPLIT distance="200" swimtime="00:02:21.54" />
                    <SPLIT distance="300" swimtime="00:03:36.06" />
                    <SPLIT distance="400" swimtime="00:04:50.04" />
                    <SPLIT distance="500" swimtime="00:06:10.40" />
                    <SPLIT distance="600" swimtime="00:07:29.87" />
                    <SPLIT distance="700" swimtime="00:08:48.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="471" swimtime="00:02:11.05" resultid="1506" heatid="2370" lane="4" entrytime="00:02:09.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Estela" lastname="Albuquerque" birthdate="2010-11-23" gender="F" nation="BRA" license="356344" swrid="5653285" athleteid="1549" externalid="356344">
              <RESULTS>
                <RESULT eventid="1060" points="470" swimtime="00:01:06.47" resultid="1550" heatid="2317" lane="6" entrytime="00:01:06.21" entrycourse="LCM" />
                <RESULT eventid="1124" points="289" swimtime="00:01:23.84" resultid="1551" heatid="2346" lane="6" />
                <RESULT eventid="1156" points="481" swimtime="00:02:24.02" resultid="1552" heatid="2364" lane="7" entrytime="00:02:21.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Zaroni" birthdate="2010-03-03" gender="F" nation="BRA" license="356345" swrid="5600282" athleteid="1470" externalid="356345">
              <RESULTS>
                <RESULT eventid="1060" points="432" swimtime="00:01:08.38" resultid="1471" heatid="2318" lane="8" entrytime="00:01:05.65" entrycourse="LCM" />
                <RESULT eventid="1076" points="428" swimtime="00:03:02.48" resultid="1472" heatid="2331" lane="3" entrytime="00:02:56.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="425" swimtime="00:01:25.23" resultid="1473" heatid="2387" lane="4" entrytime="00:01:22.19" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Leao" birthdate="2011-09-18" gender="M" nation="BRA" license="366880" swrid="5602553" athleteid="1580" externalid="366880">
              <RESULTS>
                <RESULT eventid="1132" points="279" swimtime="00:01:15.64" resultid="1581" heatid="2351" lane="2" entrytime="00:01:21.13" entrycourse="LCM" />
                <RESULT eventid="1068" points="393" swimtime="00:01:03.97" resultid="1582" heatid="2323" lane="7" entrytime="00:01:03.71" entrycourse="LCM" />
                <RESULT eventid="1164" points="407" swimtime="00:02:17.60" resultid="1583" heatid="2369" lane="1" entrytime="00:02:19.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Kraemer Geremia" birthdate="2011-07-20" gender="F" nation="BRA" license="366908" swrid="5588763" athleteid="1627" externalid="366908">
              <RESULTS>
                <RESULT eventid="1108" points="409" swimtime="00:02:45.84" resultid="1628" heatid="2342" lane="3" entrytime="00:02:39.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1092" points="450" swimtime="00:10:32.25" resultid="1629" heatid="2337" lane="6" entrytime="00:10:28.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.23" />
                    <SPLIT distance="200" swimtime="00:02:34.09" />
                    <SPLIT distance="300" swimtime="00:03:54.81" />
                    <SPLIT distance="400" swimtime="00:05:15.55" />
                    <SPLIT distance="500" swimtime="00:06:35.86" />
                    <SPLIT distance="600" swimtime="00:07:55.63" />
                    <SPLIT distance="700" swimtime="00:09:14.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="494" swimtime="00:02:22.70" resultid="1630" heatid="2364" lane="1" entrytime="00:02:22.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="346" swimtime="00:01:31.30" resultid="1631" heatid="2386" lane="8" entrytime="00:01:34.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Cury" birthdate="2005-09-28" gender="M" nation="BRA" license="329251" swrid="5600270" athleteid="1577" externalid="329251">
              <RESULTS>
                <RESULT eventid="1132" points="619" swimtime="00:00:58.00" resultid="1578" heatid="2355" lane="6" entrytime="00:00:57.21" entrycourse="LCM" />
                <RESULT eventid="1180" points="620" swimtime="00:02:09.34" resultid="1579" heatid="2374" lane="5" entrytime="00:02:08.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Vitoria Kuzmann Cercal" birthdate="2009-04-10" gender="F" nation="BRA" license="339082" swrid="5600274" athleteid="1517" externalid="339082">
              <RESULTS>
                <RESULT eventid="1060" points="524" swimtime="00:01:04.11" resultid="1518" heatid="2318" lane="2" entrytime="00:01:04.58" entrycourse="LCM" />
                <RESULT eventid="1188" points="418" swimtime="00:01:16.64" resultid="1519" heatid="2378" lane="6" entrytime="00:01:15.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Artigas Pinheiro" birthdate="2011-08-25" gender="M" nation="BRA" license="377040" swrid="5588535" athleteid="1666" externalid="377040">
              <RESULTS>
                <RESULT eventid="1084" points="340" swimtime="00:02:59.68" resultid="1667" heatid="2333" lane="4" entrytime="00:03:04.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="300" swimtime="00:06:02.07" resultid="1668" heatid="2357" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.12" />
                    <SPLIT distance="200" swimtime="00:03:02.31" />
                    <SPLIT distance="300" swimtime="00:04:38.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="310" swimtime="00:01:23.96" resultid="1669" heatid="2391" lane="2" entrytime="00:01:24.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Kremer De Aguiar" birthdate="2009-12-22" gender="F" nation="BRA" license="338987" swrid="5600196" athleteid="1510" externalid="338987">
              <RESULTS>
                <RESULT eventid="1060" points="447" swimtime="00:01:07.62" resultid="1511" heatid="2312" lane="5" />
                <RESULT eventid="1076" points="393" swimtime="00:03:07.77" resultid="1512" heatid="2330" lane="4" entrytime="00:03:02.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="437" swimtime="00:01:24.47" resultid="1513" heatid="2387" lane="6" entrytime="00:01:23.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ferreira Motta" birthdate="2008-10-24" gender="M" nation="BRA" license="378068" swrid="5600160" athleteid="1670" externalid="378068">
              <RESULTS>
                <RESULT eventid="1084" points="450" swimtime="00:02:43.69" resultid="1671" heatid="2334" lane="2" entrytime="00:02:42.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="422" swimtime="00:01:15.81" resultid="1672" heatid="2392" lane="4" entrytime="00:01:14.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="De Krinski" birthdate="2007-07-20" gender="M" nation="BRA" license="334494" swrid="5600148" athleteid="1711" externalid="334494">
              <RESULTS>
                <RESULT eventid="1116" points="476" swimtime="00:02:23.27" resultid="1712" heatid="2345" lane="3" entrytime="00:02:17.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="534" swimtime="00:01:03.58" resultid="1713" heatid="2383" lane="6" entrytime="00:01:01.36" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Clivatti" birthdate="2010-05-24" gender="M" nation="BRA" license="368007" swrid="5600139" athleteid="1444" externalid="368007">
              <RESULTS>
                <RESULT eventid="1068" points="537" swimtime="00:00:57.62" resultid="1445" heatid="2326" lane="5" entrytime="00:00:57.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Fantin Dias De Andrade" birthdate="2010-11-06" gender="F" nation="BRA" license="339262" swrid="5588684" athleteid="1649" externalid="339262">
              <RESULTS>
                <RESULT eventid="1124" points="211" swimtime="00:01:33.07" resultid="1650" heatid="2348" lane="2" entrytime="00:01:30.33" entrycourse="LCM" />
                <RESULT eventid="1156" points="345" swimtime="00:02:40.86" resultid="1651" heatid="2359" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="295" swimtime="00:01:36.28" resultid="1652" heatid="2385" lane="5" entrytime="00:01:35.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Rocha" birthdate="2011-08-25" gender="F" nation="BRA" license="366904" swrid="5602578" athleteid="1615" externalid="366904">
              <RESULTS>
                <RESULT eventid="1060" points="482" swimtime="00:01:05.93" resultid="1616" heatid="2318" lane="7" entrytime="00:01:05.12" entrycourse="LCM" />
                <RESULT eventid="1092" points="422" swimtime="00:10:45.82" resultid="1617" heatid="2337" lane="8" entrytime="00:11:05.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.38" />
                    <SPLIT distance="200" swimtime="00:02:37.11" />
                    <SPLIT distance="300" swimtime="00:03:58.36" />
                    <SPLIT distance="400" swimtime="00:05:18.92" />
                    <SPLIT distance="500" swimtime="00:06:39.68" />
                    <SPLIT distance="600" swimtime="00:08:02.19" />
                    <SPLIT distance="700" swimtime="00:09:25.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="480" swimtime="00:02:24.04" resultid="1618" heatid="2364" lane="8" entrytime="00:02:23.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorena" lastname="Mascarenhas" birthdate="2011-08-31" gender="F" nation="BRA" license="370581" swrid="5602558" athleteid="1653" externalid="370581">
              <RESULTS>
                <RESULT eventid="1060" points="426" swimtime="00:01:08.67" resultid="1654" heatid="2316" lane="5" entrytime="00:01:08.03" entrycourse="LCM" />
                <RESULT eventid="1156" points="409" swimtime="00:02:31.93" resultid="1655" heatid="2363" lane="8" entrytime="00:02:28.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="342" swimtime="00:01:31.69" resultid="1656" heatid="2386" lane="6" entrytime="00:01:31.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Fontolan Gomes" birthdate="2008-05-01" gender="M" nation="BRA" license="307667" swrid="5600166" athleteid="1489" externalid="307667">
              <RESULTS>
                <RESULT eventid="1132" status="DNS" swimtime="00:00:00.00" resultid="1490" heatid="2353" lane="3" entrytime="00:01:07.76" entrycourse="LCM" />
                <RESULT eventid="1116" points="407" swimtime="00:02:31.00" resultid="1491" heatid="2345" lane="7" entrytime="00:02:28.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="430" swimtime="00:01:08.34" resultid="1492" heatid="2382" lane="7" entrytime="00:01:08.13" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Cristina Ferreira" birthdate="2011-08-24" gender="F" nation="BRA" license="358334" swrid="5588611" athleteid="1446" externalid="358334">
              <RESULTS>
                <RESULT eventid="1204" points="482" swimtime="00:01:21.78" resultid="1447" heatid="2388" lane="6" entrytime="00:01:18.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="LIV" lastname="Carvalho" birthdate="2011-09-13" gender="F" nation="BRA" license="366899" swrid="5602524" athleteid="1603" externalid="366899">
              <RESULTS>
                <RESULT eventid="1092" points="315" swimtime="00:11:52.38" resultid="1604" heatid="2336" lane="5" entrytime="00:11:35.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.54" />
                    <SPLIT distance="200" swimtime="00:02:48.35" />
                    <SPLIT distance="300" swimtime="00:04:17.93" />
                    <SPLIT distance="400" swimtime="00:05:49.71" />
                    <SPLIT distance="500" swimtime="00:07:21.34" />
                    <SPLIT distance="600" swimtime="00:08:54.13" />
                    <SPLIT distance="700" swimtime="00:10:25.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="367" swimtime="00:02:37.49" resultid="1605" heatid="2361" lane="4" entrytime="00:02:35.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="221" swimtime="00:01:34.82" resultid="1606" heatid="2375" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Presiazniuk" birthdate="2010-10-14" gender="M" nation="BRA" license="356353" swrid="5600237" athleteid="1553" externalid="356353">
              <RESULTS>
                <RESULT eventid="1132" points="269" swimtime="00:01:16.53" resultid="1554" heatid="2350" lane="7" />
                <RESULT eventid="1068" points="501" swimtime="00:00:58.99" resultid="1555" heatid="2326" lane="2" entrytime="00:00:58.24" entrycourse="LCM" />
                <RESULT eventid="1196" points="402" swimtime="00:01:09.86" resultid="1556" heatid="2382" lane="1" entrytime="00:01:08.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Coelho" birthdate="2011-11-11" gender="M" nation="BRA" license="366889" swrid="5602527" athleteid="1584" externalid="366889">
              <RESULTS>
                <RESULT eventid="1132" points="325" swimtime="00:01:11.90" resultid="1585" heatid="2353" lane="8" entrytime="00:01:10.18" entrycourse="LCM" />
                <RESULT eventid="1068" points="376" swimtime="00:01:04.89" resultid="1586" heatid="2322" lane="6" entrytime="00:01:04.81" entrycourse="LCM" />
                <RESULT eventid="1164" points="390" swimtime="00:02:19.52" resultid="1587" heatid="2369" lane="8" entrytime="00:02:19.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Felipe Paes Feres" birthdate="2008-07-28" gender="M" nation="BRA" license="307676" swrid="5600156" athleteid="1493" externalid="307676">
              <RESULTS>
                <RESULT eventid="1116" points="422" swimtime="00:02:29.20" resultid="1494" heatid="2345" lane="6" entrytime="00:02:23.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="425" swimtime="00:01:08.60" resultid="1495" heatid="2382" lane="4" entrytime="00:01:06.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Schiavon" birthdate="2010-05-03" gender="M" nation="BRA" license="356354" swrid="5600256" athleteid="1557" externalid="356354">
              <RESULTS>
                <RESULT eventid="1116" points="402" swimtime="00:02:31.57" resultid="1558" heatid="2345" lane="8" entrytime="00:02:31.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="481" swimtime="00:02:10.10" resultid="1559" heatid="2370" lane="6" entrytime="00:02:10.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="435" swimtime="00:05:19.94" resultid="1560" heatid="2358" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                    <SPLIT distance="200" swimtime="00:02:36.96" />
                    <SPLIT distance="300" swimtime="00:04:09.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gael" lastname="Gluck" birthdate="2011-01-28" gender="M" nation="BRA" license="366891" swrid="5588726" athleteid="1588" externalid="366891">
              <RESULTS>
                <RESULT eventid="1084" points="369" swimtime="00:02:54.86" resultid="1589" heatid="2334" lane="1" entrytime="00:02:48.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="418" swimtime="00:01:02.66" resultid="1590" heatid="2324" lane="8" entrytime="00:01:02.75" entrycourse="LCM" />
                <RESULT eventid="1212" points="378" swimtime="00:01:18.66" resultid="1591" heatid="2392" lane="2" entrytime="00:01:18.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Carneiro Silva" birthdate="2011-02-21" gender="F" nation="BRA" license="390924" swrid="5602522" athleteid="1693" externalid="390924">
              <RESULTS>
                <RESULT eventid="1060" points="439" swimtime="00:01:08.01" resultid="1694" heatid="2315" lane="6" entrytime="00:01:10.50" entrycourse="LCM" />
                <RESULT eventid="1124" points="157" swimtime="00:01:42.72" resultid="1695" heatid="2347" lane="5" entrytime="00:01:44.66" entrycourse="LCM" />
                <RESULT eventid="1156" points="425" swimtime="00:02:30.02" resultid="1696" heatid="2361" lane="6" entrytime="00:02:42.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Saboia" birthdate="2009-01-25" gender="M" nation="BRA" license="342252" swrid="5600253" athleteid="1514" externalid="342252">
              <RESULTS>
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Tempo: 10:15), Na volta dos 150m." eventid="1084" status="DSQ" swimtime="00:02:40.40" resultid="1515" heatid="2334" lane="6" entrytime="00:02:40.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="468" swimtime="00:01:13.21" resultid="1516" heatid="2393" lane="1" entrytime="00:01:12.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fernandes" birthdate="2010-03-13" gender="M" nation="BRA" license="339266" swrid="5588695" athleteid="1687" externalid="339266">
              <RESULTS>
                <RESULT eventid="1116" points="433" swimtime="00:02:27.85" resultid="1688" heatid="2345" lane="2" entrytime="00:02:28.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="515" swimtime="00:00:58.45" resultid="1689" heatid="2327" lane="1" entrytime="00:00:57.58" entrycourse="LCM" />
                <RESULT eventid="1196" points="431" swimtime="00:01:08.30" resultid="1690" heatid="2382" lane="2" entrytime="00:01:07.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Emili Gomes Xavier" birthdate="2010-09-08" gender="F" nation="BRA" license="372519" swrid="5717260" athleteid="1448" externalid="372519">
              <RESULTS>
                <RESULT eventid="1204" points="437" swimtime="00:01:24.49" resultid="1449" heatid="2387" lane="8" entrytime="00:01:25.51" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thais" lastname="Mariany Bortolazzi" birthdate="2006-05-02" gender="F" nation="BRA" license="357048" swrid="5600210" athleteid="1660" externalid="357048">
              <RESULTS>
                <RESULT eventid="1092" points="590" swimtime="00:09:37.82" resultid="1661" heatid="2337" lane="4" entrytime="00:09:27.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.02" />
                    <SPLIT distance="200" swimtime="00:02:21.55" />
                    <SPLIT distance="300" swimtime="00:03:34.14" />
                    <SPLIT distance="400" swimtime="00:04:47.33" />
                    <SPLIT distance="500" swimtime="00:05:59.92" />
                    <SPLIT distance="600" swimtime="00:07:12.81" />
                    <SPLIT distance="700" swimtime="00:08:25.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="556" swimtime="00:02:17.19" resultid="1662" heatid="2364" lane="5" entrytime="00:02:16.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helen" lastname="Barato Bernardi" birthdate="2006-07-27" gender="F" nation="BRA" license="317031" swrid="5717244" athleteid="1707" externalid="317031">
              <RESULTS>
                <RESULT eventid="1076" points="573" swimtime="00:02:45.54" resultid="1708" heatid="2331" lane="5" entrytime="00:02:41.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="467" swimtime="00:02:25.43" resultid="1709" heatid="2360" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="590" swimtime="00:01:16.42" resultid="1710" heatid="2388" lane="4" entrytime="00:01:13.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Yolanda Ferreira" birthdate="2008-03-17" gender="F" nation="BRA" license="358335" swrid="5600276" athleteid="1657" externalid="358335">
              <RESULTS>
                <RESULT eventid="1060" points="483" swimtime="00:01:05.89" resultid="1658" heatid="2318" lane="6" entrytime="00:01:04.27" entrycourse="LCM" />
                <RESULT eventid="1204" points="503" swimtime="00:01:20.63" resultid="1659" heatid="2388" lane="7" entrytime="00:01:19.51" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Clara Fernandes Pereira" birthdate="2009-11-19" gender="F" nation="BRA" license="344340" swrid="5600137" athleteid="1450" externalid="344340">
              <RESULTS>
                <RESULT eventid="1124" points="350" swimtime="00:01:18.67" resultid="1451" heatid="2347" lane="1" />
                <RESULT eventid="1092" points="523" swimtime="00:10:01.63" resultid="1452" heatid="2337" lane="3" entrytime="00:09:48.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.87" />
                    <SPLIT distance="200" swimtime="00:02:27.54" />
                    <SPLIT distance="300" swimtime="00:03:44.42" />
                    <SPLIT distance="400" swimtime="00:05:00.60" />
                    <SPLIT distance="500" swimtime="00:06:16.70" />
                    <SPLIT distance="600" swimtime="00:07:31.92" />
                    <SPLIT distance="700" swimtime="00:08:47.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="546" swimtime="00:02:18.07" resultid="1453" heatid="2364" lane="3" entrytime="00:02:17.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rene" lastname="Osternack Erbe" birthdate="2011-04-03" gender="M" nation="BRA" license="366907" swrid="5588842" athleteid="1623" externalid="366907">
              <RESULTS>
                <RESULT eventid="1116" points="325" swimtime="00:02:42.63" resultid="1624" heatid="2344" lane="7" entrytime="00:02:46.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="320" swimtime="00:02:29.02" resultid="1625" heatid="2367" lane="7" entrytime="00:02:29.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="305" swimtime="00:01:16.64" resultid="1626" heatid="2381" lane="8" entrytime="00:01:16.32" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietra" lastname="Ruschel Carvalho" birthdate="2009-03-21" gender="F" nation="BRA" license="324999" swrid="5600250" athleteid="1454" externalid="324999">
              <RESULTS>
                <RESULT eventid="1188" points="451" swimtime="00:01:14.72" resultid="1455" heatid="2378" lane="2" entrytime="00:01:16.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Muxfeldt" birthdate="2011-05-13" gender="F" nation="BRA" license="366903" swrid="5602563" athleteid="1611" externalid="366903">
              <RESULTS>
                <RESULT eventid="1060" points="427" swimtime="00:01:08.64" resultid="1612" heatid="2317" lane="8" entrytime="00:01:07.77" entrycourse="LCM" />
                <RESULT eventid="1092" points="388" swimtime="00:11:04.67" resultid="1613" heatid="2335" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.71" />
                    <SPLIT distance="200" swimtime="00:02:40.17" />
                    <SPLIT distance="300" swimtime="00:04:05.12" />
                    <SPLIT distance="400" swimtime="00:05:30.45" />
                    <SPLIT distance="500" swimtime="00:06:55.70" />
                    <SPLIT distance="600" swimtime="00:08:20.52" />
                    <SPLIT distance="700" swimtime="00:09:44.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="433" swimtime="00:02:29.09" resultid="1614" heatid="2363" lane="3" entrytime="00:02:26.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Godino" birthdate="2010-04-27" gender="F" nation="BRA" license="356355" swrid="5600176" athleteid="1561" externalid="356355">
              <RESULTS>
                <RESULT eventid="1060" points="374" swimtime="00:01:11.74" resultid="1562" heatid="2316" lane="1" entrytime="00:01:09.21" entrycourse="LCM" />
                <RESULT eventid="1092" points="383" swimtime="00:11:07.32" resultid="1563" heatid="2337" lane="2" entrytime="00:10:36.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.43" />
                    <SPLIT distance="200" swimtime="00:02:43.71" />
                    <SPLIT distance="300" swimtime="00:04:07.85" />
                    <SPLIT distance="400" swimtime="00:05:32.85" />
                    <SPLIT distance="500" swimtime="00:06:57.63" />
                    <SPLIT distance="600" swimtime="00:08:21.44" />
                    <SPLIT distance="700" swimtime="00:09:44.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="422" swimtime="00:02:30.45" resultid="1564" heatid="2363" lane="6" entrytime="00:02:27.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Martynychen" birthdate="2011-12-19" gender="M" nation="BRA" license="366893" swrid="5602557" athleteid="1592" externalid="366893">
              <RESULTS>
                <RESULT eventid="1116" status="DNS" swimtime="00:00:00.00" resultid="1593" heatid="2344" lane="2" entrytime="00:02:45.19" entrycourse="LCM" />
                <RESULT eventid="1100" points="364" swimtime="00:10:32.92" resultid="1594" heatid="2340" lane="5" entrytime="00:10:02.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.58" />
                    <SPLIT distance="200" swimtime="00:02:30.23" />
                    <SPLIT distance="300" swimtime="00:03:50.87" />
                    <SPLIT distance="400" swimtime="00:05:11.05" />
                    <SPLIT distance="500" swimtime="00:06:33.01" />
                    <SPLIT distance="600" swimtime="00:07:54.60" />
                    <SPLIT distance="700" swimtime="00:09:17.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="322" swimtime="00:02:28.80" resultid="1595" heatid="2367" lane="4" entrytime="00:02:22.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Vieira Motta" birthdate="2009-09-19" gender="M" nation="BRA" license="339064" swrid="5600271" athleteid="1523" externalid="339064">
              <RESULTS>
                <RESULT eventid="1100" points="486" swimtime="00:09:34.92" resultid="1524" heatid="2340" lane="4" entrytime="00:09:25.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.94" />
                    <SPLIT distance="200" swimtime="00:02:15.21" />
                    <SPLIT distance="300" swimtime="00:03:26.79" />
                    <SPLIT distance="400" swimtime="00:04:38.61" />
                    <SPLIT distance="500" swimtime="00:05:52.96" />
                    <SPLIT distance="600" swimtime="00:07:07.94" />
                    <SPLIT distance="700" swimtime="00:08:22.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="459" swimtime="00:01:06.87" resultid="1525" heatid="2383" lane="8" entrytime="00:01:05.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Valduga Artigas" birthdate="2009-06-01" gender="M" nation="BRA" license="339569" swrid="5600268" athleteid="1520" externalid="339569">
              <RESULTS>
                <RESULT comment="SW 8.3 - Movimento alternado das pernas ou pés.  (Tempo: 12:16)" eventid="1132" status="DSQ" swimtime="00:01:17.98" resultid="1521" heatid="2352" lane="8" entrytime="00:01:15.33" entrycourse="LCM" />
                <RESULT eventid="1068" points="323" swimtime="00:01:08.26" resultid="1522" heatid="2322" lane="8" entrytime="00:01:05.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Estevao" lastname="Valduga Artigas" birthdate="2009-06-01" gender="M" nation="BRA" license="339556" swrid="5600267" athleteid="1501" externalid="339556">
              <RESULTS>
                <RESULT eventid="1100" points="387" swimtime="00:10:19.89" resultid="1502" heatid="2339" lane="3" entrytime="00:10:47.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.86" />
                    <SPLIT distance="200" swimtime="00:02:28.81" />
                    <SPLIT distance="300" swimtime="00:03:47.69" />
                    <SPLIT distance="400" swimtime="00:05:07.14" />
                    <SPLIT distance="500" swimtime="00:06:26.24" />
                    <SPLIT distance="600" swimtime="00:07:45.26" />
                    <SPLIT distance="700" swimtime="00:09:04.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="309" swimtime="00:01:16.31" resultid="1503" heatid="2380" lane="3" entrytime="00:01:18.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Pereira Galle" birthdate="2011-08-02" gender="F" nation="BRA" license="369465" swrid="5627330" athleteid="1697" externalid="369465">
              <RESULTS>
                <RESULT eventid="1060" points="463" swimtime="00:01:06.84" resultid="1698" heatid="2312" lane="6" />
                <RESULT eventid="1156" points="444" swimtime="00:02:27.84" resultid="1699" heatid="2363" lane="7" entrytime="00:02:27.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="423" swimtime="00:01:25.38" resultid="1700" heatid="2387" lane="1" entrytime="00:01:24.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Magalhaes Dos Reis" birthdate="2010-05-05" gender="M" nation="BRA" license="356361" swrid="5600207" athleteid="1565" externalid="356361">
              <RESULTS>
                <RESULT eventid="1132" points="242" swimtime="00:01:19.31" resultid="1566" heatid="2351" lane="4" entrytime="00:01:16.51" entrycourse="LCM" />
                <RESULT eventid="1068" points="461" swimtime="00:01:00.65" resultid="1567" heatid="2325" lane="2" entrytime="00:00:59.61" entrycourse="LCM" />
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="1568" heatid="2391" lane="4" entrytime="00:01:20.10" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Mattioli" birthdate="2011-10-22" gender="F" nation="BRA" license="366896" swrid="5602559" athleteid="1596" externalid="366896">
              <RESULTS>
                <RESULT eventid="1092" points="445" swimtime="00:10:34.90" resultid="1597" heatid="2336" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.47" />
                    <SPLIT distance="200" swimtime="00:02:37.08" />
                    <SPLIT distance="300" swimtime="00:03:58.43" />
                    <SPLIT distance="400" swimtime="00:05:19.34" />
                    <SPLIT distance="500" swimtime="00:06:40.31" />
                    <SPLIT distance="600" swimtime="00:08:00.84" />
                    <SPLIT distance="700" swimtime="00:09:20.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1076" points="478" swimtime="00:02:55.89" resultid="1598" heatid="2331" lane="2" entrytime="00:02:58.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="David Cella" birthdate="2008-02-17" gender="M" nation="BRA" license="341107" swrid="5634581" athleteid="1701" externalid="341107">
              <RESULTS>
                <RESULT eventid="1068" points="639" swimtime="00:00:54.38" resultid="1702" heatid="2328" lane="6" entrytime="00:00:53.76" entrycourse="LCM" />
                <RESULT eventid="1196" points="529" swimtime="00:01:03.80" resultid="1703" heatid="2383" lane="1" entrytime="00:01:04.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelo" lastname="Vanhazebrouck" birthdate="2010-01-09" gender="M" nation="BRA" license="339043" swrid="5600269" athleteid="1533" externalid="339043">
              <RESULTS>
                <RESULT eventid="1132" points="307" swimtime="00:01:13.30" resultid="1534" heatid="2352" lane="5" entrytime="00:01:11.90" entrycourse="LCM" />
                <RESULT eventid="1068" points="431" swimtime="00:01:02.03" resultid="1535" heatid="2324" lane="4" entrytime="00:01:00.30" entrycourse="LCM" />
                <RESULT eventid="1164" points="397" swimtime="00:02:18.70" resultid="1536" heatid="2369" lane="6" entrytime="00:02:15.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Lacerda" birthdate="2011-05-09" gender="M" nation="BRA" license="366909" swrid="5602550" athleteid="1632" externalid="366909">
              <RESULTS>
                <RESULT eventid="1068" points="360" swimtime="00:01:05.86" resultid="1633" heatid="2321" lane="2" entrytime="00:01:06.86" entrycourse="LCM" />
                <RESULT eventid="1164" points="311" swimtime="00:02:30.46" resultid="1634" heatid="2367" lane="5" entrytime="00:02:24.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="358" swimtime="00:05:41.21" resultid="1635" heatid="2358" lane="6" entrytime="00:05:45.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.80" />
                    <SPLIT distance="200" swimtime="00:02:50.18" />
                    <SPLIT distance="300" swimtime="00:04:26.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Braun Prado" birthdate="2008-04-07" gender="M" nation="BRA" license="307663" swrid="5484324" athleteid="1526" externalid="307663">
              <RESULTS>
                <RESULT eventid="1116" points="512" swimtime="00:02:19.89" resultid="1527" heatid="2345" lane="5" entrytime="00:02:16.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="540" swimtime="00:00:57.52" resultid="1528" heatid="2327" lane="8" entrytime="00:00:57.65" entrycourse="LCM" />
                <RESULT eventid="1196" points="557" swimtime="00:01:02.69" resultid="1529" heatid="2383" lane="7" entrytime="00:01:02.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucca" lastname="Cruz Tonin" birthdate="2004-03-19" gender="M" nation="BRA" license="270821" swrid="5622272" athleteid="1636" externalid="270821">
              <RESULTS>
                <RESULT eventid="1116" points="698" swimtime="00:02:06.15" resultid="1637" heatid="2345" lane="4" entrytime="00:02:02.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="742" swimtime="00:00:56.98" resultid="1638" heatid="2383" lane="4" entrytime="00:00:56.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pablo" lastname="Souza Tavares" birthdate="2006-05-03" gender="M" nation="BRA" license="331982" swrid="5600261" athleteid="1456" externalid="331982">
              <RESULTS>
                <RESULT eventid="1132" points="681" swimtime="00:00:56.19" resultid="1457" heatid="2355" lane="3" entrytime="00:00:57.06" entrycourse="LCM" />
                <RESULT eventid="1068" points="732" swimtime="00:00:51.98" resultid="1458" heatid="2328" lane="4" entrytime="00:00:52.43" entrycourse="LCM" />
                <RESULT eventid="1196" points="639" swimtime="00:00:59.90" resultid="1459" heatid="2383" lane="5" entrytime="00:00:59.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joshua" lastname="Gomide Capraro" birthdate="2009-01-18" gender="M" nation="BRA" license="339030" swrid="5600177" athleteid="1460" externalid="339030">
              <RESULTS>
                <RESULT eventid="1164" points="518" swimtime="00:02:06.95" resultid="1461" heatid="2371" lane="6" entrytime="00:02:02.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Fontolan Gomes" birthdate="2010-07-02" gender="M" nation="BRA" license="356245" swrid="5588705" athleteid="1537" externalid="356245">
              <RESULTS>
                <RESULT eventid="1116" points="404" swimtime="00:02:31.30" resultid="1538" heatid="2344" lane="4" entrytime="00:02:34.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="382" swimtime="00:02:20.57" resultid="1539" heatid="2368" lane="5" entrytime="00:02:20.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="396" swimtime="00:01:10.24" resultid="1540" heatid="2381" lane="3" entrytime="00:01:11.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Sachser Rocha" birthdate="2008-07-09" gender="M" nation="BRA" license="330072" swrid="5600254" athleteid="1496" externalid="330072">
              <RESULTS>
                <RESULT eventid="1132" points="581" swimtime="00:00:59.26" resultid="1497" heatid="2355" lane="2" entrytime="00:00:58.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Iglesias Vargas" birthdate="2009-01-11" gender="M" nation="BRA" license="324792" swrid="5600189" athleteid="1477" externalid="324792">
              <RESULTS>
                <RESULT eventid="1068" points="558" swimtime="00:00:56.91" resultid="1478" heatid="2327" lane="3" entrytime="00:00:56.42" entrycourse="LCM" />
                <RESULT eventid="1164" points="557" swimtime="00:02:03.95" resultid="1479" heatid="2371" lane="3" entrytime="00:02:01.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="414" swimtime="00:01:09.23" resultid="1480" heatid="2379" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Galvao" birthdate="2011-03-11" gender="M" nation="BRA" license="381989" swrid="5602541" athleteid="1673" externalid="381989">
              <RESULTS>
                <RESULT eventid="1132" points="169" swimtime="00:01:29.42" resultid="1674" heatid="2350" lane="5" />
                <RESULT eventid="1068" points="353" swimtime="00:01:06.27" resultid="1675" heatid="2321" lane="3" entrytime="00:01:06.21" entrycourse="LCM" />
                <RESULT eventid="1164" points="314" swimtime="00:02:30.00" resultid="1676" heatid="2367" lane="2" entrytime="00:02:27.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo" lastname="De Lima Cavalcanti" birthdate="2009-12-17" gender="M" nation="BRA" license="380965" swrid="5634589" athleteid="1704" externalid="380965">
              <RESULTS>
                <RESULT eventid="1132" points="534" swimtime="00:01:00.93" resultid="1705" heatid="2355" lane="7" entrytime="00:00:59.99" entrycourse="LCM" />
                <RESULT eventid="1196" points="418" swimtime="00:01:09.00" resultid="1706" heatid="2379" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="De Albuquerque" birthdate="2010-06-08" gender="F" nation="BRA" license="356249" swrid="5600145" athleteid="1541" externalid="356249">
              <RESULTS>
                <RESULT eventid="1060" points="387" swimtime="00:01:10.90" resultid="1542" heatid="2315" lane="5" entrytime="00:01:10.44" entrycourse="LCM" />
                <RESULT eventid="1108" points="407" swimtime="00:02:46.05" resultid="1543" heatid="2342" lane="6" entrytime="00:02:44.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="310" swimtime="00:01:34.69" resultid="1544" heatid="2385" lane="6" entrytime="00:01:36.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Bussmann" birthdate="2007-01-16" gender="F" nation="BRA" license="313781" swrid="5579983" athleteid="1462" externalid="313781">
              <RESULTS>
                <RESULT eventid="1076" points="484" swimtime="00:02:55.19" resultid="1463" heatid="2331" lane="4" entrytime="00:02:37.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="475" swimtime="00:05:40.60" resultid="1464" heatid="2356" lane="5" />
                <RESULT eventid="1204" points="580" swimtime="00:01:16.87" resultid="1465" heatid="2388" lane="5" entrytime="00:01:14.82" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Ramos Marcon" birthdate="2008-01-12" gender="M" nation="BRA" license="372281" swrid="5600240" athleteid="1677" externalid="372281">
              <RESULTS>
                <RESULT eventid="1068" points="573" swimtime="00:00:56.41" resultid="1678" heatid="2327" lane="4" entrytime="00:00:55.73" entrycourse="LCM" />
                <RESULT eventid="1164" points="515" swimtime="00:02:07.22" resultid="1679" heatid="2371" lane="1" entrytime="00:02:07.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolau" lastname="Neto" birthdate="2011-03-22" gender="M" nation="BRA" license="366906" swrid="5602565" athleteid="1619" externalid="366906">
              <RESULTS>
                <RESULT eventid="1068" points="445" swimtime="00:01:01.34" resultid="1620" heatid="2324" lane="5" entrytime="00:01:01.13" entrycourse="LCM" />
                <RESULT eventid="1164" points="394" swimtime="00:02:19.11" resultid="1621" heatid="2368" lane="2" entrytime="00:02:20.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="342" swimtime="00:01:21.29" resultid="1622" heatid="2392" lane="8" entrytime="00:01:19.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Fontoura" birthdate="2010-08-26" gender="M" nation="BRA" license="338922" swrid="5600167" athleteid="1569" externalid="338922">
              <RESULTS>
                <RESULT eventid="1132" points="284" swimtime="00:01:15.22" resultid="1570" heatid="2352" lane="7" entrytime="00:01:14.26" entrycourse="LCM" />
                <RESULT eventid="1068" points="395" swimtime="00:01:03.82" resultid="1571" heatid="2323" lane="2" entrytime="00:01:03.31" entrycourse="LCM" />
                <RESULT eventid="1164" points="361" swimtime="00:02:23.25" resultid="1572" heatid="2368" lane="8" entrytime="00:02:21.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Martinez Diniz" birthdate="2008-11-22" gender="M" nation="BRA" license="339400" swrid="5717283" athleteid="1498" externalid="339400">
              <RESULTS>
                <RESULT eventid="1068" points="553" swimtime="00:00:57.07" resultid="1499" heatid="2327" lane="6" entrytime="00:00:56.70" entrycourse="LCM" />
                <RESULT eventid="1164" points="478" swimtime="00:02:10.44" resultid="1500" heatid="2370" lane="5" entrytime="00:02:10.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Guimaraes E Souza" birthdate="2008-12-21" gender="M" nation="BRA" license="376972" swrid="5600182" athleteid="1663" externalid="376972">
              <RESULTS>
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Tempo: 10:15), Na volta dos 50m e 150m." eventid="1084" status="DSQ" swimtime="00:02:41.61" resultid="1664" heatid="2334" lane="3" entrytime="00:02:39.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="543" swimtime="00:01:09.71" resultid="1665" heatid="2393" lane="6" entrytime="00:01:09.22" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Brandt De Macedo" birthdate="2010-01-13" gender="M" nation="BRA" license="338925" swrid="5588565" athleteid="1573" externalid="338925">
              <RESULTS>
                <RESULT eventid="1132" points="309" swimtime="00:01:13.13" resultid="1574" heatid="2352" lane="1" entrytime="00:01:14.58" entrycourse="LCM" />
                <RESULT eventid="1068" points="461" swimtime="00:01:00.63" resultid="1575" heatid="2325" lane="7" entrytime="00:00:59.79" entrycourse="LCM" />
                <RESULT eventid="1164" points="439" swimtime="00:02:14.12" resultid="1576" heatid="2370" lane="8" entrytime="00:02:12.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Sabedotti" birthdate="2002-07-07" gender="M" nation="BRA" license="134704" swrid="5600252" athleteid="1530" externalid="134704">
              <RESULTS>
                <RESULT eventid="1132" points="660" swimtime="00:00:56.79" resultid="1531" heatid="2355" lane="4" entrytime="00:00:55.31" entrycourse="LCM" />
                <RESULT eventid="1212" points="607" swimtime="00:01:07.17" resultid="1532" heatid="2393" lane="4" entrytime="00:01:04.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Cabrera Cirino" birthdate="2011-01-28" gender="M" nation="BRA" license="369531" swrid="5588569" athleteid="1644" externalid="369531">
              <RESULTS>
                <RESULT eventid="1100" points="457" swimtime="00:09:46.72" resultid="1645" heatid="2338" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.68" />
                    <SPLIT distance="200" swimtime="00:02:24.58" />
                    <SPLIT distance="300" swimtime="00:03:38.70" />
                    <SPLIT distance="400" swimtime="00:04:52.90" />
                    <SPLIT distance="500" swimtime="00:06:07.31" />
                    <SPLIT distance="600" swimtime="00:07:21.57" />
                    <SPLIT distance="700" swimtime="00:08:35.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="473" swimtime="00:01:00.12" resultid="1646" heatid="2326" lane="8" entrytime="00:00:58.96" entrycourse="LCM" />
                <RESULT eventid="1164" points="461" swimtime="00:02:12.03" resultid="1647" heatid="2369" lane="4" entrytime="00:02:12.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="394" swimtime="00:01:10.35" resultid="1648" heatid="2382" lane="8" entrytime="00:01:08.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo" lastname="Gabriel Nascimento" birthdate="2008-11-14" gender="M" nation="BRA" license="348028" swrid="5600171" athleteid="1691" externalid="348028">
              <RESULTS>
                <RESULT eventid="1132" points="465" swimtime="00:01:03.81" resultid="1692" heatid="2354" lane="2" entrytime="00:01:03.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Fontana" birthdate="2011-12-29" gender="M" nation="BRA" license="366897" swrid="5602539" athleteid="1599" externalid="366897">
              <RESULTS>
                <RESULT eventid="1068" points="232" swimtime="00:01:16.17" resultid="1600" heatid="2320" lane="1" entrytime="00:01:17.96" entrycourse="LCM" />
                <RESULT eventid="1164" status="DNS" swimtime="00:00:00.00" resultid="1601" heatid="2365" lane="4" entrytime="00:02:57.40" entrycourse="LCM" />
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="1602" heatid="2390" lane="1" entrytime="00:01:34.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Gustavo Souza" birthdate="2011-08-24" gender="M" nation="BRA" license="366901" swrid="5588733" athleteid="1607" externalid="366901">
              <RESULTS>
                <RESULT eventid="1132" points="330" swimtime="00:01:11.51" resultid="1608" heatid="2352" lane="4" entrytime="00:01:11.45" entrycourse="LCM" />
                <RESULT eventid="1148" points="322" swimtime="00:05:53.70" resultid="1609" heatid="2358" lane="2" entrytime="00:05:46.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.32" />
                    <SPLIT distance="200" swimtime="00:02:49.21" />
                    <SPLIT distance="300" swimtime="00:04:36.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="247" swimtime="00:02:55.68" resultid="1610" heatid="2374" lane="7" entrytime="00:02:43.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nina" lastname="Rocha Ribeiro Da Silva" birthdate="2010-09-22" gender="F" nation="BRA" license="367216" swrid="5588884" athleteid="1680" externalid="367216">
              <RESULTS>
                <RESULT eventid="1060" points="448" swimtime="00:01:07.55" resultid="1681" heatid="2316" lane="2" entrytime="00:01:09.05" entrycourse="LCM" />
                <RESULT eventid="1156" points="429" swimtime="00:02:29.59" resultid="1682" heatid="2362" lane="7" entrytime="00:02:32.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="464" swimtime="00:01:22.82" resultid="1683" heatid="2388" lane="1" entrytime="00:01:20.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Heloisa Souza" birthdate="2007-01-15" gender="F" nation="BRA" license="336615" swrid="5600184" athleteid="1481" externalid="336615">
              <RESULTS>
                <RESULT eventid="1060" points="560" swimtime="00:01:02.70" resultid="1482" heatid="2318" lane="4" entrytime="00:00:59.80" entrycourse="LCM" />
                <RESULT eventid="1092" points="552" swimtime="00:09:50.78" resultid="1483" heatid="2337" lane="5" entrytime="00:09:41.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.72" />
                    <SPLIT distance="200" swimtime="00:02:23.09" />
                    <SPLIT distance="300" swimtime="00:03:37.95" />
                    <SPLIT distance="400" swimtime="00:04:53.24" />
                    <SPLIT distance="500" swimtime="00:06:07.64" />
                    <SPLIT distance="600" swimtime="00:07:21.93" />
                    <SPLIT distance="700" swimtime="00:08:36.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="591" swimtime="00:02:14.40" resultid="1484" heatid="2364" lane="4" entrytime="00:02:08.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Prosdocimo" birthdate="2010-11-23" gender="F" nation="BRA" license="356251" swrid="5600238" athleteid="1545" externalid="356251">
              <RESULTS>
                <RESULT eventid="1060" points="475" swimtime="00:01:06.24" resultid="1546" heatid="2318" lane="1" entrytime="00:01:05.28" entrycourse="LCM" />
                <RESULT eventid="1108" points="394" swimtime="00:02:47.88" resultid="1547" heatid="2342" lane="2" entrytime="00:02:47.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="431" swimtime="00:01:15.86" resultid="1548" heatid="2378" lane="3" entrytime="00:01:15.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Francisco Saldo" birthdate="2007-01-23" gender="M" nation="BRA" license="313537" swrid="5600169" athleteid="1466" externalid="313537">
              <RESULTS>
                <RESULT eventid="1132" points="596" swimtime="00:00:58.75" resultid="1467" heatid="2355" lane="5" entrytime="00:00:56.64" entrycourse="LCM" />
                <RESULT eventid="1196" status="DNS" swimtime="00:00:00.00" resultid="1468" heatid="2380" lane="8" />
                <RESULT eventid="1180" points="640" swimtime="00:02:07.98" resultid="1469" heatid="2374" lane="4" entrytime="00:02:02.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Trevisan" birthdate="2000-11-28" gender="M" nation="BRA" license="346847" swrid="5600266" athleteid="1684" externalid="346847">
              <RESULTS>
                <RESULT eventid="1068" points="604" swimtime="00:00:55.41" resultid="1685" heatid="2328" lane="7" entrytime="00:00:54.62" entrycourse="LCM" />
                <RESULT eventid="1164" points="527" swimtime="00:02:06.24" resultid="1686" heatid="2371" lane="2" entrytime="00:02:03.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2864" nation="BRA" region="PR" clubid="1220" swrid="93756" name="Associacao De Pais E Amigos Da Natacao De Ponta Gr" shortname="Apan Ponta Grossa">
          <ATHLETES>
            <ATHLETE firstname="Rafael" lastname="Gueiber Montes" birthdate="2009-03-09" gender="M" nation="BRA" license="342154" swrid="5600179" athleteid="1221" externalid="342154">
              <RESULTS>
                <RESULT eventid="1132" points="481" swimtime="00:01:03.08" resultid="1222" heatid="2349" lane="4" />
                <RESULT eventid="1068" points="652" swimtime="00:00:54.02" resultid="1223" heatid="2328" lane="2" entrytime="00:00:54.10" entrycourse="LCM" />
                <RESULT eventid="1164" points="582" swimtime="00:02:02.10" resultid="1224" heatid="2371" lane="5" entrytime="00:02:00.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="472" swimtime="00:01:06.26" resultid="1225" heatid="2383" lane="2" entrytime="00:01:01.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Allana" lastname="Lacerda" birthdate="2005-03-15" gender="F" nation="BRA" license="295186" swrid="5600197" athleteid="1232" externalid="295186">
              <RESULTS>
                <RESULT eventid="1076" points="427" swimtime="00:03:02.55" resultid="1233" heatid="2331" lane="8" entrytime="00:02:59.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="391" swimtime="00:01:27.67" resultid="1234" heatid="2387" lane="3" entrytime="00:01:22.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Delinski" birthdate="2009-11-28" gender="F" nation="BRA" license="385190" swrid="5600150" athleteid="1238" externalid="385190">
              <RESULTS>
                <RESULT eventid="1076" points="321" swimtime="00:03:20.78" resultid="1239" heatid="2330" lane="1" entrytime="00:03:21.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="399" swimtime="00:01:27.06" resultid="1240" heatid="2386" lane="5" entrytime="00:01:27.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Franca Berger" birthdate="2010-05-07" gender="F" nation="BRA" license="399692" swrid="5653290" athleteid="1251" externalid="399692">
              <RESULTS>
                <RESULT eventid="1060" points="293" swimtime="00:01:17.77" resultid="1252" heatid="2313" lane="5" entrytime="00:01:17.55" entrycourse="LCM" />
                <RESULT eventid="1204" points="222" swimtime="00:01:45.84" resultid="1253" heatid="2385" lane="8" entrytime="00:01:44.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Brenda" lastname="Gabriele Carvalho" birthdate="2010-04-11" gender="F" nation="BRA" license="399557" swrid="5658060" athleteid="1244" externalid="399557">
              <RESULTS>
                <RESULT eventid="1060" points="271" swimtime="00:01:19.90" resultid="1245" heatid="2314" lane="1" entrytime="00:01:16.26" entrycourse="LCM" />
                <RESULT eventid="1204" points="255" swimtime="00:01:41.04" resultid="1246" heatid="2385" lane="7" entrytime="00:01:43.10" entrycourse="LCM" />
                <RESULT eventid="1188" points="255" swimtime="00:01:30.30" resultid="1247" heatid="2377" lane="8" entrytime="00:01:28.44" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Augusto" lastname="Tramontin" birthdate="2011-11-29" gender="M" nation="BRA" license="399691" swrid="5652901" athleteid="1248" externalid="399691">
              <RESULTS>
                <RESULT eventid="1068" points="422" swimtime="00:01:02.43" resultid="1249" heatid="2322" lane="3" entrytime="00:01:04.15" entrycourse="LCM" />
                <RESULT eventid="1212" points="338" swimtime="00:01:21.62" resultid="1250" heatid="2391" lane="5" entrytime="00:01:23.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Pontes Mattioli" birthdate="2011-09-10" gender="F" nation="BRA" license="366914" swrid="5602572" athleteid="1254" externalid="366914">
              <RESULTS>
                <RESULT eventid="1060" points="427" swimtime="00:01:08.63" resultid="1255" heatid="2315" lane="8" entrytime="00:01:11.67" entrycourse="LCM" />
                <RESULT eventid="1108" points="351" swimtime="00:02:54.51" resultid="1256" heatid="2341" lane="4" entrytime="00:03:01.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="341" swimtime="00:01:22.03" resultid="1257" heatid="2377" lane="3" entrytime="00:01:23.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Campagnoli" birthdate="2009-04-13" gender="F" nation="BRA" license="366915" swrid="5600128" athleteid="1235" externalid="366915">
              <RESULTS>
                <RESULT eventid="1108" points="492" swimtime="00:02:35.96" resultid="1236" heatid="2342" lane="5" entrytime="00:02:36.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="457" swimtime="00:01:14.42" resultid="1237" heatid="2378" lane="5" entrytime="00:01:11.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fegert" birthdate="2009-04-13" gender="M" nation="BRA" license="353813" swrid="5622279" athleteid="1241" externalid="353813">
              <RESULTS>
                <RESULT eventid="1132" points="453" swimtime="00:01:04.36" resultid="1242" heatid="2354" lane="8" entrytime="00:01:05.20" entrycourse="LCM" />
                <RESULT eventid="1164" points="458" swimtime="00:02:12.30" resultid="1243" heatid="2365" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Chi Kravchychyn" birthdate="2009-09-27" gender="M" nation="BRA" license="344268" swrid="5600134" athleteid="1226" externalid="344268">
              <RESULTS>
                <RESULT eventid="1132" points="512" swimtime="00:01:01.78" resultid="1227" heatid="2354" lane="5" entrytime="00:01:01.32" entrycourse="LCM" />
                <RESULT eventid="1084" points="540" swimtime="00:02:34.06" resultid="1228" heatid="2334" lane="5" entrytime="00:02:30.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="488" swimtime="00:05:07.95" resultid="1229" heatid="2358" lane="4" entrytime="00:04:51.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.99" />
                    <SPLIT distance="200" swimtime="00:02:29.85" />
                    <SPLIT distance="300" swimtime="00:03:54.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="512" swimtime="00:01:11.09" resultid="1230" heatid="2393" lane="3" entrytime="00:01:09.09" entrycourse="LCM" />
                <RESULT eventid="1180" points="383" swimtime="00:02:31.84" resultid="1231" heatid="2374" lane="3" entrytime="00:02:16.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Xavier Teixeira" birthdate="2011-09-22" gender="M" nation="BRA" license="415193" athleteid="1260" externalid="415193">
              <RESULTS>
                <RESULT eventid="1068" points="269" swimtime="00:01:12.53" resultid="1261" heatid="2319" lane="5" />
                <RESULT eventid="1196" points="185" swimtime="00:01:30.53" resultid="1262" heatid="2379" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Lievore" birthdate="2010-06-07" gender="F" nation="BRA" license="414856" swrid="5757092" athleteid="1258" externalid="414856">
              <RESULTS>
                <RESULT eventid="1060" points="333" swimtime="00:01:14.59" resultid="1259" heatid="2314" lane="6" entrytime="00:01:15.00" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
