<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.79462">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Londrina" name="12º Jogos Paradesportivos 2024" course="SCM" hostclub="Secretaria do Esporte do Governo do Estado do Paraná" hostclub.url="https://www.esporte.pr.gov.br/PARAJAPS" number="S2304" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/evento/natacao/S2304" startmethod="2" timing="AUTOMATIC" touchpad="ONESIDE" masters="F" state="PR" nation="BRA">
      <AGEDATE value="2024-05-30" type="YEAR" />
      <POOL name="Associação dos Funcionários Municipais de Londrina" lanemin="1" lanemax="6" />
      <FACILITY city="Londrina" name="Associação dos Funcionários Municipais de Londrina" nation="BRA" state="PR" street="Rua dos Funcionários, 363" street2="Nikko" zip="86047-080" />
      <POINTTABLE pointtableid="3016" name="FINA Point Scoring" version="2023" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-05-30" daytime="09:00" endtime="12:36" number="1" officialmeeting="08:30" teamleadermeeting="08:50" warmupfrom="08:00" warmupuntil="08:50">
          <EVENTS>
            <EVENT eventid="1060" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="-1" agemin="-1" name="Físico-Motora S1" handicap="1" />
                <AGEGROUP agegroupid="1122" agemax="-1" agemin="-1" name="Físico-Motora S2" handicap="2" />
                <AGEGROUP agegroupid="1123" agemax="-1" agemin="-1" name="Físico-Motora S3" handicap="3" />
                <AGEGROUP agegroupid="1124" agemax="-1" agemin="-1" name="Físico-Motora S4" handicap="4" />
                <AGEGROUP agegroupid="1125" agemax="-1" agemin="-1" name="Físico-Motora S5" handicap="5" />
                <AGEGROUP agegroupid="1126" agemax="-1" agemin="-1" name="Físico-Motora S6" handicap="6">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4092" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="-1" agemin="-1" name="Físico-Motora S7" handicap="7" />
                <AGEGROUP agegroupid="1128" agemax="-1" agemin="-1" name="Físico-Motora S8" handicap="8" />
                <AGEGROUP agegroupid="1129" agemax="-1" agemin="-1" name="Físico-Motora S9" handicap="9" />
                <AGEGROUP agegroupid="1130" agemax="-1" agemin="-1" name="Físico-Motora S10" handicap="10" />
                <AGEGROUP agegroupid="1131" agemax="-1" agemin="-1" name="Visual S11" handicap="11" />
                <AGEGROUP agegroupid="1132" agemax="-1" agemin="-1" name="Visual S12" handicap="12" />
                <AGEGROUP agegroupid="1133" agemax="-1" agemin="-1" name="Visual S13" handicap="13" />
                <AGEGROUP agegroupid="1134" agemax="-1" agemin="-1" name="Intelectual S14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3966" />
                    <RANKING order="2" place="2" resultid="4040" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="-1" agemin="-1" name="Intelectual S21 (SD)" handicap="21" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4213" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1766" />
                <TIMESTANDARDREF timestandardlistid="1774" />
                <TIMESTANDARDREF timestandardlistid="1780" />
                <TIMESTANDARDREF timestandardlistid="1786" />
                <TIMESTANDARDREF timestandardlistid="1792" />
                <TIMESTANDARDREF timestandardlistid="1798" />
                <TIMESTANDARDREF timestandardlistid="1804" />
                <TIMESTANDARDREF timestandardlistid="1810" />
                <TIMESTANDARDREF timestandardlistid="1816" />
                <TIMESTANDARDREF timestandardlistid="1822" />
                <TIMESTANDARDREF timestandardlistid="1828" />
                <TIMESTANDARDREF timestandardlistid="1834" />
                <TIMESTANDARDREF timestandardlistid="1840" />
                <TIMESTANDARDREF timestandardlistid="1846" />
                <TIMESTANDARDREF timestandardlistid="1852" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1062" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1644" agemax="-1" agemin="-1" name="Físico-Motora S1" handicap="1" />
                <AGEGROUP agegroupid="1645" agemax="-1" agemin="-1" name="Físico-Motora S2" handicap="2" />
                <AGEGROUP agegroupid="1646" agemax="-1" agemin="-1" name="Físico-Motora S3" handicap="3" />
                <AGEGROUP agegroupid="1647" agemax="-1" agemin="-1" name="Físico-Motora S4" handicap="4" />
                <AGEGROUP agegroupid="1648" agemax="-1" agemin="-1" name="Físico-Motora S5" handicap="5" />
                <AGEGROUP agegroupid="1649" agemax="-1" agemin="-1" name="Físico-Motora S6" handicap="6">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3934" />
                    <RANKING order="2" place="2" resultid="3994" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1650" agemax="-1" agemin="-1" name="Físico-Motora S7" handicap="7">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4027" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1651" agemax="-1" agemin="-1" name="Físico-Motora S8" handicap="8" />
                <AGEGROUP agegroupid="1652" agemax="-1" agemin="-1" name="Físico-Motora S9" handicap="9" />
                <AGEGROUP agegroupid="1653" agemax="-1" agemin="-1" name="Físico-Motora S10" handicap="10" />
                <AGEGROUP agegroupid="1654" agemax="-1" agemin="-1" name="Visual S11" handicap="11">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4075" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1655" agemax="-1" agemin="-1" name="Visual S12" handicap="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1656" agemax="-1" agemin="-1" name="Visual S13" handicap="13" />
                <AGEGROUP agegroupid="1657" agemax="-1" agemin="-1" name="Intelectual S14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3931" />
                    <RANKING order="2" place="2" resultid="3921" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1659" agemax="-1" agemin="-1" name="Intelectual S21 (SD)" handicap="21">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3978" />
                    <RANKING order="2" place="2" resultid="3962" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4214" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4215" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1764" />
                <TIMESTANDARDREF timestandardlistid="1772" />
                <TIMESTANDARDREF timestandardlistid="1778" />
                <TIMESTANDARDREF timestandardlistid="1784" />
                <TIMESTANDARDREF timestandardlistid="1790" />
                <TIMESTANDARDREF timestandardlistid="1796" />
                <TIMESTANDARDREF timestandardlistid="1802" />
                <TIMESTANDARDREF timestandardlistid="1808" />
                <TIMESTANDARDREF timestandardlistid="1814" />
                <TIMESTANDARDREF timestandardlistid="1820" />
                <TIMESTANDARDREF timestandardlistid="1826" />
                <TIMESTANDARDREF timestandardlistid="1832" />
                <TIMESTANDARDREF timestandardlistid="1838" />
                <TIMESTANDARDREF timestandardlistid="1844" />
                <TIMESTANDARDREF timestandardlistid="1850" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1064" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1628" agemax="-1" agemin="-1" name="Físico-Motora S1" handicap="1" />
                <AGEGROUP agegroupid="1629" agemax="-1" agemin="-1" name="Físico-Motora S2" handicap="2" />
                <AGEGROUP agegroupid="1630" agemax="-1" agemin="-1" name="Físico-Motora S3" handicap="3" />
                <AGEGROUP agegroupid="1631" agemax="-1" agemin="-1" name="Físico-Motora S4" handicap="4" />
                <AGEGROUP agegroupid="1632" agemax="-1" agemin="-1" name="Físico-Motora S5" handicap="5">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1633" agemax="-1" agemin="-1" name="Físico-Motora S6" handicap="6">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4059" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1634" agemax="-1" agemin="-1" name="Físico-Motora S7" handicap="7">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4036" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1635" agemax="-1" agemin="-1" name="Físico-Motora S8" handicap="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4153" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1636" agemax="-1" agemin="-1" name="Físico-Motora S9" handicap="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4009" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1637" agemax="-1" agemin="-1" name="Físico-Motora S10" handicap="10" />
                <AGEGROUP agegroupid="1638" agemax="-1" agemin="-1" name="Visual S11" handicap="11" />
                <AGEGROUP agegroupid="1639" agemax="-1" agemin="-1" name="Visual S12" handicap="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3946" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1640" agemax="-1" agemin="-1" name="Visual S13" handicap="13" />
                <AGEGROUP agegroupid="1641" agemax="-1" agemin="-1" name="Intelectual S14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3991" />
                    <RANKING order="2" place="2" resultid="3997" />
                    <RANKING order="3" place="-1" resultid="4041" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1642" agemax="-1" agemin="-1" name="Intelectual S18 (TEA)" handicap="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4099" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1643" agemax="-1" agemin="-1" name="Intelectual S21 (SD)" handicap="21">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4002" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4216" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4217" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1766" />
                <TIMESTANDARDREF timestandardlistid="1774" />
                <TIMESTANDARDREF timestandardlistid="1780" />
                <TIMESTANDARDREF timestandardlistid="1786" />
                <TIMESTANDARDREF timestandardlistid="1792" />
                <TIMESTANDARDREF timestandardlistid="1798" />
                <TIMESTANDARDREF timestandardlistid="1804" />
                <TIMESTANDARDREF timestandardlistid="1810" />
                <TIMESTANDARDREF timestandardlistid="1816" />
                <TIMESTANDARDREF timestandardlistid="1822" />
                <TIMESTANDARDREF timestandardlistid="1828" />
                <TIMESTANDARDREF timestandardlistid="1834" />
                <TIMESTANDARDREF timestandardlistid="1840" />
                <TIMESTANDARDREF timestandardlistid="1846" />
                <TIMESTANDARDREF timestandardlistid="1852" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1066" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1612" agemax="-1" agemin="-1" name="Físico-Motora S1" handicap="1" />
                <AGEGROUP agegroupid="1613" agemax="-1" agemin="-1" name="Físico-Motora S2" handicap="2" />
                <AGEGROUP agegroupid="1614" agemax="-1" agemin="-1" name="Físico-Motora S3" handicap="3" />
                <AGEGROUP agegroupid="1615" agemax="-1" agemin="-1" name="Físico-Motora S4" handicap="4">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1616" agemax="-1" agemin="-1" name="Físico-Motora S5" handicap="5">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3884" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1617" agemax="-1" agemin="-1" name="Físico-Motora S6" handicap="6">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3858" />
                    <RANKING order="2" place="2" resultid="3949" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1618" agemax="-1" agemin="-1" name="Físico-Motora S7" handicap="7">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1619" agemax="-1" agemin="-1" name="Físico-Motora S8" handicap="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4170" />
                    <RANKING order="2" place="2" resultid="4125" />
                    <RANKING order="3" place="3" resultid="3954" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1620" agemax="-1" agemin="-1" name="Físico-Motora S9" handicap="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3867" />
                    <RANKING order="2" place="-1" resultid="3925" />
                    <RANKING order="3" place="-1" resultid="3863" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1621" agemax="-1" agemin="-1" name="Físico-Motora S10" handicap="10" />
                <AGEGROUP agegroupid="1622" agemax="-1" agemin="-1" name="Visual S11" handicap="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1623" agemax="-1" agemin="-1" name="Visual S12" handicap="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3971" />
                    <RANKING order="2" place="-1" resultid="4005" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1624" agemax="-1" agemin="-1" name="Visual S13" handicap="13" />
                <AGEGROUP agegroupid="1625" agemax="-1" agemin="-1" name="Intelectual S14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4108" />
                    <RANKING order="2" place="2" resultid="3922" />
                    <RANKING order="3" place="-1" resultid="4050" />
                    <RANKING order="4" place="-1" resultid="4180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1626" agemax="-1" agemin="-1" name="Intelectual S18 (TEA)" handicap="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4080" />
                    <RANKING order="2" place="2" resultid="3974" />
                    <RANKING order="3" place="3" resultid="4014" />
                    <RANKING order="4" place="4" resultid="4095" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1627" agemax="-1" agemin="-1" name="Intelectual S21 (SD)" handicap="21">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4157" />
                    <RANKING order="2" place="2" resultid="4088" />
                    <RANKING order="3" place="3" resultid="3979" />
                    <RANKING order="4" place="4" resultid="3871" />
                    <RANKING order="5" place="5" resultid="4020" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4218" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4219" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4220" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4221" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4222" number="5" order="5" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1764" />
                <TIMESTANDARDREF timestandardlistid="1772" />
                <TIMESTANDARDREF timestandardlistid="1778" />
                <TIMESTANDARDREF timestandardlistid="1784" />
                <TIMESTANDARDREF timestandardlistid="1790" />
                <TIMESTANDARDREF timestandardlistid="1796" />
                <TIMESTANDARDREF timestandardlistid="1802" />
                <TIMESTANDARDREF timestandardlistid="1808" />
                <TIMESTANDARDREF timestandardlistid="1814" />
                <TIMESTANDARDREF timestandardlistid="1820" />
                <TIMESTANDARDREF timestandardlistid="1826" />
                <TIMESTANDARDREF timestandardlistid="1832" />
                <TIMESTANDARDREF timestandardlistid="1838" />
                <TIMESTANDARDREF timestandardlistid="1844" />
                <TIMESTANDARDREF timestandardlistid="1850" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1068" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1599" agemax="-1" agemin="-1" name="Físico-Motora SB4" handicap="4" />
                <AGEGROUP agegroupid="1600" agemax="-1" agemin="-1" name="Físico-Motora SB5" handicap="5">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1601" agemax="-1" agemin="-1" name="Físico-Motora SB6" handicap="6" />
                <AGEGROUP agegroupid="1602" agemax="-1" agemin="-1" name="Físico-Motora SB7" handicap="7" />
                <AGEGROUP agegroupid="1603" agemax="-1" agemin="-1" name="Físico-Motora SB8" handicap="8" />
                <AGEGROUP agegroupid="1604" agemax="-1" agemin="-1" name="Físico-Motora SB9" handicap="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1605" agemax="-1" agemin="-1" name="Físico-Motora SB10" handicap="10" />
                <AGEGROUP agegroupid="1606" agemax="-1" agemin="-1" name="Visual SB11" handicap="11" />
                <AGEGROUP agegroupid="1607" agemax="-1" agemin="-1" name="Visual SB12" handicap="12" />
                <AGEGROUP agegroupid="1608" agemax="-1" agemin="-1" name="Visual SB13" handicap="13" />
                <AGEGROUP agegroupid="1609" agemax="-1" agemin="-1" name="Intelectual SB14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3990" />
                    <RANKING order="2" place="-1" resultid="4117" />
                    <RANKING order="3" place="-1" resultid="4120" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1611" agemax="-1" agemin="-1" name="Intelectual SB21 (SD)" handicap="21" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4223" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1766" />
                <TIMESTANDARDREF timestandardlistid="1774" />
                <TIMESTANDARDREF timestandardlistid="1780" />
                <TIMESTANDARDREF timestandardlistid="1786" />
                <TIMESTANDARDREF timestandardlistid="1792" />
                <TIMESTANDARDREF timestandardlistid="1798" />
                <TIMESTANDARDREF timestandardlistid="1804" />
                <TIMESTANDARDREF timestandardlistid="1810" />
                <TIMESTANDARDREF timestandardlistid="1816" />
                <TIMESTANDARDREF timestandardlistid="1822" />
                <TIMESTANDARDREF timestandardlistid="1828" />
                <TIMESTANDARDREF timestandardlistid="1834" />
                <TIMESTANDARDREF timestandardlistid="1840" />
                <TIMESTANDARDREF timestandardlistid="1846" />
                <TIMESTANDARDREF timestandardlistid="1852" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1070" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1708" agemax="-1" agemin="-1" name="Físico-Motora SB4" handicap="4" />
                <AGEGROUP agegroupid="1709" agemax="-1" agemin="-1" name="Físico-Motora SB5" handicap="5" />
                <AGEGROUP agegroupid="1710" agemax="-1" agemin="-1" name="Físico-Motora SB6" handicap="6" />
                <AGEGROUP agegroupid="1711" agemax="-1" agemin="-1" name="Físico-Motora SB7" handicap="7">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4137" />
                    <RANKING order="2" place="2" resultid="3903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1712" agemax="-1" agemin="-1" name="Físico-Motora SB8" handicap="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4114" />
                    <RANKING order="2" place="2" resultid="4024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1713" agemax="-1" agemin="-1" name="Físico-Motora SB9" handicap="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1714" agemax="-1" agemin="-1" name="Físico-Motora SB10" handicap="10" />
                <AGEGROUP agegroupid="1715" agemax="-1" agemin="-1" name="Visual SB11" handicap="11">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3910" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1716" agemax="-1" agemin="-1" name="Visual SB12" handicap="12" />
                <AGEGROUP agegroupid="1717" agemax="-1" agemin="-1" name="Visual SB13" handicap="13" />
                <AGEGROUP agegroupid="1718" agemax="-1" agemin="-1" name="Intelectual SB14" handicap="14" />
                <AGEGROUP agegroupid="1719" agemax="-1" agemin="-1" name="Intelectual SB21 (SD)" handicap="21" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4224" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1764" />
                <TIMESTANDARDREF timestandardlistid="1772" />
                <TIMESTANDARDREF timestandardlistid="1778" />
                <TIMESTANDARDREF timestandardlistid="1784" />
                <TIMESTANDARDREF timestandardlistid="1790" />
                <TIMESTANDARDREF timestandardlistid="1796" />
                <TIMESTANDARDREF timestandardlistid="1802" />
                <TIMESTANDARDREF timestandardlistid="1808" />
                <TIMESTANDARDREF timestandardlistid="1814" />
                <TIMESTANDARDREF timestandardlistid="1820" />
                <TIMESTANDARDREF timestandardlistid="1826" />
                <TIMESTANDARDREF timestandardlistid="1832" />
                <TIMESTANDARDREF timestandardlistid="1838" />
                <TIMESTANDARDREF timestandardlistid="1844" />
                <TIMESTANDARDREF timestandardlistid="1850" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1073" gender="X" number="7" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3178" agemax="-1" agemin="-1" name="MISTO">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4280" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4279" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1075" gender="F" number="8" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1564" agemax="-1" agemin="-1" name="Físico-Motora S1" handicap="1" />
                <AGEGROUP agegroupid="1565" agemax="-1" agemin="-1" name="Físico-Motora S2" handicap="2" />
                <AGEGROUP agegroupid="1566" agemax="-1" agemin="-1" name="Físico-Motora S3" handicap="3" />
                <AGEGROUP agegroupid="1567" agemax="-1" agemin="-1" name="Físico-Motora S4" handicap="4" />
                <AGEGROUP agegroupid="1568" agemax="-1" agemin="-1" name="Físico-Motora S5" handicap="5">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4066" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1569" agemax="-1" agemin="-1" name="Físico-Motora S6" handicap="6">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4161" />
                    <RANKING order="2" place="2" resultid="3938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1570" agemax="-1" agemin="-1" name="Físico-Motora S7" handicap="7" />
                <AGEGROUP agegroupid="1571" agemax="-1" agemin="-1" name="Físico-Motora S8" handicap="8" />
                <AGEGROUP agegroupid="1572" agemax="-1" agemin="-1" name="Físico-Motora S9" handicap="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1573" agemax="-1" agemin="-1" name="Físico-Motora S10" handicap="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4165" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1574" agemax="-1" agemin="-1" name="Visual S11" handicap="11" />
                <AGEGROUP agegroupid="1575" agemax="-1" agemin="-1" name="Visual S12" handicap="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3945" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1576" agemax="-1" agemin="-1" name="Visual S13" handicap="13" />
                <AGEGROUP agegroupid="1577" agemax="-1" agemin="-1" name="Intelectual S14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4104" />
                    <RANKING order="2" place="2" resultid="3967" />
                    <RANKING order="3" place="3" resultid="4141" />
                    <RANKING order="4" place="-1" resultid="4121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1578" agemax="-1" agemin="-1" name="Intelectual S18 (TEA)" handicap="18" />
                <AGEGROUP agegroupid="1579" agemax="-1" agemin="-1" name="Intelectual S21 (SD)" handicap="21" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4225" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4226" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1766" />
                <TIMESTANDARDREF timestandardlistid="1774" />
                <TIMESTANDARDREF timestandardlistid="1780" />
                <TIMESTANDARDREF timestandardlistid="1786" />
                <TIMESTANDARDREF timestandardlistid="1792" />
                <TIMESTANDARDREF timestandardlistid="1798" />
                <TIMESTANDARDREF timestandardlistid="1804" />
                <TIMESTANDARDREF timestandardlistid="1810" />
                <TIMESTANDARDREF timestandardlistid="1816" />
                <TIMESTANDARDREF timestandardlistid="1822" />
                <TIMESTANDARDREF timestandardlistid="1828" />
                <TIMESTANDARDREF timestandardlistid="1834" />
                <TIMESTANDARDREF timestandardlistid="1840" />
                <TIMESTANDARDREF timestandardlistid="1846" />
                <TIMESTANDARDREF timestandardlistid="1852" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1077" gender="M" number="9" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1548" agemax="-1" agemin="-1" name="Físico-Motora S1" handicap="1" />
                <AGEGROUP agegroupid="1549" agemax="-1" agemin="-1" name="Físico-Motora S2" handicap="2" />
                <AGEGROUP agegroupid="1550" agemax="-1" agemin="-1" name="Físico-Motora S3" handicap="3" />
                <AGEGROUP agegroupid="1551" agemax="-1" agemin="-1" name="Físico-Motora S4" handicap="4" />
                <AGEGROUP agegroupid="1552" agemax="-1" agemin="-1" name="Físico-Motora S5" handicap="5" />
                <AGEGROUP agegroupid="1553" agemax="-1" agemin="-1" name="Físico-Motora S6" handicap="6">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1554" agemax="-1" agemin="-1" name="Físico-Motora S7" handicap="7">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4149" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1555" agemax="-1" agemin="-1" name="Físico-Motora S8" handicap="8" />
                <AGEGROUP agegroupid="1556" agemax="-1" agemin="-1" name="Físico-Motora S9" handicap="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3881" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1557" agemax="-1" agemin="-1" name="Físico-Motora S10" handicap="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1558" agemax="-1" agemin="-1" name="Visual S11" handicap="11" />
                <AGEGROUP agegroupid="1559" agemax="-1" agemin="-1" name="Visual S12" handicap="12" />
                <AGEGROUP agegroupid="1560" agemax="-1" agemin="-1" name="Visual S13" handicap="13" />
                <AGEGROUP agegroupid="1561" agemax="-1" agemin="-1" name="Intelectual S14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4048" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1562" agemax="-1" agemin="-1" name="Intelectual S18 (TEA)" handicap="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4055" />
                    <RANKING order="2" place="2" resultid="3973" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1563" agemax="-1" agemin="-1" name="Intelectual S21 (SD)" handicap="21">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4087" />
                    <RANKING order="2" place="2" resultid="3958" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4227" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4228" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1764" />
                <TIMESTANDARDREF timestandardlistid="1772" />
                <TIMESTANDARDREF timestandardlistid="1778" />
                <TIMESTANDARDREF timestandardlistid="1784" />
                <TIMESTANDARDREF timestandardlistid="1790" />
                <TIMESTANDARDREF timestandardlistid="1796" />
                <TIMESTANDARDREF timestandardlistid="1802" />
                <TIMESTANDARDREF timestandardlistid="1808" />
                <TIMESTANDARDREF timestandardlistid="1814" />
                <TIMESTANDARDREF timestandardlistid="1820" />
                <TIMESTANDARDREF timestandardlistid="1826" />
                <TIMESTANDARDREF timestandardlistid="1832" />
                <TIMESTANDARDREF timestandardlistid="1838" />
                <TIMESTANDARDREF timestandardlistid="1844" />
                <TIMESTANDARDREF timestandardlistid="1850" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1079" gender="F" number="10" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1537" agemax="-1" agemin="-1" name="Físico-Motora S6" handicap="6">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4091" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1538" agemax="-1" agemin="-1" name="Físico-Motora S7" handicap="7" />
                <AGEGROUP agegroupid="1539" agemax="-1" agemin="-1" name="Físico-Motora S8" handicap="8" />
                <AGEGROUP agegroupid="1540" agemax="-1" agemin="-1" name="Físico-Motora S9" handicap="9" />
                <AGEGROUP agegroupid="1541" agemax="-1" agemin="-1" name="Físico-Motora S10" handicap="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1542" agemax="-1" agemin="-1" name="Visual S11" handicap="11" />
                <AGEGROUP agegroupid="1543" agemax="-1" agemin="-1" name="Visual S12" handicap="12" />
                <AGEGROUP agegroupid="1544" agemax="-1" agemin="-1" name="Visual S13" handicap="13" />
                <AGEGROUP agegroupid="1545" agemax="-1" agemin="-1" name="Intelectual S14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4103" />
                    <RANKING order="2" place="2" resultid="3989" />
                    <RANKING order="3" place="3" resultid="4039" />
                    <RANKING order="4" place="-1" resultid="4116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4296" agemax="-1" agemin="-1" name="Intelectual S18 (TEA)" handicap="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1547" agemax="-1" agemin="-1" name="Intelectual S21 (SD)" handicap="21" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4229" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1766" />
                <TIMESTANDARDREF timestandardlistid="1774" />
                <TIMESTANDARDREF timestandardlistid="1780" />
                <TIMESTANDARDREF timestandardlistid="1786" />
                <TIMESTANDARDREF timestandardlistid="1792" />
                <TIMESTANDARDREF timestandardlistid="1798" />
                <TIMESTANDARDREF timestandardlistid="1804" />
                <TIMESTANDARDREF timestandardlistid="1810" />
                <TIMESTANDARDREF timestandardlistid="1816" />
                <TIMESTANDARDREF timestandardlistid="1822" />
                <TIMESTANDARDREF timestandardlistid="1828" />
                <TIMESTANDARDREF timestandardlistid="1834" />
                <TIMESTANDARDREF timestandardlistid="1840" />
                <TIMESTANDARDREF timestandardlistid="1846" />
                <TIMESTANDARDREF timestandardlistid="1852" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1081" gender="M" number="11" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="4297" agemax="-1" agemin="-1" name="Físico-Motora S6" handicap="6">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4298" agemax="-1" agemin="-1" name="Físico-Motora S7" handicap="7" />
                <AGEGROUP agegroupid="4299" agemax="-1" agemin="-1" name="Físico-Motora S8" handicap="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4169" />
                    <RANKING order="2" place="2" resultid="3981" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4300" agemax="-1" agemin="-1" name="Físico-Motora S9" handicap="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4301" agemax="-1" agemin="-1" name="Físico-Motora S10" handicap="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3941" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4302" agemax="-1" agemin="-1" name="Visual S11" handicap="11">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4174" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4303" agemax="-1" agemin="-1" name="Visual S12" handicap="12" />
                <AGEGROUP agegroupid="4304" agemax="-1" agemin="-1" name="Visual S13" handicap="13" />
                <AGEGROUP agegroupid="4305" agemax="-1" agemin="-1" name="Intelectual S14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3929" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4306" agemax="-1" agemin="-1" name="Intelectual S18 (TEA)" handicap="18">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4128" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="4307" agemax="-1" agemin="-1" name="Intelectual S21 (SD)" handicap="21">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3961" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4230" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4231" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1764" />
                <TIMESTANDARDREF timestandardlistid="1772" />
                <TIMESTANDARDREF timestandardlistid="1778" />
                <TIMESTANDARDREF timestandardlistid="1784" />
                <TIMESTANDARDREF timestandardlistid="1790" />
                <TIMESTANDARDREF timestandardlistid="1796" />
                <TIMESTANDARDREF timestandardlistid="1802" />
                <TIMESTANDARDREF timestandardlistid="1808" />
                <TIMESTANDARDREF timestandardlistid="1814" />
                <TIMESTANDARDREF timestandardlistid="1820" />
                <TIMESTANDARDREF timestandardlistid="1826" />
                <TIMESTANDARDREF timestandardlistid="1832" />
                <TIMESTANDARDREF timestandardlistid="1838" />
                <TIMESTANDARDREF timestandardlistid="1844" />
                <TIMESTANDARDREF timestandardlistid="1850" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1084" gender="F" number="12" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1085" agemax="-1" agemin="-1" name="DF">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4260" />
                    <RANKING order="2" place="2" resultid="4262" />
                    <RANKING order="3" place="-1" resultid="4261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3152" agemax="-1" agemin="-1" name="DV">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4260" />
                    <RANKING order="2" place="2" resultid="4262" />
                    <RANKING order="3" place="-1" resultid="4261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3153" agemax="-1" agemin="-1" name="DI">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4260" />
                    <RANKING order="2" place="2" resultid="4262" />
                    <RANKING order="3" place="-1" resultid="4261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3155" agemax="-1" agemin="-1" name="SD">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4260" />
                    <RANKING order="2" place="2" resultid="4262" />
                    <RANKING order="3" place="-1" resultid="4261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3156" agemax="-1" agemin="-1" name="DEA">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4260" />
                    <RANKING order="2" place="2" resultid="4262" />
                    <RANKING order="3" place="-1" resultid="4261" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4259" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1766" />
                <TIMESTANDARDREF timestandardlistid="1774" />
                <TIMESTANDARDREF timestandardlistid="1780" />
                <TIMESTANDARDREF timestandardlistid="1786" />
                <TIMESTANDARDREF timestandardlistid="1792" />
                <TIMESTANDARDREF timestandardlistid="1798" />
                <TIMESTANDARDREF timestandardlistid="1804" />
                <TIMESTANDARDREF timestandardlistid="1810" />
                <TIMESTANDARDREF timestandardlistid="1816" />
                <TIMESTANDARDREF timestandardlistid="1822" />
                <TIMESTANDARDREF timestandardlistid="1828" />
                <TIMESTANDARDREF timestandardlistid="1834" />
                <TIMESTANDARDREF timestandardlistid="1840" />
                <TIMESTANDARDREF timestandardlistid="1846" />
                <TIMESTANDARDREF timestandardlistid="1852" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1086" gender="M" number="13" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3158" agemax="-1" agemin="-1" name="DF">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4266" />
                    <RANKING order="2" place="2" resultid="4267" />
                    <RANKING order="3" place="3" resultid="4265" />
                    <RANKING order="4" place="-1" resultid="4264" />
                    <RANKING order="5" place="-1" resultid="4268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3159" agemax="-1" agemin="-1" name="DV">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4266" />
                    <RANKING order="2" place="2" resultid="4267" />
                    <RANKING order="3" place="3" resultid="4265" />
                    <RANKING order="4" place="-1" resultid="4264" />
                    <RANKING order="5" place="-1" resultid="4268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3160" agemax="-1" agemin="-1" name="DI">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4266" />
                    <RANKING order="2" place="2" resultid="4267" />
                    <RANKING order="3" place="3" resultid="4265" />
                    <RANKING order="4" place="-1" resultid="4264" />
                    <RANKING order="5" place="-1" resultid="4268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3161" agemax="-1" agemin="-1" name="SD">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4266" />
                    <RANKING order="2" place="2" resultid="4267" />
                    <RANKING order="3" place="3" resultid="4265" />
                    <RANKING order="4" place="-1" resultid="4264" />
                    <RANKING order="5" place="-1" resultid="4268" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3162" agemax="-1" agemin="-1" name="DEA">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4266" />
                    <RANKING order="2" place="2" resultid="4267" />
                    <RANKING order="3" place="3" resultid="4265" />
                    <RANKING order="4" place="-1" resultid="4264" />
                    <RANKING order="5" place="-1" resultid="4268" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4263" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1764" />
                <TIMESTANDARDREF timestandardlistid="1772" />
                <TIMESTANDARDREF timestandardlistid="1778" />
                <TIMESTANDARDREF timestandardlistid="1784" />
                <TIMESTANDARDREF timestandardlistid="1790" />
                <TIMESTANDARDREF timestandardlistid="1796" />
                <TIMESTANDARDREF timestandardlistid="1802" />
                <TIMESTANDARDREF timestandardlistid="1808" />
                <TIMESTANDARDREF timestandardlistid="1814" />
                <TIMESTANDARDREF timestandardlistid="1820" />
                <TIMESTANDARDREF timestandardlistid="1826" />
                <TIMESTANDARDREF timestandardlistid="1832" />
                <TIMESTANDARDREF timestandardlistid="1838" />
                <TIMESTANDARDREF timestandardlistid="1844" />
                <TIMESTANDARDREF timestandardlistid="1850" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-05-30" daytime="15:30" endtime="17:49" number="2" officialmeeting="15:00" warmupfrom="14:30" warmupuntil="15:20">
          <EVENTS>
            <EVENT eventid="1088" gender="F" number="14" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1504" agemax="-1" agemin="-1" name="Físico-Motora SM5" handicap="5" />
                <AGEGROUP agegroupid="1505" agemax="-1" agemin="-1" name="Físico-Motora SM6" handicap="6">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4093" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1506" agemax="-1" agemin="-1" name="Físico-Motora SM7" handicap="7" />
                <AGEGROUP agegroupid="1507" agemax="-1" agemin="-1" name="Físico-Motora SM8" handicap="8" />
                <AGEGROUP agegroupid="1508" agemax="-1" agemin="-1" name="Físico-Motora SM9" handicap="9" />
                <AGEGROUP agegroupid="1509" agemax="-1" agemin="-1" name="Físico-Motora SM10" handicap="10" />
                <AGEGROUP agegroupid="1510" agemax="-1" agemin="-1" name="Visual SM11" handicap="11" />
                <AGEGROUP agegroupid="1511" agemax="-1" agemin="-1" name="Visual SM12" handicap="12" />
                <AGEGROUP agegroupid="1512" agemax="-1" agemin="-1" name="Visual SM13" handicap="13" />
                <AGEGROUP agegroupid="1513" agemax="-1" agemin="-1" name="Intelectual SM14" handicap="14" />
                <AGEGROUP agegroupid="1515" agemax="-1" agemin="-1" name="Intelectual SM21 (SD)" handicap="21" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4232" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1766" />
                <TIMESTANDARDREF timestandardlistid="1774" />
                <TIMESTANDARDREF timestandardlistid="1780" />
                <TIMESTANDARDREF timestandardlistid="1786" />
                <TIMESTANDARDREF timestandardlistid="1792" />
                <TIMESTANDARDREF timestandardlistid="1798" />
                <TIMESTANDARDREF timestandardlistid="1804" />
                <TIMESTANDARDREF timestandardlistid="1810" />
                <TIMESTANDARDREF timestandardlistid="1816" />
                <TIMESTANDARDREF timestandardlistid="1822" />
                <TIMESTANDARDREF timestandardlistid="1828" />
                <TIMESTANDARDREF timestandardlistid="1834" />
                <TIMESTANDARDREF timestandardlistid="1840" />
                <TIMESTANDARDREF timestandardlistid="1846" />
                <TIMESTANDARDREF timestandardlistid="1852" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1090" gender="M" number="15" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1730" agemax="-1" agemin="-1" name="Físico-Motora SM5" handicap="5" />
                <AGEGROUP agegroupid="1731" agemax="-1" agemin="-1" name="Físico-Motora SM6" handicap="6" />
                <AGEGROUP agegroupid="1732" agemax="-1" agemin="-1" name="Físico-Motora SM7" handicap="7" />
                <AGEGROUP agegroupid="1733" agemax="-1" agemin="-1" name="Físico-Motora SM8" handicap="8" />
                <AGEGROUP agegroupid="1734" agemax="-1" agemin="-1" name="Físico-Motora SM9" handicap="9" />
                <AGEGROUP agegroupid="1735" agemax="-1" agemin="-1" name="Físico-Motora SM10" handicap="10" />
                <AGEGROUP agegroupid="1736" agemax="-1" agemin="-1" name="Visual SM11" handicap="11" />
                <AGEGROUP agegroupid="1737" agemax="-1" agemin="-1" name="Visual SM12" handicap="12" />
                <AGEGROUP agegroupid="1738" agemax="-1" agemin="-1" name="Visual SM13" handicap="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1739" agemax="-1" agemin="-1" name="Intelectual SM14" handicap="14" />
                <AGEGROUP agegroupid="1740" agemax="-1" agemin="-1" name="Intelectual SM21 (SD)" handicap="21" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4233" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1764" />
                <TIMESTANDARDREF timestandardlistid="1772" />
                <TIMESTANDARDREF timestandardlistid="1778" />
                <TIMESTANDARDREF timestandardlistid="1784" />
                <TIMESTANDARDREF timestandardlistid="1790" />
                <TIMESTANDARDREF timestandardlistid="1796" />
                <TIMESTANDARDREF timestandardlistid="1802" />
                <TIMESTANDARDREF timestandardlistid="1808" />
                <TIMESTANDARDREF timestandardlistid="1814" />
                <TIMESTANDARDREF timestandardlistid="1820" />
                <TIMESTANDARDREF timestandardlistid="1826" />
                <TIMESTANDARDREF timestandardlistid="1832" />
                <TIMESTANDARDREF timestandardlistid="1838" />
                <TIMESTANDARDREF timestandardlistid="1844" />
                <TIMESTANDARDREF timestandardlistid="1850" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1092" gender="F" number="16" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="150" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1741" agemax="-1" agemin="-1" name="Físico-Motora SM3" handicap="3" />
                <AGEGROUP agegroupid="1742" agemax="-1" agemin="-1" name="Físico-Motora SM3" handicap="3" />
              </AGEGROUPS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1766" />
                <TIMESTANDARDREF timestandardlistid="1774" />
                <TIMESTANDARDREF timestandardlistid="1780" />
                <TIMESTANDARDREF timestandardlistid="1786" />
                <TIMESTANDARDREF timestandardlistid="1792" />
                <TIMESTANDARDREF timestandardlistid="1798" />
                <TIMESTANDARDREF timestandardlistid="1804" />
                <TIMESTANDARDREF timestandardlistid="1810" />
                <TIMESTANDARDREF timestandardlistid="1816" />
                <TIMESTANDARDREF timestandardlistid="1822" />
                <TIMESTANDARDREF timestandardlistid="1828" />
                <TIMESTANDARDREF timestandardlistid="1834" />
                <TIMESTANDARDREF timestandardlistid="1840" />
                <TIMESTANDARDREF timestandardlistid="1846" />
                <TIMESTANDARDREF timestandardlistid="1852" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1094" gender="M" number="17" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="150" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1752" agemax="-1" agemin="-1" name="Físico-Motora SM3" handicap="3" />
                <AGEGROUP agegroupid="1753" agemax="-1" agemin="-1" name="Físico-Motora SM3" handicap="3" />
              </AGEGROUPS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1764" />
                <TIMESTANDARDREF timestandardlistid="1772" />
                <TIMESTANDARDREF timestandardlistid="1778" />
                <TIMESTANDARDREF timestandardlistid="1784" />
                <TIMESTANDARDREF timestandardlistid="1790" />
                <TIMESTANDARDREF timestandardlistid="1796" />
                <TIMESTANDARDREF timestandardlistid="1802" />
                <TIMESTANDARDREF timestandardlistid="1808" />
                <TIMESTANDARDREF timestandardlistid="1814" />
                <TIMESTANDARDREF timestandardlistid="1820" />
                <TIMESTANDARDREF timestandardlistid="1826" />
                <TIMESTANDARDREF timestandardlistid="1832" />
                <TIMESTANDARDREF timestandardlistid="1838" />
                <TIMESTANDARDREF timestandardlistid="1844" />
                <TIMESTANDARDREF timestandardlistid="1850" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1096" gender="F" number="18" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1436" agemax="-1" agemin="-1" name="Físico-Motora S1" handicap="1" />
                <AGEGROUP agegroupid="1437" agemax="-1" agemin="-1" name="Físico-Motora S2" handicap="2" />
                <AGEGROUP agegroupid="1438" agemax="-1" agemin="-1" name="Físico-Motora S3" handicap="3" />
                <AGEGROUP agegroupid="1439" agemax="-1" agemin="-1" name="Físico-Motora S4" handicap="4" />
                <AGEGROUP agegroupid="1440" agemax="-1" agemin="-1" name="Físico-Motora S5" handicap="5">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1441" agemax="-1" agemin="-1" name="Físico-Motora S6" handicap="6">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4162" />
                    <RANKING order="2" place="2" resultid="4060" />
                    <RANKING order="3" place="3" resultid="3939" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1442" agemax="-1" agemin="-1" name="Físico-Motora S7" handicap="7">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4037" />
                    <RANKING order="2" place="2" resultid="3986" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1443" agemax="-1" agemin="-1" name="Físico-Motora S8" handicap="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4154" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1444" agemax="-1" agemin="-1" name="Físico-Motora S9" handicap="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4010" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1445" agemax="-1" agemin="-1" name="Físico-Motora S10" handicap="10">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4166" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1446" agemax="-1" agemin="-1" name="Visual S11" handicap="11" />
                <AGEGROUP agegroupid="1447" agemax="-1" agemin="-1" name="Visual S12" handicap="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1448" agemax="-1" agemin="-1" name="Visual S13" handicap="13" />
                <AGEGROUP agegroupid="1449" agemax="-1" agemin="-1" name="Intelectual S14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4134" />
                    <RANKING order="2" place="2" resultid="3998" />
                    <RANKING order="3" place="3" resultid="4063" />
                    <RANKING order="4" place="4" resultid="4142" />
                    <RANKING order="5" place="-1" resultid="4122" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1450" agemax="-1" agemin="-1" name="Intelectual S18 (TEA)" handicap="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4146" />
                    <RANKING order="2" place="2" resultid="4100" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1451" agemax="-1" agemin="-1" name="Intelectual S21 (SD)" handicap="21">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4003" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4234" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4235" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4236" number="3" order="3" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1766" />
                <TIMESTANDARDREF timestandardlistid="1774" />
                <TIMESTANDARDREF timestandardlistid="1780" />
                <TIMESTANDARDREF timestandardlistid="1786" />
                <TIMESTANDARDREF timestandardlistid="1792" />
                <TIMESTANDARDREF timestandardlistid="1798" />
                <TIMESTANDARDREF timestandardlistid="1804" />
                <TIMESTANDARDREF timestandardlistid="1810" />
                <TIMESTANDARDREF timestandardlistid="1816" />
                <TIMESTANDARDREF timestandardlistid="1822" />
                <TIMESTANDARDREF timestandardlistid="1828" />
                <TIMESTANDARDREF timestandardlistid="1834" />
                <TIMESTANDARDREF timestandardlistid="1840" />
                <TIMESTANDARDREF timestandardlistid="1846" />
                <TIMESTANDARDREF timestandardlistid="1852" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1098" gender="M" number="19" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1420" agemax="-1" agemin="-1" name="Físico-Motora S1" handicap="1" />
                <AGEGROUP agegroupid="1421" agemax="-1" agemin="-1" name="Físico-Motora S2" handicap="2" />
                <AGEGROUP agegroupid="1422" agemax="-1" agemin="-1" name="Físico-Motora S3" handicap="3" />
                <AGEGROUP agegroupid="1423" agemax="-1" agemin="-1" name="Físico-Motora S4" handicap="4">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3900" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1424" agemax="-1" agemin="-1" name="Físico-Motora S5" handicap="5">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1425" agemax="-1" agemin="-1" name="Físico-Motora S6" handicap="6">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3950" />
                    <RANKING order="2" place="2" resultid="3859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1426" agemax="-1" agemin="-1" name="Físico-Motora S7" handicap="7">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4150" />
                    <RANKING order="2" place="2" resultid="3904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1427" agemax="-1" agemin="-1" name="Físico-Motora S8" handicap="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4138" />
                    <RANKING order="2" place="2" resultid="4126" />
                    <RANKING order="3" place="3" resultid="4171" />
                    <RANKING order="4" place="4" resultid="3983" />
                    <RANKING order="5" place="-1" resultid="3955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1428" agemax="-1" agemin="-1" name="Físico-Motora S9" handicap="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3882" />
                    <RANKING order="2" place="2" resultid="4025" />
                    <RANKING order="3" place="3" resultid="3864" />
                    <RANKING order="4" place="4" resultid="3868" />
                    <RANKING order="5" place="5" resultid="3926" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1429" agemax="-1" agemin="-1" name="Físico-Motora S10" handicap="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3892" />
                    <RANKING order="2" place="2" resultid="3943" />
                    <RANKING order="3" place="-1" resultid="3918" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1430" agemax="-1" agemin="-1" name="Visual S11" handicap="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4083" />
                    <RANKING order="2" place="2" resultid="4072" />
                    <RANKING order="3" place="3" resultid="4176" />
                    <RANKING order="4" place="-1" resultid="3911" />
                    <RANKING order="5" place="-1" resultid="4076" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1431" agemax="-1" agemin="-1" name="Visual S12" handicap="12">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4006" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1432" agemax="-1" agemin="-1" name="Visual S13" handicap="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3877" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1433" agemax="-1" agemin="-1" name="Intelectual S14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4109" />
                    <RANKING order="2" place="2" resultid="4051" />
                    <RANKING order="3" place="3" resultid="3923" />
                    <RANKING order="4" place="4" resultid="4181" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1434" agemax="-1" agemin="-1" name="Intelectual S18 (TEA)" handicap="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4081" />
                    <RANKING order="2" place="2" resultid="3975" />
                    <RANKING order="3" place="3" resultid="4043" />
                    <RANKING order="4" place="4" resultid="4096" />
                    <RANKING order="5" place="-1" resultid="3916" />
                    <RANKING order="6" place="-1" resultid="4129" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1435" agemax="-1" agemin="-1" name="Intelectual S21 (SD)" handicap="21">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4158" />
                    <RANKING order="2" place="2" resultid="4089" />
                    <RANKING order="3" place="3" resultid="3959" />
                    <RANKING order="4" place="4" resultid="3872" />
                    <RANKING order="5" place="5" resultid="4021" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4237" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4238" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4239" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4240" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4241" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="4242" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="4243" number="7" order="7" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1764" />
                <TIMESTANDARDREF timestandardlistid="1772" />
                <TIMESTANDARDREF timestandardlistid="1778" />
                <TIMESTANDARDREF timestandardlistid="1784" />
                <TIMESTANDARDREF timestandardlistid="1790" />
                <TIMESTANDARDREF timestandardlistid="1796" />
                <TIMESTANDARDREF timestandardlistid="1802" />
                <TIMESTANDARDREF timestandardlistid="1808" />
                <TIMESTANDARDREF timestandardlistid="1814" />
                <TIMESTANDARDREF timestandardlistid="1820" />
                <TIMESTANDARDREF timestandardlistid="1826" />
                <TIMESTANDARDREF timestandardlistid="1832" />
                <TIMESTANDARDREF timestandardlistid="1838" />
                <TIMESTANDARDREF timestandardlistid="1844" />
                <TIMESTANDARDREF timestandardlistid="1850" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1100" gender="F" number="20" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1411" agemax="-1" agemin="-1" name="Físico-Motora S8" handicap="8" />
                <AGEGROUP agegroupid="1412" agemax="-1" agemin="-1" name="Físico-Motora S9" handicap="9" />
                <AGEGROUP agegroupid="1413" agemax="-1" agemin="-1" name="Físico-Motora S10" handicap="10" />
                <AGEGROUP agegroupid="1414" agemax="-1" agemin="-1" name="Visual S11" handicap="11" />
                <AGEGROUP agegroupid="1415" agemax="-1" agemin="-1" name="Visual S12" handicap="12" />
                <AGEGROUP agegroupid="1416" agemax="-1" agemin="-1" name="Visual S13" handicap="13" />
                <AGEGROUP agegroupid="1417" agemax="-1" agemin="-1" name="Intelectual S14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4132" />
                    <RANKING order="2" place="2" resultid="4102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1419" agemax="-1" agemin="-1" name="Intelectual S21 (SD)" handicap="21" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4244" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1766" />
                <TIMESTANDARDREF timestandardlistid="1774" />
                <TIMESTANDARDREF timestandardlistid="1780" />
                <TIMESTANDARDREF timestandardlistid="1786" />
                <TIMESTANDARDREF timestandardlistid="1792" />
                <TIMESTANDARDREF timestandardlistid="1798" />
                <TIMESTANDARDREF timestandardlistid="1804" />
                <TIMESTANDARDREF timestandardlistid="1810" />
                <TIMESTANDARDREF timestandardlistid="1816" />
                <TIMESTANDARDREF timestandardlistid="1822" />
                <TIMESTANDARDREF timestandardlistid="1828" />
                <TIMESTANDARDREF timestandardlistid="1834" />
                <TIMESTANDARDREF timestandardlistid="1840" />
                <TIMESTANDARDREF timestandardlistid="1846" />
                <TIMESTANDARDREF timestandardlistid="1852" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1102" gender="M" number="21" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1754" agemax="-1" agemin="-1" name="Físico-Motora S8" handicap="8" />
                <AGEGROUP agegroupid="1755" agemax="-1" agemin="-1" name="Físico-Motora S9" handicap="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4112" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1756" agemax="-1" agemin="-1" name="Físico-Motora S10" handicap="10" />
                <AGEGROUP agegroupid="1757" agemax="-1" agemin="-1" name="Visual S11" handicap="11" />
                <AGEGROUP agegroupid="1758" agemax="-1" agemin="-1" name="Visual S12" handicap="12" />
                <AGEGROUP agegroupid="1759" agemax="-1" agemin="-1" name="Visual S13" handicap="13" />
                <AGEGROUP agegroupid="1760" agemax="-1" agemin="-1" name="Intelectual S14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1761" agemax="-1" agemin="-1" name="Intelectual S21 (SD)" handicap="21" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4245" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1764" />
                <TIMESTANDARDREF timestandardlistid="1772" />
                <TIMESTANDARDREF timestandardlistid="1778" />
                <TIMESTANDARDREF timestandardlistid="1784" />
                <TIMESTANDARDREF timestandardlistid="1790" />
                <TIMESTANDARDREF timestandardlistid="1796" />
                <TIMESTANDARDREF timestandardlistid="1802" />
                <TIMESTANDARDREF timestandardlistid="1808" />
                <TIMESTANDARDREF timestandardlistid="1814" />
                <TIMESTANDARDREF timestandardlistid="1820" />
                <TIMESTANDARDREF timestandardlistid="1826" />
                <TIMESTANDARDREF timestandardlistid="1832" />
                <TIMESTANDARDREF timestandardlistid="1838" />
                <TIMESTANDARDREF timestandardlistid="1844" />
                <TIMESTANDARDREF timestandardlistid="1850" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1105" gender="F" number="22" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1676" agemax="-1" agemin="-1" name="Físico-Motora SB1" handicap="1" />
                <AGEGROUP agegroupid="1677" agemax="-1" agemin="-1" name="Físico-Motora SB2" handicap="2" />
                <AGEGROUP agegroupid="1678" agemax="-1" agemin="-1" name="Físico-Motora SB3" handicap="3" />
                <AGEGROUP agegroupid="1679" agemax="-1" agemin="-1" name="Físico-Motora SB4" handicap="4" />
                <AGEGROUP agegroupid="1680" agemax="-1" agemin="-1" name="Físico-Motora SB5" handicap="5">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1681" agemax="-1" agemin="-1" name="Físico-Motora SB6" handicap="6" />
                <AGEGROUP agegroupid="1682" agemax="-1" agemin="-1" name="Físico-Motora SB7" handicap="7" />
                <AGEGROUP agegroupid="1683" agemax="-1" agemin="-1" name="Físico-Motora SB8" handicap="8" />
                <AGEGROUP agegroupid="1684" agemax="-1" agemin="-1" name="Físico-Motora SB9" handicap="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3897" />
                    <RANKING order="2" place="2" resultid="4011" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1685" agemax="-1" agemin="-1" name="Físico-Motora SB10" handicap="10" />
                <AGEGROUP agegroupid="1686" agemax="-1" agemin="-1" name="Visual SB11" handicap="11" />
                <AGEGROUP agegroupid="1687" agemax="-1" agemin="-1" name="Visual SB12" handicap="12" />
                <AGEGROUP agegroupid="1688" agemax="-1" agemin="-1" name="Visual SB13" handicap="13" />
                <AGEGROUP agegroupid="1689" agemax="-1" agemin="-1" name="Intelectual SB14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3999" />
                    <RANKING order="2" place="2" resultid="4064" />
                    <RANKING order="3" place="-1" resultid="4118" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1690" agemax="-1" agemin="-1" name="Intelectual SB18 (TEA)" handicap="18" />
                <AGEGROUP agegroupid="1691" agemax="-1" agemin="-1" name="Intelectual SB21 (SD)" handicap="21" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4246" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1766" />
                <TIMESTANDARDREF timestandardlistid="1774" />
                <TIMESTANDARDREF timestandardlistid="1780" />
                <TIMESTANDARDREF timestandardlistid="1786" />
                <TIMESTANDARDREF timestandardlistid="1792" />
                <TIMESTANDARDREF timestandardlistid="1798" />
                <TIMESTANDARDREF timestandardlistid="1804" />
                <TIMESTANDARDREF timestandardlistid="1810" />
                <TIMESTANDARDREF timestandardlistid="1816" />
                <TIMESTANDARDREF timestandardlistid="1822" />
                <TIMESTANDARDREF timestandardlistid="1828" />
                <TIMESTANDARDREF timestandardlistid="1834" />
                <TIMESTANDARDREF timestandardlistid="1840" />
                <TIMESTANDARDREF timestandardlistid="1846" />
                <TIMESTANDARDREF timestandardlistid="1852" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1107" gender="M" number="23" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1692" agemax="-1" agemin="-1" name="Físico-Motora SB1" handicap="1" />
                <AGEGROUP agegroupid="1693" agemax="-1" agemin="-1" name="Físico-Motora SB2" handicap="2" />
                <AGEGROUP agegroupid="1694" agemax="-1" agemin="-1" name="Físico-Motora SB3" handicap="3">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3901" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1695" agemax="-1" agemin="-1" name="Físico-Motora SB4" handicap="4" />
                <AGEGROUP agegroupid="1696" agemax="-1" agemin="-1" name="Físico-Motora SB5" handicap="5">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3995" />
                    <RANKING order="2" place="-1" resultid="3951" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1697" agemax="-1" agemin="-1" name="Físico-Motora SB6" handicap="6">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4029" />
                    <RANKING order="2" place="-1" resultid="3860" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1698" agemax="-1" agemin="-1" name="Físico-Motora SB7" handicap="7">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1699" agemax="-1" agemin="-1" name="Físico-Motora SB8" handicap="8">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3927" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1700" agemax="-1" agemin="-1" name="Físico-Motora SB9" handicap="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3888" />
                    <RANKING order="2" place="-1" resultid="3869" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1701" agemax="-1" agemin="-1" name="Físico-Motora SB10" handicap="10" />
                <AGEGROUP agegroupid="1702" agemax="-1" agemin="-1" name="Visual SB11" handicap="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4084" />
                    <RANKING order="2" place="-1" resultid="3912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1703" agemax="-1" agemin="-1" name="Visual SB12" handicap="12">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4007" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1704" agemax="-1" agemin="-1" name="Visual SB13" handicap="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1705" agemax="-1" agemin="-1" name="Intelectual SB14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="4052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1706" agemax="-1" agemin="-1" name="Intelectual SB18 (TEA)" handicap="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4056" />
                    <RANKING order="2" place="2" resultid="4044" />
                    <RANKING order="3" place="-1" resultid="4130" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1707" agemax="-1" agemin="-1" name="Intelectual SB21 (SD)" handicap="21">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3873" />
                    <RANKING order="2" place="-1" resultid="3963" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4247" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4248" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4249" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4250" number="4" order="4" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1764" />
                <TIMESTANDARDREF timestandardlistid="1772" />
                <TIMESTANDARDREF timestandardlistid="1778" />
                <TIMESTANDARDREF timestandardlistid="1784" />
                <TIMESTANDARDREF timestandardlistid="1790" />
                <TIMESTANDARDREF timestandardlistid="1796" />
                <TIMESTANDARDREF timestandardlistid="1802" />
                <TIMESTANDARDREF timestandardlistid="1808" />
                <TIMESTANDARDREF timestandardlistid="1814" />
                <TIMESTANDARDREF timestandardlistid="1820" />
                <TIMESTANDARDREF timestandardlistid="1826" />
                <TIMESTANDARDREF timestandardlistid="1832" />
                <TIMESTANDARDREF timestandardlistid="1838" />
                <TIMESTANDARDREF timestandardlistid="1844" />
                <TIMESTANDARDREF timestandardlistid="1850" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1109" gender="F" number="24" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1340" agemax="-1" agemin="-1" name="Físico-Motora S1" handicap="1" />
                <AGEGROUP agegroupid="1341" agemax="-1" agemin="-1" name="Físico-Motora S2" handicap="2" />
                <AGEGROUP agegroupid="1342" agemax="-1" agemin="-1" name="Físico-Motora S3" handicap="3" />
                <AGEGROUP agegroupid="1343" agemax="-1" agemin="-1" name="Físico-Motora S4" handicap="4" />
                <AGEGROUP agegroupid="1344" agemax="-1" agemin="-1" name="Físico-Motora S5" handicap="5" />
                <AGEGROUP agegroupid="1345" agemax="-1" agemin="-1" name="Físico-Motora S6" handicap="6">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4160" />
                    <RANKING order="2" place="2" resultid="4058" />
                    <RANKING order="3" place="3" resultid="3937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1346" agemax="-1" agemin="-1" name="Físico-Motora S7" handicap="7">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4035" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1347" agemax="-1" agemin="-1" name="Físico-Motora S8" handicap="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4152" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1348" agemax="-1" agemin="-1" name="Físico-Motora S9" handicap="9" />
                <AGEGROUP agegroupid="1349" agemax="-1" agemin="-1" name="Físico-Motora S10" handicap="10" />
                <AGEGROUP agegroupid="1350" agemax="-1" agemin="-1" name="Visual S11" handicap="11" />
                <AGEGROUP agegroupid="1351" agemax="-1" agemin="-1" name="Visual S12" handicap="12" />
                <AGEGROUP agegroupid="1352" agemax="-1" agemin="-1" name="Visual S13" handicap="13" />
                <AGEGROUP agegroupid="1353" agemax="-1" agemin="-1" name="Intelectual S14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4133" />
                    <RANKING order="2" place="2" resultid="3965" />
                    <RANKING order="3" place="3" resultid="4140" />
                    <RANKING order="4" place="4" resultid="4062" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1354" agemax="-1" agemin="-1" name="Intelectual S18 (TEA)" handicap="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4145" />
                    <RANKING order="2" place="2" resultid="4098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1355" agemax="-1" agemin="-1" name="Intelectual S21 (SD)" handicap="21">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4001" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4251" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4252" number="2" order="2" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1766" />
                <TIMESTANDARDREF timestandardlistid="1774" />
                <TIMESTANDARDREF timestandardlistid="1780" />
                <TIMESTANDARDREF timestandardlistid="1786" />
                <TIMESTANDARDREF timestandardlistid="1792" />
                <TIMESTANDARDREF timestandardlistid="1798" />
                <TIMESTANDARDREF timestandardlistid="1804" />
                <TIMESTANDARDREF timestandardlistid="1810" />
                <TIMESTANDARDREF timestandardlistid="1816" />
                <TIMESTANDARDREF timestandardlistid="1822" />
                <TIMESTANDARDREF timestandardlistid="1828" />
                <TIMESTANDARDREF timestandardlistid="1834" />
                <TIMESTANDARDREF timestandardlistid="1840" />
                <TIMESTANDARDREF timestandardlistid="1846" />
                <TIMESTANDARDREF timestandardlistid="1852" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1111" gender="M" number="25" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1324" agemax="-1" agemin="-1" name="Físico-Motora S1" handicap="1" />
                <AGEGROUP agegroupid="1325" agemax="-1" agemin="-1" name="Físico-Motora S2" handicap="2" />
                <AGEGROUP agegroupid="1326" agemax="-1" agemin="-1" name="Físico-Motora S3" handicap="3" />
                <AGEGROUP agegroupid="1327" agemax="-1" agemin="-1" name="Físico-Motora S4" handicap="4" />
                <AGEGROUP agegroupid="1328" agemax="-1" agemin="-1" name="Físico-Motora S5" handicap="5" />
                <AGEGROUP agegroupid="1329" agemax="-1" agemin="-1" name="Físico-Motora S6" handicap="6">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1330" agemax="-1" agemin="-1" name="Físico-Motora S7" handicap="7">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4148" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1331" agemax="-1" agemin="-1" name="Físico-Motora S8" handicap="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4136" />
                    <RANKING order="2" place="2" resultid="4124" />
                    <RANKING order="3" place="3" resultid="3982" />
                    <RANKING order="4" place="4" resultid="3953" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1332" agemax="-1" agemin="-1" name="Físico-Motora S9" handicap="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4113" />
                    <RANKING order="2" place="2" resultid="3880" />
                    <RANKING order="3" place="-1" resultid="3862" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1333" agemax="-1" agemin="-1" name="Físico-Motora S10" handicap="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3890" />
                    <RANKING order="2" place="2" resultid="3942" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1334" agemax="-1" agemin="-1" name="Visual S11" handicap="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4070" />
                    <RANKING order="2" place="2" resultid="4175" />
                    <RANKING order="3" place="-1" resultid="4074" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1335" agemax="-1" agemin="-1" name="Visual S12" handicap="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1336" agemax="-1" agemin="-1" name="Visual S13" handicap="13" />
                <AGEGROUP agegroupid="1337" agemax="-1" agemin="-1" name="Intelectual S14" handicap="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4047" />
                    <RANKING order="2" place="2" resultid="4107" />
                    <RANKING order="3" place="3" resultid="3930" />
                    <RANKING order="4" place="-1" resultid="4179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1338" agemax="-1" agemin="-1" name="Intelectual S18 (TEA)" handicap="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4054" />
                    <RANKING order="2" place="2" resultid="4079" />
                    <RANKING order="3" place="3" resultid="4013" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1339" agemax="-1" agemin="-1" name="Intelectual S21 (SD)" handicap="21">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4156" />
                    <RANKING order="2" place="2" resultid="3977" />
                    <RANKING order="3" place="3" resultid="3957" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4253" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="4254" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="4255" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="4256" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="4257" number="5" order="5" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1764" />
                <TIMESTANDARDREF timestandardlistid="1772" />
                <TIMESTANDARDREF timestandardlistid="1778" />
                <TIMESTANDARDREF timestandardlistid="1784" />
                <TIMESTANDARDREF timestandardlistid="1790" />
                <TIMESTANDARDREF timestandardlistid="1796" />
                <TIMESTANDARDREF timestandardlistid="1802" />
                <TIMESTANDARDREF timestandardlistid="1808" />
                <TIMESTANDARDREF timestandardlistid="1814" />
                <TIMESTANDARDREF timestandardlistid="1820" />
                <TIMESTANDARDREF timestandardlistid="1826" />
                <TIMESTANDARDREF timestandardlistid="1832" />
                <TIMESTANDARDREF timestandardlistid="1838" />
                <TIMESTANDARDREF timestandardlistid="1844" />
                <TIMESTANDARDREF timestandardlistid="1850" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1114" gender="F" number="26" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3163" agemax="-1" agemin="-1" name="DF">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4270" />
                    <RANKING order="2" place="2" resultid="4272" />
                    <RANKING order="3" place="-1" resultid="4271" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3164" agemax="-1" agemin="-1" name="DV">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4270" />
                    <RANKING order="2" place="2" resultid="4272" />
                    <RANKING order="3" place="-1" resultid="4271" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3165" agemax="-1" agemin="-1" name="DI">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4270" />
                    <RANKING order="2" place="2" resultid="4272" />
                    <RANKING order="3" place="-1" resultid="4271" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3166" agemax="-1" agemin="-1" name="SD">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4270" />
                    <RANKING order="2" place="2" resultid="4272" />
                    <RANKING order="3" place="-1" resultid="4271" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3167" agemax="-1" agemin="-1" name="TEA">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4270" />
                    <RANKING order="2" place="2" resultid="4272" />
                    <RANKING order="3" place="-1" resultid="4271" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4269" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1766" />
                <TIMESTANDARDREF timestandardlistid="1774" />
                <TIMESTANDARDREF timestandardlistid="1780" />
                <TIMESTANDARDREF timestandardlistid="1786" />
                <TIMESTANDARDREF timestandardlistid="1792" />
                <TIMESTANDARDREF timestandardlistid="1798" />
                <TIMESTANDARDREF timestandardlistid="1804" />
                <TIMESTANDARDREF timestandardlistid="1810" />
                <TIMESTANDARDREF timestandardlistid="1816" />
                <TIMESTANDARDREF timestandardlistid="1822" />
                <TIMESTANDARDREF timestandardlistid="1828" />
                <TIMESTANDARDREF timestandardlistid="1834" />
                <TIMESTANDARDREF timestandardlistid="1840" />
                <TIMESTANDARDREF timestandardlistid="1846" />
                <TIMESTANDARDREF timestandardlistid="1852" />
              </TIMESTANDARDREFS>
            </EVENT>
            <EVENT eventid="1116" gender="M" number="27" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="3168" agemax="-1" agemin="-1" name="DF">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4278" />
                    <RANKING order="2" place="2" resultid="4277" />
                    <RANKING order="3" place="3" resultid="4275" />
                    <RANKING order="4" place="-1" resultid="4276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3169" agemax="-1" agemin="-1" name="DV">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4278" />
                    <RANKING order="2" place="2" resultid="4277" />
                    <RANKING order="3" place="3" resultid="4275" />
                    <RANKING order="4" place="-1" resultid="4276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3170" agemax="-1" agemin="-1" name="DI">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4278" />
                    <RANKING order="2" place="2" resultid="4277" />
                    <RANKING order="3" place="3" resultid="4275" />
                    <RANKING order="4" place="-1" resultid="4276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3171" agemax="-1" agemin="-1" name="SD">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4278" />
                    <RANKING order="2" place="2" resultid="4277" />
                    <RANKING order="3" place="3" resultid="4275" />
                    <RANKING order="4" place="-1" resultid="4276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="3172" agemax="-1" agemin="-1" name="TEA">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4278" />
                    <RANKING order="2" place="2" resultid="4277" />
                    <RANKING order="3" place="3" resultid="4275" />
                    <RANKING order="4" place="-1" resultid="4276" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="4274" number="1" order="1" status="OFFICIAL" />
              </HEATS>
              <TIMESTANDARDREFS>
                <TIMESTANDARDREF timestandardlistid="1764" />
                <TIMESTANDARDREF timestandardlistid="1772" />
                <TIMESTANDARDREF timestandardlistid="1778" />
                <TIMESTANDARDREF timestandardlistid="1784" />
                <TIMESTANDARDREF timestandardlistid="1790" />
                <TIMESTANDARDREF timestandardlistid="1796" />
                <TIMESTANDARDREF timestandardlistid="1802" />
                <TIMESTANDARDREF timestandardlistid="1808" />
                <TIMESTANDARDREF timestandardlistid="1814" />
                <TIMESTANDARDREF timestandardlistid="1820" />
                <TIMESTANDARDREF timestandardlistid="1826" />
                <TIMESTANDARDREF timestandardlistid="1832" />
                <TIMESTANDARDREF timestandardlistid="1838" />
                <TIMESTANDARDREF timestandardlistid="1844" />
                <TIMESTANDARDREF timestandardlistid="1850" />
              </TIMESTANDARDREFS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="1488" nation="BRA" region="PR" clubid="4110" name="Seleção de Maringá" shortname="Maringá">
          <ATHLETES>
            <ATHLETE firstname="Matheus" lastname="Junio Brambilla" birthdate="2004-10-07" gender="M" nation="BRA" athleteid="4147">
              <HANDICAP exception="DF" free="7" />
              <RESULTS>
                <RESULT eventid="1111" points="201" swimtime="00:01:16.53" resultid="4148" heatid="4256" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="283" swimtime="00:00:33.12" resultid="4149" heatid="4228" lane="3" />
                <RESULT eventid="1098" points="252" swimtime="00:00:31.89" resultid="4150" heatid="4241" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Gomes Da Silva" birthdate="2000-06-09" gender="M" nation="BRA" athleteid="4123">
              <HANDICAP exception="DF" free="8" />
              <RESULTS>
                <RESULT eventid="1111" points="158" swimtime="00:01:22.90" resultid="4124" heatid="4253" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="96" swimtime="00:00:48.19" resultid="4125" heatid="4220" lane="5" />
                <RESULT eventid="1098" points="154" swimtime="00:00:37.61" resultid="4126" heatid="4240" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Sanches Da Silva Ghelere" birthdate="2008-08-06" gender="F" nation="BRA" athleteid="4131">
              <HANDICAP exception="DI" free="14" />
              <RESULTS>
                <RESULT eventid="1100" points="369" swimtime="00:01:15.31" resultid="4132" heatid="4244" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="444" swimtime="00:01:05.86" resultid="4133" heatid="4251" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="462" swimtime="00:00:29.65" resultid="4134" heatid="4234" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jonathan" lastname="Marcos Barros Drews" birthdate="1990-10-26" gender="M" nation="BRA" athleteid="4127">
              <HANDICAP exception="TEA" breast="18" free="18" />
              <RESULTS>
                <RESULT eventid="1081" status="DNS" swimtime="00:00:00.00" resultid="4128" heatid="4231" lane="3" />
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="4129" heatid="4239" lane="4" />
                <RESULT eventid="1107" status="DNS" swimtime="00:00:00.00" resultid="4130" heatid="4250" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Felipe Sakaguti" birthdate="2007-06-22" gender="M" nation="BRA" athleteid="4155">
              <HANDICAP exception="SD" free="21" />
              <RESULTS>
                <RESULT eventid="1111" points="69" swimtime="00:01:49.12" resultid="4156" heatid="4257" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="66" swimtime="00:00:54.45" resultid="4157" heatid="4221" lane="4" />
                <RESULT eventid="1098" points="86" swimtime="00:00:45.59" resultid="4158" heatid="4242" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Pauloski Murante" birthdate="1997-06-06" gender="M" nation="BRA" athleteid="4135">
              <HANDICAP exception="DF" breast="7" free="8" />
              <RESULTS>
                <RESULT eventid="1111" points="260" swimtime="00:01:10.25" resultid="4136" heatid="4254" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1070" points="176" swimtime="00:01:38.62" resultid="4137" heatid="4224" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="262" swimtime="00:00:31.50" resultid="4138" heatid="4240" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Lopes Ferreira" birthdate="2008-12-03" gender="F" nation="BRA" athleteid="4163">
              <HANDICAP exception="DF" breast="9" free="10" medley="10" />
              <RESULTS>
                <RESULT eventid="1079" points="181" swimtime="00:01:36.92" resultid="4164" heatid="4229" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="85" swimtime="00:00:55.37" resultid="4165" heatid="4226" lane="4" />
                <RESULT eventid="1096" status="DSQ" swimtime="00:00:38.67" resultid="4166" heatid="4235" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Henrique Vieira Góes" birthdate="2008-10-26" gender="M" nation="BRA" athleteid="4111">
              <HANDICAP exception="DF" breast="8" free="9" />
              <RESULTS>
                <RESULT eventid="1102" points="194" swimtime="00:01:22.53" resultid="4112" heatid="4245" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="271" swimtime="00:01:09.29" resultid="4113" heatid="4256" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1070" points="227" swimtime="00:01:30.52" resultid="4114" heatid="4224" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Débora" lastname="Borges Carneiro" birthdate="1998-05-07" gender="F" nation="BRA" athleteid="4119">
              <HANDICAP exception="DI" breast="14" free="14" />
              <RESULTS>
                <RESULT eventid="1068" status="WDR" swimtime="00:00:00.00" resultid="4120" />
                <RESULT eventid="1075" status="WDR" swimtime="00:00:00.00" resultid="4121" />
                <RESULT eventid="1096" status="WDR" swimtime="00:00:00.00" resultid="4122" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Roslaine" lastname="Da Silva Volpato" birthdate="1975-10-18" gender="F" nation="BRA" athleteid="4159">
              <HANDICAP exception="DF" free="6" />
              <RESULTS>
                <RESULT eventid="1109" points="192" swimtime="00:01:27.01" resultid="4160" heatid="4252" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="114" swimtime="00:00:50.14" resultid="4161" heatid="4225" lane="4" />
                <RESULT eventid="1096" points="100" swimtime="00:00:49.26" resultid="4162" heatid="4236" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Isabel Henriques" birthdate="2007-09-05" gender="F" nation="BRA" athleteid="4143">
              <HANDICAP exception="TEA" free="18" />
              <RESULTS>
                <RESULT eventid="1079" points="87" swimtime="00:02:03.47" resultid="4144" heatid="4229" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1109" points="128" swimtime="00:01:39.67" resultid="4145" heatid="4252" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="135" swimtime="00:00:44.61" resultid="4146" heatid="4235" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Da Silva Garcia Cateburcio" birthdate="2004-01-18" gender="F" nation="BRA" athleteid="4151">
              <HANDICAP exception="DF" free="8" />
              <RESULTS>
                <RESULT eventid="1109" points="58" swimtime="00:02:09.13" resultid="4152" heatid="4251" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" points="36" swimtime="00:01:16.07" resultid="4153" heatid="4216" lane="5" />
                <RESULT eventid="1096" points="71" swimtime="00:00:55.20" resultid="4154" heatid="4234" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Borges Carneiro" birthdate="1998-05-07" gender="F" nation="BRA" athleteid="4115">
              <HANDICAP exception="DI" breast="14" free="14" />
              <RESULTS>
                <RESULT eventid="1079" status="WDR" swimtime="00:00:00.00" resultid="4116" />
                <RESULT eventid="1068" status="WDR" swimtime="00:00:00.00" resultid="4117" />
                <RESULT eventid="1105" status="WDR" swimtime="00:00:00.00" resultid="4118" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Aparecida Pedro Souza" birthdate="2005-08-19" gender="F" nation="BRA" athleteid="4139">
              <HANDICAP exception="DI" free="14" />
              <RESULTS>
                <RESULT eventid="1109" points="46" swimtime="00:02:19.99" resultid="4140" heatid="4251" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="34" swimtime="00:01:15.05" resultid="4141" heatid="4226" lane="5" />
                <RESULT eventid="1096" points="43" swimtime="00:01:05.01" resultid="4142" heatid="4235" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="MARINGÁ &quot;A&quot;">
              <RESULTS>
                <RESULT eventid="1086" points="243" swimtime="00:02:11.08" resultid="4266" heatid="4263" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                    <SPLIT distance="100" swimtime="00:01:09.28" />
                    <SPLIT distance="150" swimtime="00:01:40.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4111" number="1" />
                    <RELAYPOSITION athleteid="4123" number="2" />
                    <RELAYPOSITION athleteid="4147" number="3" />
                    <RELAYPOSITION athleteid="4135" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1116" points="198" swimtime="00:02:33.89" resultid="4278" heatid="4274" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.41" />
                    <SPLIT distance="100" swimtime="00:01:31.05" />
                    <SPLIT distance="150" swimtime="00:02:03.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4123" number="1" />
                    <RELAYPOSITION athleteid="4111" number="2" />
                    <RELAYPOSITION athleteid="4147" number="3" />
                    <RELAYPOSITION athleteid="4135" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="MARINGÁ &quot;A&quot;">
              <RESULTS>
                <RESULT eventid="1084" status="WDR" swimtime="00:00:00.00" resultid="4261" heatid="4259" lane="3">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4115" number="1" />
                    <RELAYPOSITION athleteid="4119" number="2" />
                    <RELAYPOSITION athleteid="4131" number="3" />
                    <RELAYPOSITION athleteid="4139" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1114" status="WDR" swimtime="00:00:00.00" resultid="4271" heatid="4269" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4115" number="1" />
                    <RELAYPOSITION athleteid="4119" number="2" />
                    <RELAYPOSITION athleteid="4131" number="3" />
                    <RELAYPOSITION athleteid="4139" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="18108" nation="BRA" region="PR" clubid="3856" name="Seleção de Astorga" shortname="Astorga">
          <ATHLETES>
            <ATHLETE firstname="Jonatan" lastname="Rafael Nerys" birthdate="1985-05-13" gender="M" nation="BRA" athleteid="3861">
              <HANDICAP exception="DF" free="9" />
              <RESULTS>
                <RESULT eventid="1111" status="DNS" swimtime="00:00:00.00" resultid="3862" heatid="4256" lane="4" />
                <RESULT eventid="1066" status="DNS" swimtime="00:00:00.00" resultid="3863" heatid="4219" lane="2" />
                <RESULT eventid="1098" points="62" swimtime="00:00:50.75" resultid="3864" heatid="4238" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emerson" lastname="Moizes Ribeiro" birthdate="1986-10-16" gender="M" nation="BRA" athleteid="3857">
              <HANDICAP exception="DF" breast="6" free="6" />
              <RESULTS>
                <RESULT eventid="1066" points="24" swimtime="00:01:15.69" resultid="3858" heatid="4218" lane="2" />
                <RESULT eventid="1098" points="44" swimtime="00:00:56.94" resultid="3859" heatid="4242" lane="3" />
                <RESULT eventid="1107" status="DNS" swimtime="00:00:00.00" resultid="3860" heatid="4250" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1490" nation="BRA" region="PR" clubid="4167" name="Seleção de Ponta Grossa" shortname="Ponta Grossa">
          <ATHLETES>
            <ATHLETE firstname="Renan" lastname="André Araújo Cruz" birthdate="1993-10-02" gender="M" nation="BRA" athleteid="4168">
              <HANDICAP exception="DF" breast="7" free="8" medley="8" />
              <RESULTS>
                <RESULT eventid="1081" points="101" swimtime="00:01:43.62" resultid="4169" heatid="4231" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="108" swimtime="00:00:46.41" resultid="4170" heatid="4218" lane="3" />
                <RESULT eventid="1098" points="102" swimtime="00:00:43.13" resultid="4171" heatid="4241" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18116" nation="BRA" region="PR" clubid="4177" name="Seleção de Sertanópolis" shortname="Sertanópolis">
          <ATHLETES>
            <ATHLETE firstname="Renan" lastname="Soares De Freitas" birthdate="1997-10-14" gender="M" nation="BRA" athleteid="4178">
              <HANDICAP exception="DI" free="14" />
              <RESULTS>
                <RESULT eventid="1111" status="DSQ" swimtime="00:00:00.00" resultid="4179" heatid="4255" lane="1" />
                <RESULT eventid="1066" status="DSQ" swimtime="00:01:04.00" resultid="4180" heatid="4219" lane="3" />
                <RESULT eventid="1098" points="71" swimtime="00:00:48.47" resultid="4181" heatid="4237" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="689" nation="BRA" region="PR" clubid="3893" name="Seleção de Cascavel" shortname="Cascavel">
          <ATHLETES>
            <ATHLETE firstname="Carlos" lastname="Augusto Alencar De Carvalho" birthdate="2002-10-16" gender="M" nation="BRA" athleteid="3898">
              <HANDICAP exception="DF" breast="3" free="4" />
              <RESULTS>
                <RESULT eventid="1066" points="16" swimtime="00:01:26.62" resultid="3899" heatid="4219" lane="6" />
                <RESULT eventid="1098" points="29" swimtime="00:01:04.95" resultid="3900" heatid="4240" lane="2" />
                <RESULT eventid="1107" points="25" swimtime="00:01:24.33" resultid="3901" heatid="4250" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Paulo Kall" birthdate="2003-06-27" gender="M" nation="BRA" athleteid="3917">
              <HANDICAP exception="DF" free="10" />
              <RESULTS>
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="3918" heatid="4240" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Pereira Gonçalves" birthdate="2006-08-19" gender="F" nation="BRA" athleteid="3894">
              <HANDICAP exception="DF" breast="9" free="9" />
              <RESULTS>
                <RESULT eventid="1068" points="89" swimtime="00:02:19.25" resultid="3895" heatid="4223" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="63" swimtime="00:01:01.05" resultid="3896" heatid="4225" lane="3" />
                <RESULT eventid="1105" points="92" swimtime="00:01:02.71" resultid="3897" heatid="4246" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Paulo Ribeiro Dos Santos" birthdate="2007-06-22" gender="M" nation="BRA" athleteid="3913">
              <HANDICAP exception="DF" />
              <RESULTS>
                <RESULT eventid="1098" status="WDR" swimtime="00:00:00.00" resultid="3914" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Bento Da Silva" birthdate="1991-10-01" gender="M" nation="BRA" athleteid="3909">
              <HANDICAP exception="DV" breast="11" free="11" />
              <RESULTS>
                <RESULT eventid="1070" status="DNS" swimtime="00:00:00.00" resultid="3910" heatid="4224" lane="1" />
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="3911" heatid="4243" lane="1" />
                <RESULT eventid="1107" status="DNS" swimtime="00:00:00.00" resultid="3912" heatid="4248" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dany" lastname="Joel Hernandez Mujica" birthdate="2004-02-20" gender="M" nation="BRA" athleteid="3906">
              <HANDICAP exception="DV" />
              <RESULTS>
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="3907" heatid="4238" lane="1" />
                <RESULT eventid="1107" status="DNS" swimtime="00:00:00.00" resultid="3908" heatid="4249" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Gabriel Canan Phillpesen" birthdate="2007-03-29" gender="M" nation="BRA" athleteid="3915">
              <HANDICAP exception="TEA" free="18" />
              <RESULTS>
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="3916" heatid="4239" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cleoni" lastname="Vilas Boas Da Silva" birthdate="1985-11-12" gender="M" nation="BRA" athleteid="3902">
              <HANDICAP exception="DF" breast="7" free="7" />
              <RESULTS>
                <RESULT eventid="1070" points="39" swimtime="00:02:41.92" resultid="3903" heatid="4224" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="15" swimtime="00:01:20.92" resultid="3904" heatid="4241" lane="6" />
                <RESULT eventid="1107" points="36" swimtime="00:01:15.54" resultid="3905" heatid="4249" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18109" nation="BRA" region="PR" clubid="4085" name="Seleção de Mandaguari" shortname="Mandaguari">
          <ATHLETES>
            <ATHLETE firstname="Alessandro" lastname="Bula Balan" birthdate="1984-04-10" gender="M" nation="BRA" athleteid="4086">
              <HANDICAP exception="SD" free="21" />
              <RESULTS>
                <RESULT eventid="1077" points="43" swimtime="00:01:01.77" resultid="4087" heatid="4228" lane="5" />
                <RESULT eventid="1066" points="64" swimtime="00:00:55.23" resultid="4088" heatid="4221" lane="2" />
                <RESULT eventid="1098" points="59" swimtime="00:00:51.70" resultid="4089" heatid="4242" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jana" lastname="Beidoun" birthdate="1998-12-11" gender="F" nation="BRA" athleteid="4097">
              <HANDICAP exception="TEA" free="18" />
              <RESULTS>
                <RESULT eventid="1109" points="32" swimtime="00:02:36.71" resultid="4098" heatid="4251" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" points="38" swimtime="00:01:14.80" resultid="4099" heatid="4216" lane="2" />
                <RESULT eventid="1096" points="46" swimtime="00:01:03.99" resultid="4100" heatid="4235" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Murilo Fante" birthdate="2001-04-03" gender="M" nation="BRA" athleteid="4094">
              <HANDICAP exception="TEA" free="18" />
              <RESULTS>
                <RESULT eventid="1066" points="19" swimtime="00:01:22.51" resultid="4095" heatid="4220" lane="2" />
                <RESULT eventid="1098" points="41" swimtime="00:00:58.30" resultid="4096" heatid="4239" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mirian" lastname="Rose Garcia Gouvea" birthdate="1989-10-25" gender="F" nation="BRA" athleteid="4101">
              <HANDICAP exception="DI" free="14" />
              <RESULTS>
                <RESULT eventid="1100" points="258" swimtime="00:01:24.87" resultid="4102" heatid="4244" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="240" swimtime="00:01:28.29" resultid="4103" heatid="4229" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="317" swimtime="00:00:35.73" resultid="4104" heatid="4226" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emanuelle" lastname="Victória Sá De Araújo" birthdate="2007-03-24" gender="F" nation="BRA" athleteid="4090">
              <HANDICAP exception="DF" free="6" medley="6" />
              <RESULTS>
                <RESULT eventid="1079" points="89" swimtime="00:02:02.92" resultid="4091" heatid="4229" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="175" swimtime="00:03:17.05" resultid="4092" heatid="4213" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.67" />
                    <SPLIT distance="100" swimtime="00:01:33.20" />
                    <SPLIT distance="150" swimtime="00:02:24.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1088" points="99" swimtime="00:04:23.26" resultid="4093" heatid="4232" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.59" />
                    <SPLIT distance="100" swimtime="00:02:04.75" />
                    <SPLIT distance="150" swimtime="00:03:30.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="10975" nation="BRA" region="PR" clubid="3865" name="Seleção de Campo Largo" shortname="Campo Largo">
          <ATHLETES>
            <ATHLETE firstname="Jhonatan" lastname="Lechenski Estevam" birthdate="1992-07-15" gender="M" nation="BRA" athleteid="3866">
              <HANDICAP exception="DF" breast="9" free="9" medley="9" />
              <RESULTS>
                <RESULT eventid="1066" points="12" swimtime="00:01:35.14" resultid="3867" heatid="4219" lane="5" />
                <RESULT eventid="1098" points="46" swimtime="00:00:55.95" resultid="3868" heatid="4238" lane="5" />
                <RESULT eventid="1107" status="DSQ" swimtime="00:01:23.94" resultid="3869" heatid="4250" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Henrique Krupa" birthdate="2002-06-14" gender="M" nation="BRA" athleteid="3870">
              <HANDICAP exception="SD" breast="21" free="21" />
              <RESULTS>
                <RESULT eventid="1066" points="24" swimtime="00:01:16.36" resultid="3871" heatid="4222" lane="3" />
                <RESULT eventid="1098" points="32" swimtime="00:01:02.95" resultid="3872" heatid="4242" lane="2" />
                <RESULT eventid="1107" points="22" swimtime="00:01:27.79" resultid="3873" heatid="4249" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6462" nation="BRA" region="PR" clubid="4172" name="Seleção de São José dos Pinhais" shortname="São José dos Pinhais">
          <ATHLETES>
            <ATHLETE firstname="Juan" lastname="Marcelo Da Silva Santos" birthdate="2001-04-04" gender="M" nation="BRA" athleteid="4173">
              <HANDICAP exception="DV" breast="11" free="11" medley="11" />
              <RESULTS>
                <RESULT eventid="1081" status="DSQ" swimtime="00:02:26.05" resultid="4174" heatid="4230" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="63" swimtime="00:01:52.64" resultid="4175" heatid="4257" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="71" swimtime="00:00:48.57" resultid="4176" heatid="4243" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1492" nation="BRA" region="PR" clubid="3919" name="Seleção de Curitiba" shortname="Curitiba">
          <ATHLETES>
            <ATHLETE firstname="Adriano" lastname="Braune" birthdate="1998-11-23" gender="M" nation="BRA" athleteid="3920">
              <HANDICAP exception="DI" free="14" />
              <RESULTS>
                <RESULT eventid="1062" points="77" swimtime="00:03:53.11" resultid="3921" heatid="4215" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.19" />
                    <SPLIT distance="100" swimtime="00:01:43.12" />
                    <SPLIT distance="150" swimtime="00:02:47.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="49" swimtime="00:01:00.40" resultid="3922" heatid="4221" lane="5" />
                <RESULT eventid="1098" points="89" swimtime="00:00:45.04" resultid="3923" heatid="4237" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jéssica" lastname="Eloisa Pedroso" birthdate="1997-02-12" gender="F" nation="BRA" athleteid="3988">
              <HANDICAP exception="DI" breast="14" free="14" />
              <RESULTS>
                <RESULT eventid="1079" points="79" swimtime="00:02:07.47" resultid="3989" heatid="4229" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="77" swimtime="00:02:26.55" resultid="3990" heatid="4223" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" points="77" swimtime="00:00:59.29" resultid="3991" heatid="4216" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Lima Cardoso" birthdate="2000-06-12" gender="M" nation="BRA" athleteid="4069">
              <HANDICAP exception="DV" free="11" />
              <RESULTS>
                <RESULT eventid="1111" points="113" swimtime="00:01:32.51" resultid="4070" heatid="4257" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="84" swimtime="00:00:50.41" resultid="4071" heatid="4220" lane="1" />
                <RESULT eventid="1098" points="149" swimtime="00:00:37.99" resultid="4072" heatid="4243" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorena" lastname="Isabel Bylnoski" birthdate="1984-07-13" gender="F" nation="BRA" athleteid="4008">
              <HANDICAP exception="DF" breast="9" free="9" />
              <RESULTS>
                <RESULT eventid="1064" points="22" swimtime="00:01:29.43" resultid="4009" heatid="4216" lane="4" />
                <RESULT eventid="1096" points="36" swimtime="00:01:09.01" resultid="4010" heatid="4236" lane="5" />
                <RESULT eventid="1105" points="22" swimtime="00:01:40.30" resultid="4011" heatid="4246" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Gustavo Lopes Nonato" birthdate="2004-07-26" gender="M" nation="BRA" athleteid="4019">
              <HANDICAP exception="SD" free="21" />
              <RESULTS>
                <RESULT eventid="1066" points="20" swimtime="00:01:21.30" resultid="4020" heatid="4222" lane="6" />
                <RESULT eventid="1098" points="14" swimtime="00:01:23.63" resultid="4021" heatid="4242" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Lubian" birthdate="2007-12-14" gender="F" nation="BRA" athleteid="3936">
              <HANDICAP exception="DF" free="6" />
              <RESULTS>
                <RESULT eventid="1109" points="38" swimtime="00:02:28.59" resultid="3937" heatid="4252" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="39" swimtime="00:01:11.39" resultid="3938" heatid="4225" lane="2" />
                <RESULT eventid="1096" points="40" swimtime="00:01:06.57" resultid="3939" heatid="4235" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leandro" lastname="Vosne Da Rosa" birthdate="1987-06-26" gender="M" nation="BRA" athleteid="4004">
              <HANDICAP exception="DV" breast="12" free="12" />
              <RESULTS>
                <RESULT eventid="1066" status="DNS" swimtime="00:00:00.00" resultid="4005" heatid="4221" lane="1" />
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="4006" heatid="4241" lane="1" />
                <RESULT eventid="1107" status="DNS" swimtime="00:00:00.00" resultid="4007" heatid="4249" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Miguel Dos Santos Ferreira" birthdate="2005-07-26" gender="M" nation="BRA" athleteid="3932">
              <HANDICAP exception="DF" free="6" />
              <RESULTS>
                <RESULT eventid="1111" points="112" swimtime="00:01:32.78" resultid="3933" heatid="4256" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1062" points="133" swimtime="00:03:14.32" resultid="3934" heatid="4214" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.15" />
                    <SPLIT distance="100" swimtime="00:01:34.16" />
                    <SPLIT distance="150" swimtime="00:02:24.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="98" swimtime="00:00:47.15" resultid="3935" heatid="4227" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Flaviano" lastname="Fagundes" birthdate="1992-12-26" gender="M" nation="BRA" athleteid="3952">
              <HANDICAP exception="DF" breast="7" free="8" medley="8" />
              <RESULTS>
                <RESULT eventid="1111" points="65" swimtime="00:01:51.43" resultid="3953" heatid="4253" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="37" swimtime="00:01:06.34" resultid="3954" heatid="4220" lane="6" />
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="3955" heatid="4241" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Erick" lastname="Campos Arruda" birthdate="2004-05-17" gender="M" nation="BRA" athleteid="3948">
              <HANDICAP exception="DF" breast="5" free="6" />
              <RESULTS>
                <RESULT eventid="1066" points="18" swimtime="00:01:24.18" resultid="3949" heatid="4218" lane="4" />
                <RESULT eventid="1098" points="49" swimtime="00:00:54.81" resultid="3950" heatid="4238" lane="4" />
                <RESULT eventid="1107" status="DNS" swimtime="00:00:00.00" resultid="3951" heatid="4248" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovani" lastname="Mayer" birthdate="1972-10-28" gender="M" nation="BRA" athleteid="3968">
              <HANDICAP exception="DV" free="12" />
              <RESULTS>
                <RESULT eventid="1111" points="69" swimtime="00:01:49.11" resultid="3969" heatid="4256" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1062" points="69" swimtime="00:04:01.30" resultid="3970" heatid="4215" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.36" />
                    <SPLIT distance="100" swimtime="00:01:53.38" />
                    <SPLIT distance="150" swimtime="00:02:58.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="29" swimtime="00:01:11.79" resultid="3971" heatid="4222" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Renato" lastname="Lucas Da Cunha Constantino" birthdate="2005-09-15" gender="M" nation="BRA" athleteid="4049">
              <HANDICAP exception="DI" breast="14" free="14" />
              <RESULTS>
                <RESULT eventid="1066" status="DSQ" swimtime="00:00:50.82" resultid="4050" heatid="4221" lane="6" />
                <RESULT eventid="1098" points="132" swimtime="00:00:39.55" resultid="4051" heatid="4237" lane="6" />
                <RESULT eventid="1107" status="DSQ" swimtime="00:01:08.91" resultid="4052" heatid="4248" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelo" lastname="De França" birthdate="1975-12-10" gender="M" nation="BRA" athleteid="4026">
              <HANDICAP exception="DF" breast="6" free="7" />
              <RESULTS>
                <RESULT eventid="1062" points="35" swimtime="00:05:02.78" resultid="4027" heatid="4215" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.65" />
                    <SPLIT distance="100" swimtime="00:02:22.97" />
                    <SPLIT distance="150" swimtime="00:03:47.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="28" swimtime="00:01:12.19" resultid="4028" heatid="4222" lane="2" />
                <RESULT eventid="1107" points="13" swimtime="00:01:44.40" resultid="4029" heatid="4248" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anderson" lastname="Andrade Leal" birthdate="1987-08-06" gender="M" nation="BRA" athleteid="3928">
              <HANDICAP exception="DI" free="14" />
              <RESULTS>
                <RESULT eventid="1081" points="66" swimtime="00:01:59.45" resultid="3929" heatid="4231" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="123" swimtime="00:01:30.00" resultid="3930" heatid="4254" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1062" points="91" swimtime="00:03:40.29" resultid="3931" heatid="4215" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.79" />
                    <SPLIT distance="100" swimtime="00:01:35.84" />
                    <SPLIT distance="150" swimtime="00:02:34.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Marina Dantas Novaes" birthdate="1984-09-04" gender="F" nation="BRA" athleteid="4015">
              <HANDICAP exception="DF" />
              <RESULTS>
                <RESULT eventid="1075" status="WDR" swimtime="00:00:00.00" resultid="4016" />
                <RESULT eventid="1064" status="WDR" swimtime="00:00:00.00" resultid="4017" />
                <RESULT eventid="1096" status="WDR" swimtime="00:00:00.00" resultid="4018" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Da Silva Fabris" birthdate="1993-04-21" gender="F" nation="BRA" athleteid="3964">
              <HANDICAP exception="DI" free="14" />
              <RESULTS>
                <RESULT eventid="1109" points="135" swimtime="00:01:37.76" resultid="3965" heatid="4251" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="145" swimtime="00:03:29.65" resultid="3966" heatid="4213" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.22" />
                    <SPLIT distance="100" swimtime="00:01:46.05" />
                    <SPLIT distance="150" swimtime="00:02:41.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="85" swimtime="00:00:55.30" resultid="3967" heatid="4226" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicollas" lastname="Henrique Kaguimoto Ferreira" birthdate="1994-05-23" gender="M" nation="BRA" athleteid="4045">
              <HANDICAP exception="DI" free="14" />
              <RESULTS>
                <RESULT eventid="1102" points="131" swimtime="00:01:34.03" resultid="4046" heatid="4245" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="246" swimtime="00:01:11.55" resultid="4047" heatid="4254" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="158" swimtime="00:00:40.15" resultid="4048" heatid="4228" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Damásio Nascimento" birthdate="2008-08-25" gender="F" nation="BRA" athleteid="3984">
              <HANDICAP exception="DF" breast="5" free="7" />
              <RESULTS>
                <RESULT eventid="1068" status="DSQ" swimtime="00:05:41.32" resultid="3985" heatid="4223" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:02:40.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="28" swimtime="00:01:14.89" resultid="3986" heatid="4236" lane="3" />
                <RESULT eventid="1105" status="DSQ" swimtime="00:02:51.51" resultid="3987" heatid="4246" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tisbe" lastname="De Souza Andrade" birthdate="1998-07-21" gender="F" nation="BRA" athleteid="4065">
              <HANDICAP exception="DF" free="5" />
              <RESULTS>
                <RESULT eventid="1075" points="46" swimtime="00:01:07.97" resultid="4066" heatid="4226" lane="2" />
                <RESULT eventid="1064" points="81" swimtime="00:00:58.31" resultid="4067" heatid="4217" lane="2" />
                <RESULT eventid="1096" points="57" swimtime="00:00:59.52" resultid="4068" heatid="4234" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Felipe De Souza" birthdate="1994-04-27" gender="M" nation="BRA" athleteid="4022">
              <HANDICAP exception="DF" breast="8" free="9" />
              <RESULTS>
                <RESULT eventid="1081" points="152" swimtime="00:01:30.53" resultid="4023" heatid="4231" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1070" points="170" swimtime="00:01:39.78" resultid="4024" heatid="4224" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="174" swimtime="00:00:36.08" resultid="4025" heatid="4238" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Altamir" lastname="Pereira" birthdate="1958-03-13" gender="M" nation="BRA" athleteid="3924">
              <HANDICAP exception="DF" breast="8" free="9" />
              <RESULTS>
                <RESULT eventid="1066" status="DSQ" swimtime="00:01:34.93" resultid="3925" heatid="4219" lane="1" />
                <RESULT eventid="1098" points="29" swimtime="00:01:05.38" resultid="3926" heatid="4238" lane="2" />
                <RESULT eventid="1107" status="DSQ" swimtime="00:01:42.89" resultid="3927" heatid="4247" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Delgado Carvalho" birthdate="2007-09-03" gender="M" nation="BRA" athleteid="4042">
              <HANDICAP exception="TEA" breast="18" free="18" />
              <RESULTS>
                <RESULT eventid="1098" points="44" swimtime="00:00:57.06" resultid="4043" heatid="4239" lane="6" />
                <RESULT eventid="1107" points="83" swimtime="00:00:57.10" resultid="4044" heatid="4250" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dayane" lastname="Esther Pinheiro" birthdate="1996-04-12" gender="F" nation="BRA" athleteid="3944">
              <HANDICAP exception="DV" free="12" />
              <RESULTS>
                <RESULT eventid="1075" points="19" swimtime="00:01:30.03" resultid="3945" heatid="4226" lane="1" />
                <RESULT eventid="1064" points="18" swimtime="00:01:36.22" resultid="3946" heatid="4217" lane="1" />
                <RESULT eventid="1096" points="38" swimtime="00:01:07.97" resultid="3947" heatid="4236" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Felipe Domingues Masena" birthdate="2004-11-29" gender="M" nation="BRA" athleteid="3980">
              <HANDICAP exception="DF" free="8" />
              <RESULTS>
                <RESULT eventid="1081" points="56" swimtime="00:02:05.84" resultid="3981" heatid="4231" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="73" swimtime="00:01:46.81" resultid="3982" heatid="4253" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="84" swimtime="00:00:45.86" resultid="3983" heatid="4240" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Talita" lastname="Aparecida Cuceravai" birthdate="1986-09-05" gender="F" nation="BRA" athleteid="4061">
              <HANDICAP exception="DI" breast="14" free="14" />
              <RESULTS>
                <RESULT eventid="1109" points="38" swimtime="00:02:29.04" resultid="4062" heatid="4251" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="61" swimtime="00:00:57.96" resultid="4063" heatid="4234" lane="4" />
                <RESULT eventid="1105" points="22" swimtime="00:01:40.70" resultid="4064" heatid="4246" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ketlyn" lastname="Padilha Veitex" birthdate="2001-03-04" gender="F" nation="BRA" athleteid="4000">
              <HANDICAP exception="SD" free="21" />
              <RESULTS>
                <RESULT eventid="1109" points="47" swimtime="00:02:19.22" resultid="4001" heatid="4252" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" points="33" swimtime="00:01:18.09" resultid="4002" heatid="4217" lane="5" />
                <RESULT eventid="1096" status="DSQ" swimtime="00:00:57.96" resultid="4003" heatid="4235" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Melissa" lastname="Karla De Oliveira" birthdate="1980-07-07" gender="F" nation="BRA" athleteid="4038">
              <HANDICAP exception="DI" free="14" />
              <RESULTS>
                <RESULT eventid="1079" points="21" swimtime="00:03:16.81" resultid="4039" heatid="4229" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:34.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="24" swimtime="00:06:20.81" resultid="4040" heatid="4213" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:22.56" />
                    <SPLIT distance="100" swimtime="00:02:55.78" />
                    <SPLIT distance="150" swimtime="00:04:37.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" status="DNS" swimtime="00:00:00.00" resultid="4041" heatid="4217" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cleverson" lastname="Ribeiro Dos Santos" birthdate="1996-11-12" gender="M" nation="BRA" athleteid="3940">
              <HANDICAP exception="DF" free="10" />
              <RESULTS>
                <RESULT eventid="1081" points="178" swimtime="00:01:25.81" resultid="3941" heatid="4231" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1111" points="259" swimtime="00:01:10.34" resultid="3942" heatid="4255" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="240" swimtime="00:00:32.40" resultid="3943" heatid="4240" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Inacio Berti" birthdate="1991-08-20" gender="M" nation="BRA" athleteid="3960">
              <HANDICAP exception="SD" breast="21" free="21" />
              <RESULTS>
                <RESULT eventid="1081" points="15" swimtime="00:03:15.86" resultid="3961" heatid="4230" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:34.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1062" points="27" swimtime="00:05:28.30" resultid="3962" heatid="4215" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:15.86" />
                    <SPLIT distance="100" swimtime="00:02:37.69" />
                    <SPLIT distance="150" swimtime="00:04:02.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" status="DSQ" swimtime="00:01:37.97" resultid="3963" heatid="4249" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Romano Sartor" birthdate="1994-06-29" gender="F" nation="BRA" athleteid="3996">
              <HANDICAP exception="DI" breast="14" free="14" />
              <RESULTS>
                <RESULT eventid="1064" points="51" swimtime="00:01:07.66" resultid="3997" heatid="4217" lane="6" />
                <RESULT eventid="1096" points="135" swimtime="00:00:44.59" resultid="3998" heatid="4234" lane="2" />
                <RESULT eventid="1105" points="93" swimtime="00:01:02.43" resultid="3999" heatid="4246" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Dos Santos Ferreira" birthdate="1999-09-28" gender="M" nation="BRA" athleteid="3956">
              <HANDICAP exception="SD" free="21" />
              <RESULTS>
                <RESULT eventid="1111" points="35" swimtime="00:02:16.51" resultid="3957" heatid="4257" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="26" swimtime="00:01:13.02" resultid="3958" heatid="4228" lane="2" />
                <RESULT eventid="1098" points="42" swimtime="00:00:57.94" resultid="3959" heatid="4239" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrike" lastname="Furquim Barbosa" birthdate="2007-08-09" gender="M" nation="BRA" athleteid="3976">
              <HANDICAP exception="SD" free="21" />
              <RESULTS>
                <RESULT eventid="1111" points="37" swimtime="00:02:14.09" resultid="3977" heatid="4257" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1062" points="40" swimtime="00:04:50.32" resultid="3978" heatid="4215" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.57" />
                    <SPLIT distance="100" swimtime="00:02:12.60" />
                    <SPLIT distance="150" swimtime="00:03:32.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="28" swimtime="00:01:12.77" resultid="3979" heatid="4221" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Suzana" lastname="De Almeida Pinheiro" birthdate="1986-04-21" gender="F" nation="BRA" athleteid="4057">
              <HANDICAP exception="DF" breast="6" free="6" medley="6" />
              <RESULTS>
                <RESULT eventid="1109" points="63" swimtime="00:02:05.80" resultid="4058" heatid="4252" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" points="59" swimtime="00:01:04.51" resultid="4059" heatid="4216" lane="1" />
                <RESULT eventid="1096" points="83" swimtime="00:00:52.53" resultid="4060" heatid="4236" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luan" lastname="Neo São Marcos" birthdate="2002-05-01" gender="M" nation="BRA" athleteid="4012">
              <HANDICAP exception="TEA" free="18" />
              <RESULTS>
                <RESULT eventid="1111" points="81" swimtime="00:01:43.48" resultid="4013" heatid="4255" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="57" swimtime="00:00:57.23" resultid="4014" heatid="4220" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariana" lastname="Oliva" birthdate="1993-06-20" gender="F" nation="BRA" athleteid="4034">
              <HANDICAP exception="DF" free="7" />
              <RESULTS>
                <RESULT eventid="1109" points="49" swimtime="00:02:16.85" resultid="4035" heatid="4252" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" status="DSQ" swimtime="00:01:09.94" resultid="4036" heatid="4217" lane="4" />
                <RESULT eventid="1096" points="50" swimtime="00:01:02.13" resultid="4037" heatid="4236" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Manassés Da Silva De Oliveira" birthdate="2007-04-27" gender="M" nation="BRA" athleteid="3972">
              <HANDICAP exception="TEA" free="18" />
              <RESULTS>
                <RESULT eventid="1077" points="66" swimtime="00:00:53.63" resultid="3973" heatid="4227" lane="3" />
                <RESULT eventid="1066" points="93" swimtime="00:00:48.71" resultid="3974" heatid="4220" lane="3" />
                <RESULT eventid="1098" points="130" swimtime="00:00:39.72" resultid="3975" heatid="4237" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Saimon" lastname="Rodrigues Stang" birthdate="2008-02-23" gender="M" nation="BRA" athleteid="4053">
              <HANDICAP exception="TEA" breast="18" free="18" />
              <RESULTS>
                <RESULT eventid="1111" points="182" swimtime="00:01:19.04" resultid="4054" heatid="4255" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="137" swimtime="00:00:42.15" resultid="4055" heatid="4227" lane="4" />
                <RESULT eventid="1107" points="180" swimtime="00:00:44.16" resultid="4056" heatid="4250" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose" lastname="Carlos Mendonça" birthdate="1981-10-04" gender="M" nation="BRA" athleteid="3992">
              <HANDICAP exception="DF" breast="5" free="6" />
              <RESULTS>
                <RESULT eventid="1081" points="26" swimtime="00:02:43.09" resultid="3993" heatid="4230" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:17.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1062" points="52" swimtime="00:04:25.24" resultid="3994" heatid="4214" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.47" />
                    <SPLIT distance="100" swimtime="00:02:03.62" />
                    <SPLIT distance="150" swimtime="00:03:16.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="62" swimtime="00:01:02.87" resultid="3995" heatid="4248" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wagner" lastname="Bitencourt" birthdate="1986-01-13" gender="M" nation="BRA" athleteid="4073">
              <HANDICAP exception="DV" free="11" />
              <RESULTS>
                <RESULT eventid="1111" status="DNS" swimtime="00:00:00.00" resultid="4074" heatid="4257" lane="2" />
                <RESULT eventid="1062" status="DNS" swimtime="00:00:00.00" resultid="4075" heatid="4214" lane="1" />
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="4076" heatid="4243" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Isabel Kfuri Dos Santos" birthdate="2005-12-20" gender="F" nation="BRA" athleteid="4030">
              <HANDICAP exception="DF" />
              <RESULTS>
                <RESULT eventid="1100" status="DSQ" swimtime="00:00:00.00" resultid="4031" heatid="4244" lane="5" late="yes" />
                <RESULT eventid="1060" points="267" status="EXH" swimtime="00:02:51.27" resultid="4032" heatid="4213" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.59" />
                    <SPLIT distance="100" swimtime="00:01:21.30" />
                    <SPLIT distance="150" swimtime="00:02:06.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="203" status="EXH" swimtime="00:00:41.43" resultid="4033" heatid="4225" lane="5" late="yes" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBA &quot;A&quot;">
              <RESULTS>
                <RESULT eventid="1086" status="WDR" swimtime="00:00:00.00" resultid="4268" heatid="4263" lane="1">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3968" number="1" />
                    <RELAYPOSITION athleteid="4004" number="2" />
                    <RELAYPOSITION athleteid="4069" number="3" />
                    <RELAYPOSITION athleteid="4073" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1116" points="136" swimtime="00:02:54.10" resultid="4277" heatid="4274" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.23" />
                    <SPLIT distance="100" swimtime="00:01:39.03" />
                    <SPLIT distance="150" swimtime="00:02:14.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3980" number="1" />
                    <RELAYPOSITION athleteid="4022" number="2" />
                    <RELAYPOSITION athleteid="3940" number="3" />
                    <RELAYPOSITION athleteid="3932" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1086" points="133" swimtime="00:02:40.05" resultid="4267" heatid="4263" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.61" />
                    <SPLIT distance="100" swimtime="00:01:21.59" />
                    <SPLIT distance="150" swimtime="00:02:06.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4049" number="1" />
                    <RELAYPOSITION athleteid="3928" number="2" />
                    <RELAYPOSITION athleteid="3920" number="3" />
                    <RELAYPOSITION athleteid="4045" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1116" points="81" swimtime="00:03:26.87" resultid="4275" heatid="4274" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.46" />
                    <SPLIT distance="100" swimtime="00:02:04.49" />
                    <SPLIT distance="150" swimtime="00:02:42.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4049" number="1" />
                    <RELAYPOSITION athleteid="3928" number="2" />
                    <RELAYPOSITION athleteid="4045" number="3" />
                    <RELAYPOSITION athleteid="3920" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBA &quot;A&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1086" points="126" swimtime="00:02:42.78" resultid="4265" heatid="4263" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.42" />
                    <SPLIT distance="100" swimtime="00:01:23.13" />
                    <SPLIT distance="150" swimtime="00:02:06.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3940" number="1" />
                    <RELAYPOSITION athleteid="3992" number="2" />
                    <RELAYPOSITION athleteid="3980" number="3" />
                    <RELAYPOSITION athleteid="4022" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBA &quot;A&quot;">
              <RESULTS>
                <RESULT eventid="1084" points="104" swimtime="00:03:16.12" resultid="4260" heatid="4259" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.07" />
                    <SPLIT distance="100" swimtime="00:01:35.38" />
                    <SPLIT distance="150" swimtime="00:02:35.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3996" number="1" />
                    <RELAYPOSITION athleteid="3988" number="2" />
                    <RELAYPOSITION athleteid="4061" number="3" />
                    <RELAYPOSITION athleteid="3964" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1114" points="53" swimtime="00:04:32.25" resultid="4270" heatid="4269" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.94" />
                    <SPLIT distance="100" swimtime="00:02:50.37" />
                    <SPLIT distance="150" swimtime="00:03:47.01" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3996" number="1" />
                    <RELAYPOSITION athleteid="4061" number="2" />
                    <RELAYPOSITION athleteid="3964" number="3" />
                    <RELAYPOSITION athleteid="3988" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1084" points="43" swimtime="00:04:22.73" resultid="4262" heatid="4259" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.30" />
                    <SPLIT distance="100" swimtime="00:02:19.79" />
                    <SPLIT distance="150" swimtime="00:03:20.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3936" number="1" />
                    <RELAYPOSITION athleteid="4008" number="2" />
                    <RELAYPOSITION athleteid="4034" number="3" />
                    <RELAYPOSITION athleteid="4065" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1114" points="44" swimtime="00:04:48.31" resultid="4272" heatid="4269" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.52" />
                    <SPLIT distance="100" swimtime="00:02:41.38" />
                    <SPLIT distance="150" swimtime="00:03:57.23" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4065" number="1" />
                    <RELAYPOSITION athleteid="4008" number="2" />
                    <RELAYPOSITION athleteid="3936" number="3" />
                    <RELAYPOSITION athleteid="4057" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBA &quot;A&quot;">
              <RESULTS>
                <RESULT eventid="1073" points="36" swimtime="00:04:24.10" resultid="4280" heatid="4279" lane="3" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.60" />
                    <SPLIT distance="100" swimtime="00:02:11.91" />
                    <SPLIT distance="150" swimtime="00:03:33.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3944" number="1" />
                    <RELAYPOSITION athleteid="3976" number="2" />
                    <RELAYPOSITION athleteid="4038" number="3" />
                    <RELAYPOSITION athleteid="3952" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="18111" nation="BRA" region="PR" clubid="4105" name="Seleção de Marilândia do Sul" shortname="Marilândia do Sul">
          <ATHLETES>
            <ATHLETE firstname="Lucas" lastname="Gutierres" birthdate="1995-05-19" gender="M" nation="BRA" athleteid="4106">
              <HANDICAP exception="DI" free="14" />
              <RESULTS>
                <RESULT eventid="1111" points="140" swimtime="00:01:26.32" resultid="4107" heatid="4255" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="112" swimtime="00:00:45.82" resultid="4108" heatid="4219" lane="4" />
                <RESULT eventid="1098" points="140" swimtime="00:00:38.78" resultid="4109" heatid="4237" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1493" nation="BRA" region="PR" clubid="4077" name="Seleção de Londrina" shortname="Londrina">
          <ATHLETES>
            <ATHLETE firstname="Thiago" lastname="Stela Bornia" birthdate="1981-07-01" gender="M" nation="BRA" athleteid="4082">
              <HANDICAP exception="DV" breast="11" free="11" />
              <RESULTS>
                <RESULT eventid="1098" points="149" swimtime="00:00:37.98" resultid="4083" heatid="4243" lane="3" />
                <RESULT eventid="1107" points="133" swimtime="00:00:48.85" resultid="4084" heatid="4247" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Tenório De Almeida" birthdate="2003-12-13" gender="M" nation="BRA" athleteid="4078">
              <HANDICAP exception="TEA" free="18" />
              <RESULTS>
                <RESULT eventid="1111" points="145" swimtime="00:01:25.16" resultid="4079" heatid="4254" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="137" swimtime="00:00:42.82" resultid="4080" heatid="4222" lane="4" />
                <RESULT eventid="1098" points="170" swimtime="00:00:36.39" resultid="4081" heatid="4237" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1485" nation="BRA" region="PR" clubid="3874" name="Seleção de Campo Mourão" shortname="Campo Mourão">
          <ATHLETES>
            <ATHLETE firstname="Antonio" lastname="Paulino De Oliveira Junior" birthdate="1987-12-14" gender="M" nation="BRA" athleteid="3875">
              <HANDICAP exception="DV" breast="13" free="13" medley="13" />
              <RESULTS>
                <RESULT eventid="1090" points="109" swimtime="00:03:49.08" resultid="3876" heatid="4233" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.93" />
                    <SPLIT distance="100" swimtime="00:01:44.44" />
                    <SPLIT distance="150" swimtime="00:02:54.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1098" points="148" swimtime="00:00:38.11" resultid="3877" heatid="4239" lane="1" />
                <RESULT eventid="1107" points="131" swimtime="00:00:49.06" resultid="3878" heatid="4247" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tharcys" lastname="Gustavo Cussolin Batista" birthdate="2000-09-16" gender="M" nation="BRA" athleteid="3889">
              <HANDICAP exception="DF" free="10" />
              <RESULTS>
                <RESULT eventid="1111" points="294" swimtime="00:01:07.36" resultid="3890" heatid="4255" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="299" swimtime="00:00:32.51" resultid="3891" heatid="4228" lane="4" />
                <RESULT eventid="1098" points="290" swimtime="00:00:30.44" resultid="3892" heatid="4243" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Narciso De Melo" birthdate="2000-02-21" gender="M" nation="BRA" athleteid="3883">
              <HANDICAP exception="DF" free="5" />
              <RESULTS>
                <RESULT eventid="1066" status="DNS" swimtime="00:00:00.00" resultid="3884" heatid="4222" lane="5" />
                <RESULT eventid="1098" status="DNS" swimtime="00:00:00.00" resultid="3885" heatid="4241" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Erick" lastname="Campos De Jesus" birthdate="2008-03-14" gender="M" nation="BRA" athleteid="3879">
              <HANDICAP exception="DF" free="9" />
              <RESULTS>
                <RESULT eventid="1111" points="252" swimtime="00:01:10.92" resultid="3880" heatid="4256" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="233" swimtime="00:00:35.31" resultid="3881" heatid="4228" lane="6" />
                <RESULT eventid="1098" points="302" swimtime="00:00:30.04" resultid="3882" heatid="4242" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauê" lastname="Chagas" birthdate="2005-06-29" gender="M" nation="BRA" athleteid="3886">
              <HANDICAP exception="DF" breast="9" />
              <RESULTS>
                <RESULT eventid="1070" points="233" swimtime="00:01:29.83" resultid="3887" heatid="4224" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="246" swimtime="00:00:39.78" resultid="3888" heatid="4249" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CAMPO MOURÃO &quot;A&quot;">
              <RESULTS>
                <RESULT eventid="1086" status="WDR" swimtime="00:00:00.00" resultid="4264" heatid="4263" lane="4">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3879" number="1" />
                    <RELAYPOSITION athleteid="3883" number="2" />
                    <RELAYPOSITION athleteid="3886" number="3" />
                    <RELAYPOSITION athleteid="3889" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1116" status="WDR" swimtime="00:00:00.00" resultid="4276" heatid="4274" lane="2">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3879" number="1" />
                    <RELAYPOSITION athleteid="3883" number="2" />
                    <RELAYPOSITION athleteid="3886" number="3" />
                    <RELAYPOSITION athleteid="3889" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
  <TIMESTANDARDLISTS>
    <TIMESTANDARDLIST timestandardlistid="1764" code="S1" course="SCM" gender="M" handicap="1" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:03:07.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:17:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1766" code="S1" course="SCM" gender="F" handicap="1" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:05:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:22.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:20:00.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:22.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:22.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:22.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1820" code="S10" course="SCM" gender="M" handicap="10" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:33.45">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:33.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:21.15">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:01.15">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:43.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:37.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1822" code="S10" course="SCM" gender="F" handicap="10" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:11.15">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:26.15">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:21.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:56.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:46.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:11.15">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1826" code="S11" course="SCM" gender="M" handicap="11" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:27.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:01.15">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:37.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:35.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:41.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:02.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:41.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1828" code="S11" course="SCM" gender="F" handicap="11" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:42.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:08.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:42.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:58.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1832" code="S12" course="SCM" gender="M" handicap="12" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:58.45">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:21.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:58.45">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:32.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:28.45">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:56.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:58.45">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1834" code="S12" course="SCM" gender="F" handicap="12" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:23.45">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:56.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:13.45">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:08.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:47.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:52.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:36.15">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1838" code="S13" course="SCM" gender="M" handicap="13" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:52.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:22.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:36.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:38.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:58.45">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1840" code="S13" course="SCM" gender="F" handicap="13" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:11.15">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:52.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:07.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:02.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:43.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:47.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:11.15">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1844" code="S14" course="SCM" gender="M" handicap="14" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:45.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1846" code="S14" course="SCM" gender="F" handicap="14" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:20.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1772" code="S2" course="SCM" gender="M" handicap="2" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:09:35.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:07.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1774" code="S2" course="SCM" gender="F" handicap="2" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:03:57.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:15.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:12:30.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:20.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:07.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1850" code="S21" course="SCM" gender="M" handicap="21" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:25.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:10.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1852" code="S21" course="SCM" gender="F" handicap="21" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:03:00.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:45.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:20.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1778" code="S3" course="SCM" gender="M" handicap="3" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:11.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:55.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:46.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:46.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1780" code="S3" course="SCM" gender="F" handicap="3" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:50.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:11:52.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:07.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:07.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:55.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1784" code="S4" course="SCM" gender="M" handicap="4" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:42.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:07:05.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:11.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:33.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:27.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1786" code="S4" course="SCM" gender="F" handicap="4" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:57.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:10.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:08:20.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:11.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:58.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1790" code="S5" course="SCM" gender="M" handicap="5" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:58.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:36.15">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:11.15">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:06.15">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1792" code="S5" course="SCM" gender="F" handicap="5" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:52.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:45.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:42.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:33.45">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:33.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:18.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1796" code="S6" course="SCM" gender="M" handicap="6" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:56.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:52.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:06:33.45">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:56.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:08.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:11.15">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1798" code="S6" course="SCM" gender="F" handicap="6" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:33.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:32.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:18.45">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:56.15">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:27.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:05.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:42.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1802" code="S7" course="SCM" gender="M" handicap="7" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:58.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:17.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:42.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:53.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:02.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:46.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1804" code="S7" course="SCM" gender="F" handicap="7" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:03:26.15">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:17.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:05:18.45">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:21.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:03.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:36.15">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1808" code="S8" course="SCM" gender="M" handicap="8" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:52.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:05.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:35.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:22.30">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:52.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:56.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:42.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:58.45">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1810" code="S8" course="SCM" gender="F" handicap="8" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:15.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:55.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:11.15">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:41.15">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:33.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:08.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:00.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:30.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1814" code="S9" course="SCM" gender="M" handicap="9" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:01:37.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:46.15">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:58.45">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:23.45">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:10.00">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:48.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:50.00">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:37.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:40.00">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
    <TIMESTANDARDLIST timestandardlistid="1816" code="S9" course="SCM" gender="F" handicap="9" name="Índice para Pontuação (PARAJAPS)" type="MAXIMUM">
      <TIMESTANDARDS>
        <TIMESTANDARD swimtime="00:02:17.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:08.45">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:42.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:46.15">
          <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:04:03.45">
          <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:27.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:01:02.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:00:47.30">
          <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
        </TIMESTANDARD>
        <TIMESTANDARD swimtime="00:02:17.30">
          <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
        </TIMESTANDARD>
      </TIMESTANDARDS>
    </TIMESTANDARDLIST>
  </TIMESTANDARDLISTS>
</LENEX>
