<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.79125">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Curitiba" name="Torneio Regional da 1ª Região (Pré-Mirim/Sênior)" course="SCM" deadline="2024-02-26" entrystartdate="2024-02-16" entrytype="INVITATION" hostclub="Clube Curitibano" hostclub.url="https://clubecuritibano.com.br/" number="38296" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/evento/natacao/38296" startmethod="1" timing="AUTOMATIC" masters="F" withdrawuntil="2024-02-28" state="PR" nation="BRA">
      <AGEDATE value="2024-03-01" type="YEAR" />
      <POOL name="Parque Aquático do Clube Curitibano" lanemin="1" lanemax="8" />
      <FACILITY city="Curitiba" name="Parque Aquático do Clube Curitibano" nation="BRA" state="PR" street="Avenida Presidente Getúlio Vargas, 2857" street2="Água Verde" zip="80240-040" />
      <POINTTABLE pointtableid="3016" name="FINA Point Scoring" version="2023" />
      <QUALIFY from="2023-03-01" until="2024-02-29" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-03-01" daytime="15:10" endtime="18:14" name="1ª Etapa (Pré-Mirim/Petiz)" number="1" officialmeeting="15:30" warmupfrom="14:00" warmupuntil="15:00">
          <EVENTS>
            <EVENT eventid="1062" daytime="15:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1063" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2172" />
                    <RANKING order="2" place="2" resultid="2715" />
                    <RANKING order="3" place="3" resultid="2333" />
                    <RANKING order="4" place="4" resultid="1413" />
                    <RANKING order="5" place="5" resultid="2207" />
                    <RANKING order="6" place="6" resultid="2482" />
                    <RANKING order="7" place="7" resultid="3295" />
                    <RANKING order="8" place="8" resultid="2226" />
                    <RANKING order="9" place="-1" resultid="3201" />
                    <RANKING order="10" place="-1" resultid="2420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1064" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2116" />
                    <RANKING order="2" place="2" resultid="2076" />
                    <RANKING order="3" place="3" resultid="2081" />
                    <RANKING order="4" place="4" resultid="2477" />
                    <RANKING order="5" place="5" resultid="2141" />
                    <RANKING order="6" place="6" resultid="3324" />
                    <RANKING order="7" place="7" resultid="2343" />
                    <RANKING order="8" place="8" resultid="2277" />
                    <RANKING order="9" place="9" resultid="2798" />
                    <RANKING order="10" place="10" resultid="3345" />
                    <RANKING order="11" place="-1" resultid="2686" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3392" daytime="15:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3393" daytime="15:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3394" daytime="15:16" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1065" daytime="15:20" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1066" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2283" />
                    <RANKING order="2" place="2" resultid="1601" />
                    <RANKING order="3" place="3" resultid="2309" />
                    <RANKING order="4" place="4" resultid="2273" />
                    <RANKING order="5" place="5" resultid="2218" />
                    <RANKING order="6" place="6" resultid="2298" />
                    <RANKING order="7" place="7" resultid="3261" />
                    <RANKING order="8" place="8" resultid="2319" />
                    <RANKING order="9" place="9" resultid="2270" />
                    <RANKING order="10" place="10" resultid="3269" />
                    <RANKING order="11" place="11" resultid="2329" />
                    <RANKING order="12" place="12" resultid="2255" />
                    <RANKING order="13" place="13" resultid="2823" />
                    <RANKING order="14" place="-1" resultid="2237" />
                    <RANKING order="15" place="-1" resultid="3214" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2102" />
                    <RANKING order="2" place="2" resultid="3169" />
                    <RANKING order="3" place="3" resultid="2132" />
                    <RANKING order="4" place="4" resultid="2147" />
                    <RANKING order="5" place="5" resultid="2339" />
                    <RANKING order="6" place="6" resultid="2097" />
                    <RANKING order="7" place="7" resultid="2223" />
                    <RANKING order="8" place="8" resultid="2314" />
                    <RANKING order="9" place="9" resultid="3247" />
                    <RANKING order="10" place="10" resultid="3291" />
                    <RANKING order="11" place="11" resultid="2288" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3395" daytime="15:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3396" daytime="15:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3397" daytime="15:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3398" daytime="15:30" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1068" daytime="15:34" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1069" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2552" />
                    <RANKING order="2" place="2" resultid="2517" />
                    <RANKING order="3" place="3" resultid="2577" />
                    <RANKING order="4" place="4" resultid="2537" />
                    <RANKING order="5" place="5" resultid="2582" />
                    <RANKING order="6" place="6" resultid="3387" />
                    <RANKING order="7" place="7" resultid="2682" />
                    <RANKING order="8" place="8" resultid="2726" />
                    <RANKING order="9" place="9" resultid="2512" />
                    <RANKING order="10" place="10" resultid="2650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3193" />
                    <RANKING order="2" place="2" resultid="2370" />
                    <RANKING order="3" place="3" resultid="3364" />
                    <RANKING order="4" place="4" resultid="2498" />
                    <RANKING order="5" place="5" resultid="2473" />
                    <RANKING order="6" place="6" resultid="1714" />
                    <RANKING order="7" place="7" resultid="1404" />
                    <RANKING order="8" place="8" resultid="2375" />
                    <RANKING order="9" place="9" resultid="3300" />
                    <RANKING order="10" place="10" resultid="3018" />
                    <RANKING order="11" place="11" resultid="1665" />
                    <RANKING order="12" place="12" resultid="3353" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3399" daytime="15:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3400" daytime="15:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3401" daytime="15:38" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1071" daytime="15:40" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1072" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2507" />
                    <RANKING order="2" place="2" resultid="2677" />
                    <RANKING order="3" place="3" resultid="3278" />
                    <RANKING order="4" place="4" resultid="2557" />
                    <RANKING order="5" place="5" resultid="2645" />
                    <RANKING order="6" place="6" resultid="2700" />
                    <RANKING order="7" place="7" resultid="2730" />
                    <RANKING order="8" place="8" resultid="2672" />
                    <RANKING order="9" place="9" resultid="2658" />
                    <RANKING order="10" place="10" resultid="2734" />
                    <RANKING order="11" place="-1" resultid="2635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2390" />
                    <RANKING order="2" place="2" resultid="3242" />
                    <RANKING order="3" place="3" resultid="3317" />
                    <RANKING order="4" place="4" resultid="1422" />
                    <RANKING order="5" place="5" resultid="2443" />
                    <RANKING order="6" place="6" resultid="2963" />
                    <RANKING order="7" place="7" resultid="3321" />
                    <RANKING order="8" place="8" resultid="2385" />
                    <RANKING order="9" place="9" resultid="2453" />
                    <RANKING order="10" place="-1" resultid="2426" />
                    <RANKING order="11" place="-1" resultid="2430" />
                    <RANKING order="12" place="-1" resultid="2503" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3402" daytime="15:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3403" daytime="15:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3404" daytime="15:46" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1074" daytime="15:48" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1075" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2250" />
                    <RANKING order="2" place="2" resultid="2168" />
                    <RANKING order="3" place="3" resultid="2242" />
                    <RANKING order="4" place="4" resultid="2782" />
                    <RANKING order="5" place="5" resultid="1586" />
                    <RANKING order="6" place="6" resultid="2354" />
                    <RANKING order="7" place="7" resultid="2265" />
                    <RANKING order="8" place="8" resultid="1489" />
                    <RANKING order="9" place="9" resultid="2260" />
                    <RANKING order="10" place="10" resultid="2903" />
                    <RANKING order="11" place="11" resultid="1414" />
                    <RANKING order="12" place="12" resultid="3250" />
                    <RANKING order="13" place="13" resultid="2438" />
                    <RANKING order="14" place="14" resultid="3264" />
                    <RANKING order="15" place="15" resultid="3390" />
                    <RANKING order="16" place="16" resultid="3056" />
                    <RANKING order="17" place="17" resultid="3296" />
                    <RANKING order="18" place="-1" resultid="3228" />
                    <RANKING order="19" place="-1" resultid="1485" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1076" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2293" />
                    <RANKING order="2" place="2" resultid="2478" />
                    <RANKING order="3" place="3" resultid="2213" />
                    <RANKING order="4" place="4" resultid="2082" />
                    <RANKING order="5" place="5" resultid="2203" />
                    <RANKING order="6" place="6" resultid="2127" />
                    <RANKING order="7" place="7" resultid="3223" />
                    <RANKING order="8" place="8" resultid="3325" />
                    <RANKING order="9" place="9" resultid="2122" />
                    <RANKING order="10" place="10" resultid="3188" />
                    <RANKING order="11" place="11" resultid="2142" />
                    <RANKING order="12" place="12" resultid="1475" />
                    <RANKING order="13" place="13" resultid="2278" />
                    <RANKING order="14" place="14" resultid="2771" />
                    <RANKING order="15" place="15" resultid="1396" />
                    <RANKING order="16" place="16" resultid="1426" />
                    <RANKING order="17" place="17" resultid="2344" />
                    <RANKING order="18" place="18" resultid="3037" />
                    <RANKING order="19" place="19" resultid="1654" />
                    <RANKING order="20" place="20" resultid="3346" />
                    <RANKING order="21" place="-1" resultid="1717" />
                    <RANKING order="22" place="-1" resultid="2654" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3405" daytime="15:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3406" daytime="15:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3407" daytime="15:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3408" daytime="15:56" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3409" daytime="16:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3410" daytime="16:02" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1077" daytime="16:04" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1078" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1386" />
                    <RANKING order="2" place="2" resultid="3273" />
                    <RANKING order="3" place="3" resultid="2163" />
                    <RANKING order="4" place="4" resultid="3206" />
                    <RANKING order="5" place="5" resultid="2493" />
                    <RANKING order="6" place="6" resultid="2324" />
                    <RANKING order="7" place="7" resultid="2232" />
                    <RANKING order="8" place="8" resultid="3268" />
                    <RANKING order="9" place="9" resultid="3253" />
                    <RANKING order="10" place="10" resultid="3238" />
                    <RANKING order="11" place="11" resultid="3336" />
                    <RANKING order="12" place="-1" resultid="2822" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2101" />
                    <RANKING order="2" place="2" resultid="2879" />
                    <RANKING order="3" place="3" resultid="2062" />
                    <RANKING order="4" place="4" resultid="2107" />
                    <RANKING order="5" place="5" resultid="2092" />
                    <RANKING order="6" place="6" resultid="2067" />
                    <RANKING order="7" place="7" resultid="2087" />
                    <RANKING order="8" place="7" resultid="2112" />
                    <RANKING order="9" place="9" resultid="1498" />
                    <RANKING order="10" place="10" resultid="2072" />
                    <RANKING order="11" place="11" resultid="2137" />
                    <RANKING order="12" place="12" resultid="3211" />
                    <RANKING order="13" place="13" resultid="2131" />
                    <RANKING order="14" place="14" resultid="2158" />
                    <RANKING order="15" place="15" resultid="3313" />
                    <RANKING order="16" place="16" resultid="2313" />
                    <RANKING order="17" place="17" resultid="1590" />
                    <RANKING order="18" place="18" resultid="1516" />
                    <RANKING order="19" place="19" resultid="2222" />
                    <RANKING order="20" place="20" resultid="3349" />
                    <RANKING order="21" place="21" resultid="2287" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3411" daytime="16:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3412" daytime="16:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3413" daytime="16:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3414" daytime="16:12" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3415" daytime="16:14" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1080" daytime="16:18" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1081" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2984" />
                    <RANKING order="2" place="2" resultid="2998" />
                    <RANKING order="3" place="3" resultid="2562" />
                    <RANKING order="4" place="4" resultid="2640" />
                    <RANKING order="5" place="5" resultid="2667" />
                    <RANKING order="6" place="6" resultid="3386" />
                    <RANKING order="7" place="7" resultid="1508" />
                    <RANKING order="8" place="8" resultid="2527" />
                    <RANKING order="9" place="9" resultid="2572" />
                    <RANKING order="10" place="10" resultid="2725" />
                    <RANKING order="11" place="11" resultid="2649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3299" />
                    <RANKING order="2" place="2" resultid="1391" />
                    <RANKING order="3" place="3" resultid="2488" />
                    <RANKING order="4" place="4" resultid="3363" />
                    <RANKING order="5" place="5" resultid="2542" />
                    <RANKING order="6" place="6" resultid="2587" />
                    <RANKING order="7" place="7" resultid="3305" />
                    <RANKING order="8" place="8" resultid="2374" />
                    <RANKING order="9" place="9" resultid="2458" />
                    <RANKING order="10" place="10" resultid="2463" />
                    <RANKING order="11" place="11" resultid="3017" />
                    <RANKING order="12" place="12" resultid="3003" />
                    <RANKING order="13" place="13" resultid="3352" />
                    <RANKING order="14" place="-1" resultid="2434" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3416" daytime="16:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3417" daytime="16:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3418" daytime="16:22" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3419" daytime="16:26" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1083" daytime="16:28" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1084" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2522" />
                    <RANKING order="2" place="2" resultid="2567" />
                    <RANKING order="3" place="3" resultid="2556" />
                    <RANKING order="4" place="4" resultid="2644" />
                    <RANKING order="5" place="5" resultid="2721" />
                    <RANKING order="6" place="6" resultid="2657" />
                    <RANKING order="7" place="7" resultid="2634" />
                    <RANKING order="8" place="8" resultid="2671" />
                    <RANKING order="9" place="9" resultid="2733" />
                    <RANKING order="10" place="10" resultid="2729" />
                    <RANKING order="11" place="11" resultid="2705" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2349" />
                    <RANKING order="2" place="2" resultid="2615" />
                    <RANKING order="3" place="3" resultid="1409" />
                    <RANKING order="4" place="4" resultid="2380" />
                    <RANKING order="5" place="5" resultid="1502" />
                    <RANKING order="6" place="6" resultid="2384" />
                    <RANKING order="7" place="7" resultid="2547" />
                    <RANKING order="8" place="8" resultid="3233" />
                    <RANKING order="9" place="9" resultid="3309" />
                    <RANKING order="10" place="10" resultid="2532" />
                    <RANKING order="11" place="11" resultid="3316" />
                    <RANKING order="12" place="12" resultid="2468" />
                    <RANKING order="13" place="13" resultid="2663" />
                    <RANKING order="14" place="14" resultid="3257" />
                    <RANKING order="15" place="15" resultid="2452" />
                    <RANKING order="16" place="16" resultid="3334" />
                    <RANKING order="17" place="-1" resultid="2448" />
                    <RANKING order="18" place="-1" resultid="2502" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3420" daytime="16:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3421" daytime="16:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3422" daytime="16:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3423" daytime="16:38" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1086" daytime="16:40" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1087" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2781" />
                    <RANKING order="2" place="2" resultid="2167" />
                    <RANKING order="3" place="3" resultid="2173" />
                    <RANKING order="4" place="4" resultid="2716" />
                    <RANKING order="5" place="5" resultid="3227" />
                    <RANKING order="6" place="6" resultid="2208" />
                    <RANKING order="7" place="7" resultid="2249" />
                    <RANKING order="8" place="8" resultid="2334" />
                    <RANKING order="9" place="9" resultid="3202" />
                    <RANKING order="10" place="10" resultid="1585" />
                    <RANKING order="11" place="11" resultid="2353" />
                    <RANKING order="12" place="12" resultid="2241" />
                    <RANKING order="13" place="13" resultid="2264" />
                    <RANKING order="14" place="14" resultid="2437" />
                    <RANKING order="15" place="15" resultid="1488" />
                    <RANKING order="16" place="16" resultid="2483" />
                    <RANKING order="17" place="17" resultid="2902" />
                    <RANKING order="18" place="18" resultid="2421" />
                    <RANKING order="19" place="19" resultid="2259" />
                    <RANKING order="20" place="20" resultid="1484" />
                    <RANKING order="21" place="21" resultid="2227" />
                    <RANKING order="22" place="22" resultid="3055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2292" />
                    <RANKING order="2" place="2" resultid="2077" />
                    <RANKING order="3" place="3" resultid="2212" />
                    <RANKING order="4" place="4" resultid="2121" />
                    <RANKING order="5" place="5" resultid="2126" />
                    <RANKING order="6" place="6" resultid="2202" />
                    <RANKING order="7" place="7" resultid="3222" />
                    <RANKING order="8" place="8" resultid="1641" />
                    <RANKING order="9" place="9" resultid="3187" />
                    <RANKING order="10" place="10" resultid="2687" />
                    <RANKING order="11" place="11" resultid="2117" />
                    <RANKING order="12" place="12" resultid="1395" />
                    <RANKING order="13" place="13" resultid="3036" />
                    <RANKING order="14" place="14" resultid="1425" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3424" daytime="16:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3425" daytime="16:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3426" daytime="16:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3427" daytime="16:56" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3428" daytime="17:00" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1089" daytime="17:04" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1090" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1385" />
                    <RANKING order="2" place="2" resultid="1600" />
                    <RANKING order="3" place="3" resultid="3272" />
                    <RANKING order="4" place="4" resultid="2308" />
                    <RANKING order="5" place="5" resultid="2272" />
                    <RANKING order="6" place="6" resultid="2297" />
                    <RANKING order="7" place="7" resultid="2162" />
                    <RANKING order="8" place="8" resultid="2323" />
                    <RANKING order="9" place="9" resultid="2282" />
                    <RANKING order="10" place="10" resultid="2492" />
                    <RANKING order="11" place="11" resultid="2217" />
                    <RANKING order="12" place="12" resultid="2254" />
                    <RANKING order="13" place="13" resultid="2231" />
                    <RANKING order="14" place="14" resultid="2328" />
                    <RANKING order="15" place="15" resultid="3260" />
                    <RANKING order="16" place="16" resultid="2318" />
                    <RANKING order="17" place="17" resultid="2269" />
                    <RANKING order="18" place="18" resultid="3237" />
                    <RANKING order="19" place="-1" resultid="2236" />
                    <RANKING order="20" place="-1" resultid="3213" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2111" />
                    <RANKING order="2" place="2" resultid="2061" />
                    <RANKING order="3" place="3" resultid="2136" />
                    <RANKING order="4" place="4" resultid="3168" />
                    <RANKING order="5" place="5" resultid="2106" />
                    <RANKING order="6" place="6" resultid="2066" />
                    <RANKING order="7" place="7" resultid="2091" />
                    <RANKING order="8" place="8" resultid="2071" />
                    <RANKING order="9" place="9" resultid="2146" />
                    <RANKING order="10" place="10" resultid="2086" />
                    <RANKING order="11" place="11" resultid="2338" />
                    <RANKING order="12" place="12" resultid="2878" />
                    <RANKING order="13" place="13" resultid="3210" />
                    <RANKING order="14" place="14" resultid="2157" />
                    <RANKING order="15" place="15" resultid="1497" />
                    <RANKING order="16" place="16" resultid="2096" />
                    <RANKING order="17" place="17" resultid="3290" />
                    <RANKING order="18" place="18" resultid="3360" />
                    <RANKING order="19" place="19" resultid="3246" />
                    <RANKING order="20" place="20" resultid="1515" />
                    <RANKING order="21" place="-1" resultid="1645" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3429" daytime="17:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3430" daytime="17:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3431" daytime="17:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3432" daytime="17:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3433" daytime="17:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3434" daytime="17:28" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1092" daytime="17:32" gender="F" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1093" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2983" />
                    <RANKING order="2" place="2" resultid="2536" />
                    <RANKING order="3" place="3" resultid="2997" />
                    <RANKING order="4" place="4" resultid="2561" />
                    <RANKING order="5" place="5" resultid="2576" />
                    <RANKING order="6" place="6" resultid="2581" />
                    <RANKING order="7" place="7" resultid="2516" />
                    <RANKING order="8" place="8" resultid="2666" />
                    <RANKING order="9" place="9" resultid="2639" />
                    <RANKING order="10" place="10" resultid="2551" />
                    <RANKING order="11" place="11" resultid="2571" />
                    <RANKING order="12" place="12" resultid="2511" />
                    <RANKING order="13" place="13" resultid="2681" />
                    <RANKING order="14" place="14" resultid="2526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3192" />
                    <RANKING order="2" place="2" resultid="2369" />
                    <RANKING order="3" place="3" resultid="1390" />
                    <RANKING order="4" place="4" resultid="2457" />
                    <RANKING order="5" place="5" resultid="2472" />
                    <RANKING order="6" place="6" resultid="2586" />
                    <RANKING order="7" place="7" resultid="1403" />
                    <RANKING order="8" place="8" resultid="2497" />
                    <RANKING order="9" place="9" resultid="2487" />
                    <RANKING order="10" place="10" resultid="2541" />
                    <RANKING order="11" place="11" resultid="2462" />
                    <RANKING order="12" place="12" resultid="3304" />
                    <RANKING order="13" place="13" resultid="3002" />
                    <RANKING order="14" place="-1" resultid="2433" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3435" daytime="17:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3436" daytime="17:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3437" daytime="17:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3438" daytime="17:42" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1095" daytime="17:46" gender="M" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1096" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2521" />
                    <RANKING order="2" place="2" resultid="3277" />
                    <RANKING order="3" place="3" resultid="2506" />
                    <RANKING order="4" place="4" resultid="2566" />
                    <RANKING order="5" place="5" resultid="2676" />
                    <RANKING order="6" place="6" resultid="2699" />
                    <RANKING order="7" place="7" resultid="2720" />
                    <RANKING order="8" place="-1" resultid="2704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2348" />
                    <RANKING order="2" place="2" resultid="2389" />
                    <RANKING order="3" place="3" resultid="1408" />
                    <RANKING order="4" place="4" resultid="2379" />
                    <RANKING order="5" place="5" resultid="3241" />
                    <RANKING order="6" place="6" resultid="2546" />
                    <RANKING order="7" place="7" resultid="1421" />
                    <RANKING order="8" place="8" resultid="3232" />
                    <RANKING order="9" place="9" resultid="1501" />
                    <RANKING order="10" place="10" resultid="2447" />
                    <RANKING order="11" place="11" resultid="2614" />
                    <RANKING order="12" place="12" resultid="2962" />
                    <RANKING order="13" place="13" resultid="2467" />
                    <RANKING order="14" place="14" resultid="2442" />
                    <RANKING order="15" place="15" resultid="3308" />
                    <RANKING order="16" place="16" resultid="2531" />
                    <RANKING order="17" place="17" resultid="3320" />
                    <RANKING order="18" place="18" resultid="3256" />
                    <RANKING order="19" place="19" resultid="2662" />
                    <RANKING order="20" place="20" resultid="3333" />
                    <RANKING order="21" place="-1" resultid="2425" />
                    <RANKING order="22" place="-1" resultid="2429" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3439" daytime="17:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3440" daytime="17:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3441" daytime="17:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3442" daytime="17:56" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-03-02" daytime="09:10" endtime="11:07" name="2ª Etapa (Pré-Mirim/Petiz)" number="2" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1098" daytime="09:10" gender="F" number="13" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1099" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1100" daytime="09:10" gender="M" number="14" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1101" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1102" daytime="09:10" gender="F" number="15" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1103" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2174" />
                    <RANKING order="2" place="2" resultid="2783" />
                    <RANKING order="3" place="3" resultid="2209" />
                    <RANKING order="4" place="4" resultid="2169" />
                    <RANKING order="5" place="5" resultid="2335" />
                    <RANKING order="6" place="6" resultid="3229" />
                    <RANKING order="7" place="7" resultid="2243" />
                    <RANKING order="8" place="8" resultid="1587" />
                    <RANKING order="9" place="9" resultid="1415" />
                    <RANKING order="10" place="10" resultid="2266" />
                    <RANKING order="11" place="11" resultid="2355" />
                    <RANKING order="12" place="12" resultid="2484" />
                    <RANKING order="13" place="13" resultid="2422" />
                    <RANKING order="14" place="14" resultid="3057" />
                    <RANKING order="15" place="15" resultid="2228" />
                    <RANKING order="16" place="-1" resultid="2251" />
                    <RANKING order="17" place="-1" resultid="2261" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1104" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2083" />
                    <RANKING order="2" place="2" resultid="2078" />
                    <RANKING order="3" place="3" resultid="2123" />
                    <RANKING order="4" place="4" resultid="2214" />
                    <RANKING order="5" place="5" resultid="2479" />
                    <RANKING order="6" place="6" resultid="2204" />
                    <RANKING order="7" place="7" resultid="2118" />
                    <RANKING order="8" place="8" resultid="2143" />
                    <RANKING order="9" place="9" resultid="3189" />
                    <RANKING order="10" place="10" resultid="3224" />
                    <RANKING order="11" place="11" resultid="2799" />
                    <RANKING order="12" place="12" resultid="2688" />
                    <RANKING order="13" place="13" resultid="3326" />
                    <RANKING order="14" place="14" resultid="1718" />
                    <RANKING order="15" place="15" resultid="2279" />
                    <RANKING order="16" place="16" resultid="2345" />
                    <RANKING order="17" place="17" resultid="3038" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3443" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3444" daytime="09:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3445" daytime="09:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3446" daytime="09:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3447" daytime="09:22" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1105" daytime="09:26" gender="M" number="16" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1106" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1602" />
                    <RANKING order="2" place="2" resultid="2310" />
                    <RANKING order="3" place="3" resultid="2284" />
                    <RANKING order="4" place="4" resultid="3274" />
                    <RANKING order="5" place="5" resultid="2274" />
                    <RANKING order="6" place="6" resultid="3215" />
                    <RANKING order="7" place="7" resultid="2325" />
                    <RANKING order="8" place="8" resultid="2494" />
                    <RANKING order="9" place="9" resultid="3207" />
                    <RANKING order="10" place="10" resultid="2233" />
                    <RANKING order="11" place="11" resultid="2320" />
                    <RANKING order="12" place="12" resultid="2824" />
                    <RANKING order="13" place="13" resultid="2330" />
                    <RANKING order="14" place="-1" resultid="2238" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1107" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2103" />
                    <RANKING order="2" place="2" resultid="2093" />
                    <RANKING order="3" place="3" resultid="3170" />
                    <RANKING order="4" place="4" resultid="2133" />
                    <RANKING order="5" place="5" resultid="2108" />
                    <RANKING order="6" place="6" resultid="2148" />
                    <RANKING order="7" place="7" resultid="2088" />
                    <RANKING order="8" place="8" resultid="2880" />
                    <RANKING order="9" place="9" resultid="1646" />
                    <RANKING order="10" place="10" resultid="2098" />
                    <RANKING order="11" place="11" resultid="1591" />
                    <RANKING order="12" place="12" resultid="2315" />
                    <RANKING order="13" place="13" resultid="2289" />
                    <RANKING order="14" place="-1" resultid="2159" />
                    <RANKING order="15" place="-1" resultid="3046" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3448" daytime="09:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3449" daytime="09:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3450" daytime="09:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3451" daytime="09:34" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1108" daytime="09:38" gender="F" number="17" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1109" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2985" />
                    <RANKING order="2" place="2" resultid="2563" />
                    <RANKING order="3" place="3" resultid="2538" />
                    <RANKING order="4" place="4" resultid="2999" />
                    <RANKING order="5" place="5" resultid="2518" />
                    <RANKING order="6" place="6" resultid="2578" />
                    <RANKING order="7" place="7" resultid="2583" />
                    <RANKING order="8" place="8" resultid="2573" />
                    <RANKING order="9" place="9" resultid="2668" />
                    <RANKING order="10" place="10" resultid="2641" />
                    <RANKING order="11" place="11" resultid="2513" />
                    <RANKING order="12" place="12" resultid="2683" />
                    <RANKING order="13" place="13" resultid="2553" />
                    <RANKING order="14" place="14" resultid="2528" />
                    <RANKING order="15" place="15" resultid="2651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1110" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2371" />
                    <RANKING order="2" place="2" resultid="3194" />
                    <RANKING order="3" place="3" resultid="2588" />
                    <RANKING order="4" place="4" resultid="2459" />
                    <RANKING order="5" place="5" resultid="2474" />
                    <RANKING order="6" place="6" resultid="3301" />
                    <RANKING order="7" place="7" resultid="3365" />
                    <RANKING order="8" place="8" resultid="2543" />
                    <RANKING order="9" place="9" resultid="2499" />
                    <RANKING order="10" place="10" resultid="2376" />
                    <RANKING order="11" place="11" resultid="2464" />
                    <RANKING order="12" place="12" resultid="1392" />
                    <RANKING order="13" place="13" resultid="1405" />
                    <RANKING order="14" place="14" resultid="2489" />
                    <RANKING order="15" place="15" resultid="3019" />
                    <RANKING order="16" place="16" resultid="3354" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3452" daytime="09:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3453" daytime="09:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3454" daytime="09:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3455" daytime="09:44" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1111" daytime="09:48" gender="M" number="18" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1112" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2523" />
                    <RANKING order="2" place="2" resultid="3279" />
                    <RANKING order="3" place="3" resultid="2558" />
                    <RANKING order="4" place="4" resultid="2568" />
                    <RANKING order="5" place="5" resultid="2678" />
                    <RANKING order="6" place="6" resultid="2508" />
                    <RANKING order="7" place="7" resultid="2646" />
                    <RANKING order="8" place="8" resultid="2701" />
                    <RANKING order="9" place="9" resultid="2673" />
                    <RANKING order="10" place="10" resultid="2735" />
                    <RANKING order="11" place="11" resultid="2722" />
                    <RANKING order="12" place="12" resultid="2659" />
                    <RANKING order="13" place="13" resultid="2706" />
                    <RANKING order="14" place="-1" resultid="2636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2350" />
                    <RANKING order="2" place="2" resultid="2391" />
                    <RANKING order="3" place="3" resultid="2381" />
                    <RANKING order="4" place="4" resultid="2548" />
                    <RANKING order="5" place="5" resultid="2386" />
                    <RANKING order="6" place="6" resultid="2449" />
                    <RANKING order="7" place="7" resultid="2469" />
                    <RANKING order="8" place="8" resultid="3243" />
                    <RANKING order="9" place="9" resultid="1410" />
                    <RANKING order="10" place="10" resultid="2444" />
                    <RANKING order="11" place="11" resultid="3234" />
                    <RANKING order="12" place="12" resultid="2616" />
                    <RANKING order="13" place="13" resultid="3310" />
                    <RANKING order="14" place="14" resultid="2533" />
                    <RANKING order="15" place="15" resultid="2454" />
                    <RANKING order="16" place="-1" resultid="2964" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3456" daytime="09:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3457" daytime="09:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3458" daytime="09:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3459" daytime="09:54" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1114" daytime="09:56" gender="F" number="19" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1115" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1662" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3460" daytime="09:56" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1116" daytime="09:58" gender="M" number="20" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1117" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1118" daytime="09:58" gender="F" number="21" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1119" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2784" />
                    <RANKING order="2" place="2" resultid="2175" />
                    <RANKING order="3" place="3" resultid="2717" />
                    <RANKING order="4" place="4" resultid="3203" />
                    <RANKING order="5" place="5" resultid="2244" />
                    <RANKING order="6" place="6" resultid="2356" />
                    <RANKING order="7" place="7" resultid="3265" />
                    <RANKING order="8" place="-1" resultid="2170" />
                    <RANKING order="9" place="-1" resultid="2439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2294" />
                    <RANKING order="2" place="2" resultid="2128" />
                    <RANKING order="3" place="3" resultid="2084" />
                    <RANKING order="4" place="4" resultid="2144" />
                    <RANKING order="5" place="5" resultid="1642" />
                    <RANKING order="6" place="6" resultid="1476" />
                    <RANKING order="7" place="7" resultid="2800" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3461" daytime="09:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3462" daytime="10:02" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1121" daytime="10:06" gender="M" number="22" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1122" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1387" />
                    <RANKING order="2" place="2" resultid="2164" />
                    <RANKING order="3" place="3" resultid="2219" />
                    <RANKING order="4" place="4" resultid="3216" />
                    <RANKING order="5" place="5" resultid="2256" />
                    <RANKING order="6" place="-1" resultid="2299" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1123" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2138" />
                    <RANKING order="2" place="2" resultid="2063" />
                    <RANKING order="3" place="3" resultid="2113" />
                    <RANKING order="4" place="4" resultid="2340" />
                    <RANKING order="5" place="5" resultid="2068" />
                    <RANKING order="6" place="6" resultid="2073" />
                    <RANKING order="7" place="-1" resultid="3292" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3463" daytime="10:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3464" daytime="10:08" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1124" daytime="10:12" gender="F" number="23" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1125" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1126" daytime="10:12" gender="M" number="24" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1127" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1128" daytime="10:12" gender="F" number="25" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1129" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2986" />
                    <RANKING order="2" place="2" resultid="3000" />
                    <RANKING order="3" place="3" resultid="2539" />
                    <RANKING order="4" place="4" resultid="2564" />
                    <RANKING order="5" place="5" resultid="2579" />
                    <RANKING order="6" place="6" resultid="2519" />
                    <RANKING order="7" place="7" resultid="2584" />
                    <RANKING order="8" place="8" resultid="3388" />
                    <RANKING order="9" place="9" resultid="2669" />
                    <RANKING order="10" place="10" resultid="1509" />
                    <RANKING order="11" place="11" resultid="2574" />
                    <RANKING order="12" place="12" resultid="2642" />
                    <RANKING order="13" place="13" resultid="2514" />
                    <RANKING order="14" place="14" resultid="2554" />
                    <RANKING order="15" place="15" resultid="2652" />
                    <RANKING order="16" place="16" resultid="2727" />
                    <RANKING order="17" place="17" resultid="2529" />
                    <RANKING order="18" place="-1" resultid="2684" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3195" />
                    <RANKING order="2" place="2" resultid="2372" />
                    <RANKING order="3" place="3" resultid="3302" />
                    <RANKING order="4" place="4" resultid="1393" />
                    <RANKING order="5" place="5" resultid="2475" />
                    <RANKING order="6" place="6" resultid="3366" />
                    <RANKING order="7" place="7" resultid="2490" />
                    <RANKING order="8" place="8" resultid="2544" />
                    <RANKING order="9" place="9" resultid="2460" />
                    <RANKING order="10" place="10" resultid="1406" />
                    <RANKING order="11" place="11" resultid="3306" />
                    <RANKING order="12" place="12" resultid="2465" />
                    <RANKING order="13" place="12" resultid="2500" />
                    <RANKING order="14" place="14" resultid="2377" />
                    <RANKING order="15" place="15" resultid="3004" />
                    <RANKING order="16" place="16" resultid="1715" />
                    <RANKING order="17" place="17" resultid="1666" />
                    <RANKING order="18" place="18" resultid="2435" />
                    <RANKING order="19" place="19" resultid="3355" />
                    <RANKING order="20" place="20" resultid="3020" />
                    <RANKING order="21" place="21" resultid="2995" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3465" daytime="10:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3466" daytime="10:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3467" daytime="10:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3468" daytime="10:18" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3469" daytime="10:20" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1131" daytime="10:24" gender="M" number="26" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1132" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2524" />
                    <RANKING order="2" place="2" resultid="3280" />
                    <RANKING order="3" place="3" resultid="2509" />
                    <RANKING order="4" place="4" resultid="2569" />
                    <RANKING order="5" place="5" resultid="2559" />
                    <RANKING order="6" place="6" resultid="2647" />
                    <RANKING order="7" place="7" resultid="2674" />
                    <RANKING order="8" place="8" resultid="2679" />
                    <RANKING order="9" place="9" resultid="2660" />
                    <RANKING order="10" place="10" resultid="2637" />
                    <RANKING order="11" place="11" resultid="2723" />
                    <RANKING order="12" place="12" resultid="2731" />
                    <RANKING order="13" place="13" resultid="2702" />
                    <RANKING order="14" place="14" resultid="2707" />
                    <RANKING order="15" place="15" resultid="2736" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1133" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2392" />
                    <RANKING order="2" place="2" resultid="2351" />
                    <RANKING order="3" place="3" resultid="1411" />
                    <RANKING order="4" place="4" resultid="2382" />
                    <RANKING order="5" place="5" resultid="3244" />
                    <RANKING order="6" place="6" resultid="1423" />
                    <RANKING order="7" place="7" resultid="2549" />
                    <RANKING order="8" place="8" resultid="1503" />
                    <RANKING order="9" place="9" resultid="2617" />
                    <RANKING order="10" place="10" resultid="2450" />
                    <RANKING order="11" place="11" resultid="3235" />
                    <RANKING order="12" place="12" resultid="2387" />
                    <RANKING order="13" place="13" resultid="2445" />
                    <RANKING order="14" place="14" resultid="2470" />
                    <RANKING order="15" place="15" resultid="2534" />
                    <RANKING order="16" place="16" resultid="3318" />
                    <RANKING order="17" place="17" resultid="3311" />
                    <RANKING order="18" place="18" resultid="3258" />
                    <RANKING order="19" place="19" resultid="3322" />
                    <RANKING order="20" place="20" resultid="2664" />
                    <RANKING order="21" place="21" resultid="2455" />
                    <RANKING order="22" place="-1" resultid="2427" />
                    <RANKING order="23" place="-1" resultid="2431" />
                    <RANKING order="24" place="-1" resultid="2504" />
                    <RANKING order="25" place="-1" resultid="2965" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3470" daytime="10:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3471" daytime="10:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3472" daytime="10:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3473" daytime="10:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3474" daytime="10:32" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1134" daytime="10:34" gender="F" number="27" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1135" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1663" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3475" daytime="10:34" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1136" daytime="10:36" gender="M" number="28" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="25" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1137" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1138" daytime="10:36" gender="F" number="29" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1139" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2210" />
                    <RANKING order="2" place="2" resultid="2252" />
                    <RANKING order="3" place="3" resultid="2718" />
                    <RANKING order="4" place="4" resultid="2336" />
                    <RANKING order="5" place="5" resultid="3230" />
                    <RANKING order="6" place="6" resultid="1588" />
                    <RANKING order="7" place="7" resultid="3204" />
                    <RANKING order="8" place="8" resultid="1416" />
                    <RANKING order="9" place="9" resultid="2267" />
                    <RANKING order="10" place="10" resultid="1490" />
                    <RANKING order="11" place="11" resultid="2904" />
                    <RANKING order="12" place="12" resultid="2423" />
                    <RANKING order="13" place="13" resultid="3251" />
                    <RANKING order="14" place="14" resultid="1486" />
                    <RANKING order="15" place="15" resultid="3266" />
                    <RANKING order="16" place="16" resultid="2485" />
                    <RANKING order="17" place="17" resultid="2814" />
                    <RANKING order="18" place="18" resultid="2440" />
                    <RANKING order="19" place="19" resultid="3058" />
                    <RANKING order="20" place="20" resultid="2229" />
                    <RANKING order="21" place="21" resultid="3391" />
                    <RANKING order="22" place="22" resultid="3297" />
                    <RANKING order="23" place="-1" resultid="2262" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1140" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2295" />
                    <RANKING order="2" place="2" resultid="2079" />
                    <RANKING order="3" place="3" resultid="2215" />
                    <RANKING order="4" place="4" resultid="2129" />
                    <RANKING order="5" place="5" resultid="2205" />
                    <RANKING order="6" place="6" resultid="2124" />
                    <RANKING order="7" place="7" resultid="2480" />
                    <RANKING order="8" place="8" resultid="3190" />
                    <RANKING order="9" place="9" resultid="3225" />
                    <RANKING order="10" place="10" resultid="2689" />
                    <RANKING order="11" place="11" resultid="2119" />
                    <RANKING order="12" place="12" resultid="1643" />
                    <RANKING order="13" place="12" resultid="3327" />
                    <RANKING order="14" place="14" resultid="1477" />
                    <RANKING order="15" place="15" resultid="1719" />
                    <RANKING order="16" place="16" resultid="2280" />
                    <RANKING order="17" place="17" resultid="2346" />
                    <RANKING order="18" place="18" resultid="3039" />
                    <RANKING order="19" place="19" resultid="2772" />
                    <RANKING order="20" place="20" resultid="1427" />
                    <RANKING order="21" place="21" resultid="1655" />
                    <RANKING order="22" place="22" resultid="3347" />
                    <RANKING order="23" place="-1" resultid="2655" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3476" daytime="10:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3477" daytime="10:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3478" daytime="10:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3479" daytime="10:42" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3480" daytime="10:42" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3481" daytime="10:44" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1141" daytime="10:46" gender="M" number="30" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1142" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1388" />
                    <RANKING order="2" place="2" resultid="2311" />
                    <RANKING order="3" place="3" resultid="1603" />
                    <RANKING order="4" place="4" resultid="3275" />
                    <RANKING order="5" place="5" resultid="2326" />
                    <RANKING order="6" place="6" resultid="2165" />
                    <RANKING order="7" place="7" resultid="2285" />
                    <RANKING order="8" place="8" resultid="2275" />
                    <RANKING order="9" place="9" resultid="2300" />
                    <RANKING order="10" place="10" resultid="3208" />
                    <RANKING order="11" place="11" resultid="2220" />
                    <RANKING order="12" place="12" resultid="2495" />
                    <RANKING order="13" place="13" resultid="2234" />
                    <RANKING order="14" place="14" resultid="3262" />
                    <RANKING order="15" place="15" resultid="2257" />
                    <RANKING order="16" place="16" resultid="2825" />
                    <RANKING order="17" place="17" resultid="3254" />
                    <RANKING order="18" place="18" resultid="2321" />
                    <RANKING order="19" place="19" resultid="2331" />
                    <RANKING order="20" place="20" resultid="3270" />
                    <RANKING order="21" place="21" resultid="2922" />
                    <RANKING order="22" place="22" resultid="3337" />
                    <RANKING order="23" place="23" resultid="3239" />
                    <RANKING order="24" place="-1" resultid="2239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1143" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2104" />
                    <RANKING order="2" place="2" resultid="2114" />
                    <RANKING order="3" place="3" resultid="3171" />
                    <RANKING order="4" place="4" resultid="2094" />
                    <RANKING order="5" place="5" resultid="2139" />
                    <RANKING order="6" place="6" resultid="2069" />
                    <RANKING order="7" place="7" resultid="2134" />
                    <RANKING order="8" place="8" resultid="2881" />
                    <RANKING order="9" place="9" resultid="1647" />
                    <RANKING order="10" place="10" resultid="2089" />
                    <RANKING order="11" place="11" resultid="2064" />
                    <RANKING order="12" place="12" resultid="2074" />
                    <RANKING order="13" place="13" resultid="2149" />
                    <RANKING order="14" place="14" resultid="2109" />
                    <RANKING order="15" place="15" resultid="1499" />
                    <RANKING order="16" place="16" resultid="2341" />
                    <RANKING order="17" place="17" resultid="2099" />
                    <RANKING order="18" place="18" resultid="1592" />
                    <RANKING order="19" place="19" resultid="2160" />
                    <RANKING order="20" place="20" resultid="2316" />
                    <RANKING order="21" place="21" resultid="3361" />
                    <RANKING order="22" place="22" resultid="3293" />
                    <RANKING order="23" place="23" resultid="3248" />
                    <RANKING order="24" place="24" resultid="3314" />
                    <RANKING order="25" place="25" resultid="1517" />
                    <RANKING order="26" place="26" resultid="3350" />
                    <RANKING order="27" place="27" resultid="2290" />
                    <RANKING order="28" place="-1" resultid="3047" />
                    <RANKING order="29" place="-1" resultid="2224" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3482" daytime="10:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3483" daytime="10:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3484" daytime="10:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3485" daytime="10:52" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3486" daytime="10:54" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3487" daytime="10:56" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="3488" daytime="10:56" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-03-02" daytime="15:10" endtime="18:28" name="3ª Etapa (Infantil/Sênior)" number="3" officialmeeting="15:30" warmupfrom="14:00" warmupuntil="15:00">
          <EVENTS>
            <EVENT eventid="1144" daytime="15:10" gender="F" number="31" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1145" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2194" />
                    <RANKING order="2" place="2" resultid="2029" />
                    <RANKING order="3" place="3" resultid="2011" />
                    <RANKING order="4" place="4" resultid="1981" />
                    <RANKING order="5" place="5" resultid="2601" />
                    <RANKING order="6" place="6" resultid="2005" />
                    <RANKING order="7" place="7" resultid="2595" />
                    <RANKING order="8" place="8" resultid="2183" />
                    <RANKING order="9" place="9" resultid="2868" />
                    <RANKING order="10" place="10" resultid="1993" />
                    <RANKING order="11" place="11" resultid="3127" />
                    <RANKING order="12" place="12" resultid="3180" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1935" />
                    <RANKING order="2" place="2" resultid="1893" />
                    <RANKING order="3" place="3" resultid="1887" />
                    <RANKING order="4" place="4" resultid="1899" />
                    <RANKING order="5" place="5" resultid="1923" />
                    <RANKING order="6" place="6" resultid="3155" />
                    <RANKING order="7" place="7" resultid="1947" />
                    <RANKING order="8" place="8" resultid="1780" />
                    <RANKING order="9" place="9" resultid="3218" />
                    <RANKING order="10" place="10" resultid="3197" />
                    <RANKING order="11" place="11" resultid="2892" />
                    <RANKING order="12" place="12" resultid="1882" />
                    <RANKING order="13" place="13" resultid="2044" />
                    <RANKING order="14" place="14" resultid="2709" />
                    <RANKING order="15" place="15" resultid="1435" />
                    <RANKING order="16" place="16" resultid="3378" />
                    <RANKING order="17" place="17" resultid="2945" />
                    <RANKING order="18" place="18" resultid="2951" />
                    <RANKING order="19" place="-1" resultid="3382" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1730" />
                    <RANKING order="2" place="2" resultid="3061" />
                    <RANKING order="3" place="3" resultid="1777" />
                    <RANKING order="4" place="4" resultid="1851" />
                    <RANKING order="5" place="5" resultid="2775" />
                    <RANKING order="6" place="6" resultid="1669" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1148" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2836" />
                    <RANKING order="2" place="2" resultid="2977" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1149" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1793" />
                    <RANKING order="2" place="2" resultid="2808" />
                    <RANKING order="3" place="3" resultid="1615" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3075" />
                    <RANKING order="2" place="2" resultid="2873" />
                    <RANKING order="3" place="3" resultid="2930" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1151" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2414" />
                    <RANKING order="2" place="2" resultid="2590" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3489" daytime="15:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3490" daytime="15:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3491" daytime="15:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3492" daytime="15:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3493" daytime="15:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3494" daytime="15:48" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1152" daytime="15:54" gender="M" number="32" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1153" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1964" />
                    <RANKING order="2" place="2" resultid="2152" />
                    <RANKING order="3" place="3" resultid="1958" />
                    <RANKING order="4" place="4" resultid="1976" />
                    <RANKING order="5" place="5" resultid="2036" />
                    <RANKING order="6" place="6" resultid="2000" />
                    <RANKING order="7" place="7" resultid="3173" />
                    <RANKING order="8" place="8" resultid="3144" />
                    <RANKING order="9" place="9" resultid="1685" />
                    <RANKING order="10" place="10" resultid="3132" />
                    <RANKING order="11" place="11" resultid="2024" />
                    <RANKING order="12" place="12" resultid="2304" />
                    <RANKING order="13" place="13" resultid="3140" />
                    <RANKING order="14" place="14" resultid="2364" />
                    <RANKING order="15" place="15" resultid="2924" />
                    <RANKING order="16" place="16" resultid="3184" />
                    <RANKING order="17" place="-1" resultid="3330" />
                    <RANKING order="18" place="-1" resultid="3136" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1906" />
                    <RANKING order="2" place="2" resultid="2051" />
                    <RANKING order="3" place="3" resultid="1918" />
                    <RANKING order="4" place="4" resultid="1566" />
                    <RANKING order="5" place="5" resultid="1871" />
                    <RANKING order="6" place="6" resultid="1912" />
                    <RANKING order="7" place="7" resultid="3148" />
                    <RANKING order="8" place="8" resultid="1942" />
                    <RANKING order="9" place="9" resultid="1690" />
                    <RANKING order="10" place="-1" resultid="2854" />
                    <RANKING order="11" place="-1" resultid="1596" />
                    <RANKING order="12" place="-1" resultid="3283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1755" />
                    <RANKING order="2" place="2" resultid="1790" />
                    <RANKING order="3" place="3" resultid="2848" />
                    <RANKING order="4" place="4" resultid="1359" />
                    <RANKING order="5" place="5" resultid="3031" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2056" />
                    <RANKING order="2" place="2" resultid="2696" />
                    <RANKING order="3" place="3" resultid="2888" />
                    <RANKING order="4" place="4" resultid="1721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1796" />
                    <RANKING order="2" place="2" resultid="3070" />
                    <RANKING order="3" place="3" resultid="2972" />
                    <RANKING order="4" place="4" resultid="2917" />
                    <RANKING order="5" place="5" resultid="3375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2627" />
                    <RANKING order="2" place="2" resultid="2631" />
                    <RANKING order="3" place="3" resultid="3119" />
                    <RANKING order="4" place="4" resultid="2897" />
                    <RANKING order="5" place="5" resultid="2833" />
                    <RANKING order="6" place="6" resultid="1809" />
                    <RANKING order="7" place="7" resultid="2936" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2907" />
                    <RANKING order="2" place="2" resultid="1544" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3495" daytime="15:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3496" daytime="16:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3497" daytime="16:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3498" daytime="16:16" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3499" daytime="16:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3500" daytime="16:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="3501" daytime="16:36" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1160" daytime="16:42" gender="F" number="33" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1161" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2195" />
                    <RANKING order="2" place="2" resultid="2602" />
                    <RANKING order="3" place="3" resultid="2007" />
                    <RANKING order="4" place="4" resultid="1983" />
                    <RANKING order="5" place="5" resultid="2185" />
                    <RANKING order="6" place="6" resultid="2031" />
                    <RANKING order="7" place="7" resultid="2803" />
                    <RANKING order="8" place="8" resultid="1994" />
                    <RANKING order="9" place="9" resultid="2013" />
                    <RANKING order="10" place="10" resultid="3129" />
                    <RANKING order="11" place="11" resultid="2760" />
                    <RANKING order="12" place="12" resultid="2597" />
                    <RANKING order="13" place="13" resultid="1480" />
                    <RANKING order="14" place="14" resultid="3340" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1162" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2399" />
                    <RANKING order="2" place="2" resultid="1782" />
                    <RANKING order="3" place="3" resultid="2711" />
                    <RANKING order="4" place="4" resultid="2178" />
                    <RANKING order="5" place="5" resultid="1884" />
                    <RANKING order="6" place="6" resultid="1369" />
                    <RANKING order="7" place="7" resultid="1381" />
                    <RANKING order="8" place="8" resultid="3029" />
                    <RANKING order="9" place="-1" resultid="1936" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1163" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1576" />
                    <RANKING order="2" place="2" resultid="1839" />
                    <RANKING order="3" place="3" resultid="1843" />
                    <RANKING order="4" place="4" resultid="1786" />
                    <RANKING order="5" place="5" resultid="1352" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1164" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1726" />
                    <RANKING order="2" place="2" resultid="2190" />
                    <RANKING order="3" place="3" resultid="2979" />
                    <RANKING order="4" place="4" resultid="1446" />
                    <RANKING order="5" place="-1" resultid="3084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1766" />
                    <RANKING order="2" place="2" resultid="1611" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2623" />
                    <RANKING order="2" place="2" resultid="1338" />
                    <RANKING order="3" place="3" resultid="2743" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2591" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3502" daytime="16:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3503" daytime="16:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3504" daytime="16:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3505" daytime="16:52" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3506" daytime="16:54" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1168" daytime="16:56" gender="M" number="34" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1169" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2017" />
                    <RANKING order="2" place="2" resultid="1970" />
                    <RANKING order="3" place="3" resultid="2035" />
                    <RANKING order="4" place="4" resultid="3143" />
                    <RANKING order="5" place="5" resultid="3139" />
                    <RANKING order="6" place="6" resultid="2303" />
                    <RANKING order="7" place="7" resultid="1988" />
                    <RANKING order="8" place="8" resultid="1605" />
                    <RANKING order="9" place="9" resultid="3012" />
                    <RANKING order="10" place="-1" resultid="3342" />
                    <RANKING order="11" place="-1" resultid="3135" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1565" />
                    <RANKING order="2" place="2" resultid="2409" />
                    <RANKING order="3" place="3" resultid="1929" />
                    <RANKING order="4" place="4" resultid="1870" />
                    <RANKING order="5" place="5" resultid="1905" />
                    <RANKING order="6" place="6" resultid="2853" />
                    <RANKING order="7" place="7" resultid="1877" />
                    <RANKING order="8" place="8" resultid="3023" />
                    <RANKING order="9" place="-1" resultid="1595" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1329" />
                    <RANKING order="2" place="2" resultid="2863" />
                    <RANKING order="3" place="3" resultid="3287" />
                    <RANKING order="4" place="4" resultid="1834" />
                    <RANKING order="5" place="5" resultid="1847" />
                    <RANKING order="6" place="6" resultid="3113" />
                    <RANKING order="7" place="7" resultid="1554" />
                    <RANKING order="8" place="8" resultid="1624" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1763" />
                    <RANKING order="2" place="2" resultid="1752" />
                    <RANKING order="3" place="3" resultid="2358" />
                    <RANKING order="4" place="4" resultid="2246" />
                    <RANKING order="5" place="5" resultid="1825" />
                    <RANKING order="6" place="6" resultid="1817" />
                    <RANKING order="7" place="7" resultid="2695" />
                    <RANKING order="8" place="8" resultid="2887" />
                    <RANKING order="9" place="9" resultid="2739" />
                    <RANKING order="10" place="10" resultid="1694" />
                    <RANKING order="11" place="11" resultid="1460" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1173" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1800" />
                    <RANKING order="2" place="2" resultid="3088" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1770" />
                    <RANKING order="2" place="2" resultid="1744" />
                    <RANKING order="3" place="3" resultid="3159" />
                    <RANKING order="4" place="4" resultid="2828" />
                    <RANKING order="5" place="5" resultid="2935" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1804" />
                    <RANKING order="2" place="2" resultid="1866" />
                    <RANKING order="3" place="3" resultid="3616" />
                    <RANKING order="4" place="4" resultid="1334" />
                    <RANKING order="5" place="5" resultid="1547" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3507" daytime="16:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3508" daytime="17:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3509" daytime="17:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3510" daytime="17:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3511" daytime="17:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3512" daytime="17:10" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="3513" daytime="17:14" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1176" daytime="17:16" gender="F" number="35" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1177" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1399" />
                    <RANKING order="2" place="-1" resultid="1471" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3368" />
                    <RANKING order="2" place="2" resultid="3156" />
                    <RANKING order="3" place="3" resultid="2953" />
                    <RANKING order="4" place="4" resultid="3379" />
                    <RANKING order="5" place="5" resultid="2947" />
                    <RANKING order="6" place="-1" resultid="3383" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1179" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1739" />
                    <RANKING order="2" place="2" resultid="1581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1180" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1734" />
                    <RANKING order="2" place="2" resultid="1441" />
                    <RANKING order="3" place="3" resultid="1466" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1181" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1610" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3076" />
                    <RANKING order="2" place="2" resultid="1337" />
                    <RANKING order="3" place="3" resultid="2883" />
                    <RANKING order="4" place="4" resultid="2931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1183" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3117" />
                    <RANKING order="2" place="2" resultid="2941" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3514" daytime="17:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3515" daytime="17:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3516" daytime="17:20" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1184" daytime="17:22" gender="M" number="36" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1185" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1684" />
                    <RANKING order="2" place="2" resultid="3329" />
                    <RANKING order="3" place="3" resultid="1559" />
                    <RANKING order="4" place="4" resultid="2968" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3147" />
                    <RANKING order="2" place="2" resultid="2050" />
                    <RANKING order="3" place="3" resultid="1941" />
                    <RANKING order="4" place="4" resultid="3022" />
                    <RANKING order="5" place="-1" resultid="1594" />
                    <RANKING order="6" place="-1" resultid="1689" />
                    <RANKING order="7" place="-1" resultid="3282" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1328" />
                    <RANKING order="2" place="2" resultid="3092" />
                    <RANKING order="3" place="3" resultid="2619" />
                    <RANKING order="4" place="4" resultid="1356" />
                    <RANKING order="5" place="5" resultid="3371" />
                    <RANKING order="6" place="6" resultid="1856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1188" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1759" />
                    <RANKING order="2" place="2" resultid="1820" />
                    <RANKING order="3" place="3" resultid="2417" />
                    <RANKING order="4" place="4" resultid="3079" />
                    <RANKING order="5" place="5" resultid="3105" />
                    <RANKING order="6" place="6" resultid="2750" />
                    <RANKING order="7" place="7" resultid="1451" />
                    <RANKING order="8" place="8" resultid="1824" />
                    <RANKING order="9" place="9" resultid="1650" />
                    <RANKING order="10" place="10" resultid="3049" />
                    <RANKING order="11" place="11" resultid="1633" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1189" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2842" />
                    <RANKING order="2" place="2" resultid="3087" />
                    <RANKING order="3" place="3" resultid="3041" />
                    <RANKING order="4" place="4" resultid="3006" />
                    <RANKING order="5" place="5" resultid="2916" />
                    <RANKING order="6" place="6" resultid="2792" />
                    <RANKING order="7" place="7" resultid="1708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1953" />
                    <RANKING order="2" place="2" resultid="3163" />
                    <RANKING order="3" place="3" resultid="1363" />
                    <RANKING order="4" place="4" resultid="1539" />
                    <RANKING order="5" place="5" resultid="1673" />
                    <RANKING order="6" place="6" resultid="1700" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2403" />
                    <RANKING order="2" place="2" resultid="1550" />
                    <RANKING order="3" place="3" resultid="2906" />
                    <RANKING order="4" place="4" resultid="1535" />
                    <RANKING order="5" place="5" resultid="1543" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3517" daytime="17:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3518" daytime="17:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3519" daytime="17:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3520" daytime="17:28" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3521" daytime="17:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3522" daytime="17:30" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1192" daytime="17:32" gender="F" number="37" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1193" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2030" />
                    <RANKING order="2" place="2" resultid="2012" />
                    <RANKING order="3" place="3" resultid="2184" />
                    <RANKING order="4" place="4" resultid="1982" />
                    <RANKING order="5" place="5" resultid="2596" />
                    <RANKING order="6" place="6" resultid="2006" />
                    <RANKING order="7" place="7" resultid="1658" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1456" />
                    <RANKING order="2" place="2" resultid="1894" />
                    <RANKING order="3" place="3" resultid="1883" />
                    <RANKING order="4" place="4" resultid="1901" />
                    <RANKING order="5" place="5" resultid="2710" />
                    <RANKING order="6" place="6" resultid="1925" />
                    <RANKING order="7" place="7" resultid="2893" />
                    <RANKING order="8" place="8" resultid="2398" />
                    <RANKING order="9" place="9" resultid="2177" />
                    <RANKING order="10" place="10" resultid="1948" />
                    <RANKING order="11" place="11" resultid="2946" />
                    <RANKING order="12" place="12" resultid="3028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1195" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1521" />
                    <RANKING order="2" place="2" resultid="1343" />
                    <RANKING order="3" place="3" resultid="1852" />
                    <RANKING order="4" place="4" resultid="2989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1196" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1733" />
                    <RANKING order="2" place="2" resultid="3152" />
                    <RANKING order="3" place="3" resultid="2837" />
                    <RANKING order="4" place="4" resultid="2912" />
                    <RANKING order="5" place="5" resultid="2958" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1197" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3066" />
                    <RANKING order="2" place="2" resultid="1348" />
                    <RANKING order="3" place="3" resultid="2810" />
                    <RANKING order="4" place="4" resultid="1616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1431" />
                    <RANKING order="2" place="2" resultid="2874" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1199" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3523" daytime="17:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3524" daytime="17:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3525" daytime="17:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3526" daytime="17:42" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3527" daytime="17:46" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1200" daytime="17:48" gender="M" number="38" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1201" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2151" />
                    <RANKING order="2" place="2" resultid="1492" />
                    <RANKING order="3" place="3" resultid="3131" />
                    <RANKING order="4" place="4" resultid="1374" />
                    <RANKING order="5" place="5" resultid="2023" />
                    <RANKING order="6" place="6" resultid="1963" />
                    <RANKING order="7" place="7" resultid="1975" />
                    <RANKING order="8" place="8" resultid="1957" />
                    <RANKING order="9" place="9" resultid="1969" />
                    <RANKING order="10" place="10" resultid="1999" />
                    <RANKING order="11" place="11" resultid="2302" />
                    <RANKING order="12" place="12" resultid="2816" />
                    <RANKING order="13" place="13" resultid="1987" />
                    <RANKING order="14" place="14" resultid="2363" />
                    <RANKING order="15" place="15" resultid="2967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2408" />
                    <RANKING order="2" place="2" resultid="1564" />
                    <RANKING order="3" place="3" resultid="1911" />
                    <RANKING order="4" place="4" resultid="1876" />
                    <RANKING order="5" place="5" resultid="1917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1203" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1524" />
                    <RANKING order="2" place="2" resultid="1322" />
                    <RANKING order="3" place="3" resultid="3286" />
                    <RANKING order="4" place="4" resultid="3097" />
                    <RANKING order="5" place="5" resultid="2862" />
                    <RANKING order="6" place="6" resultid="1859" />
                    <RANKING order="7" place="-1" resultid="2847" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1204" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1747" />
                    <RANKING order="2" place="2" resultid="1862" />
                    <RANKING order="3" place="3" resultid="1828" />
                    <RANKING order="4" place="4" resultid="1751" />
                    <RANKING order="5" place="5" resultid="1816" />
                    <RANKING order="6" place="6" resultid="1812" />
                    <RANKING order="7" place="7" resultid="1450" />
                    <RANKING order="8" place="8" resultid="1649" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1205" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2691" />
                    <RANKING order="2" place="2" resultid="2786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1206" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1743" />
                    <RANKING order="2" place="2" resultid="1808" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3528" daytime="17:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3529" daytime="17:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3530" daytime="17:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3531" daytime="17:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3532" daytime="18:02" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1208" daytime="18:04" gender="F" number="39" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1209" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1398" />
                    <RANKING order="2" place="2" resultid="2802" />
                    <RANKING order="3" place="3" resultid="1679" />
                    <RANKING order="4" place="4" resultid="2869" />
                    <RANKING order="5" place="5" resultid="3128" />
                    <RANKING order="6" place="6" resultid="3181" />
                    <RANKING order="7" place="7" resultid="2759" />
                    <RANKING order="8" place="8" resultid="1657" />
                    <RANKING order="9" place="9" resultid="1470" />
                    <RANKING order="10" place="10" resultid="1479" />
                    <RANKING order="11" place="11" resultid="1511" />
                    <RANKING order="12" place="12" resultid="3357" />
                    <RANKING order="13" place="13" resultid="2992" />
                    <RANKING order="14" place="14" resultid="3339" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1210" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1888" />
                    <RANKING order="2" place="2" resultid="1455" />
                    <RANKING order="3" place="3" resultid="2397" />
                    <RANKING order="4" place="4" resultid="1781" />
                    <RANKING order="5" place="5" resultid="1900" />
                    <RANKING order="6" place="6" resultid="2045" />
                    <RANKING order="7" place="7" resultid="3198" />
                    <RANKING order="8" place="8" resultid="1924" />
                    <RANKING order="9" place="9" resultid="1436" />
                    <RANKING order="10" place="10" resultid="1380" />
                    <RANKING order="11" place="11" resultid="2952" />
                    <RANKING order="12" place="12" resultid="1368" />
                    <RANKING order="13" place="13" resultid="2766" />
                    <RANKING order="14" place="14" resultid="1505" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1738" />
                    <RANKING order="2" place="2" resultid="1342" />
                    <RANKING order="3" place="3" resultid="2776" />
                    <RANKING order="4" place="4" resultid="3109" />
                    <RANKING order="5" place="5" resultid="1520" />
                    <RANKING order="6" place="6" resultid="1580" />
                    <RANKING order="7" place="7" resultid="3101" />
                    <RANKING order="8" place="8" resultid="3123" />
                    <RANKING order="9" place="9" resultid="1575" />
                    <RANKING order="10" place="10" resultid="1670" />
                    <RANKING order="11" place="11" resultid="2988" />
                    <RANKING order="12" place="12" resultid="2755" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1212" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2978" />
                    <RANKING order="2" place="2" resultid="2189" />
                    <RANKING order="3" place="3" resultid="1440" />
                    <RANKING order="4" place="4" resultid="1445" />
                    <RANKING order="5" place="5" resultid="3083" />
                    <RANKING order="6" place="6" resultid="3151" />
                    <RANKING order="7" place="7" resultid="2957" />
                    <RANKING order="8" place="8" resultid="2769" />
                    <RANKING order="9" place="9" resultid="1465" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1213" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3065" />
                    <RANKING order="2" place="2" resultid="1347" />
                    <RANKING order="3" place="3" resultid="2809" />
                    <RANKING order="4" place="4" resultid="1609" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1430" />
                    <RANKING order="2" place="2" resultid="2742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2940" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3533" daytime="18:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3534" daytime="18:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3535" daytime="18:08" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3536" daytime="18:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3537" daytime="18:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3538" daytime="18:12" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="3539" daytime="18:14" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1216" daytime="18:16" gender="M" number="40" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1217" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2153" />
                    <RANKING order="2" place="2" resultid="3174" />
                    <RANKING order="3" place="3" resultid="1686" />
                    <RANKING order="4" place="4" resultid="2018" />
                    <RANKING order="5" place="5" resultid="1375" />
                    <RANKING order="6" place="6" resultid="1971" />
                    <RANKING order="7" place="7" resultid="3145" />
                    <RANKING order="8" place="8" resultid="2025" />
                    <RANKING order="9" place="9" resultid="2365" />
                    <RANKING order="10" place="10" resultid="3331" />
                    <RANKING order="11" place="11" resultid="1977" />
                    <RANKING order="12" place="12" resultid="1606" />
                    <RANKING order="13" place="13" resultid="2925" />
                    <RANKING order="14" place="14" resultid="1560" />
                    <RANKING order="15" place="15" resultid="3013" />
                    <RANKING order="16" place="16" resultid="1620" />
                    <RANKING order="17" place="17" resultid="2817" />
                    <RANKING order="18" place="18" resultid="1711" />
                    <RANKING order="19" place="19" resultid="1493" />
                    <RANKING order="20" place="20" resultid="3343" />
                    <RANKING order="21" place="-1" resultid="3137" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2410" />
                    <RANKING order="2" place="2" resultid="1872" />
                    <RANKING order="3" place="3" resultid="2052" />
                    <RANKING order="4" place="4" resultid="1930" />
                    <RANKING order="5" place="5" resultid="1907" />
                    <RANKING order="6" place="6" resultid="1629" />
                    <RANKING order="7" place="7" resultid="3024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1756" />
                    <RANKING order="2" place="2" resultid="1570" />
                    <RANKING order="3" place="3" resultid="1525" />
                    <RANKING order="4" place="4" resultid="1323" />
                    <RANKING order="5" place="5" resultid="2620" />
                    <RANKING order="6" place="6" resultid="1835" />
                    <RANKING order="7" place="7" resultid="3098" />
                    <RANKING order="8" place="8" resultid="3093" />
                    <RANKING order="9" place="9" resultid="3114" />
                    <RANKING order="10" place="10" resultid="1357" />
                    <RANKING order="11" place="11" resultid="1555" />
                    <RANKING order="12" place="12" resultid="3288" />
                    <RANKING order="13" place="13" resultid="1360" />
                    <RANKING order="14" place="14" resultid="1625" />
                    <RANKING order="15" place="15" resultid="3372" />
                    <RANKING order="16" place="16" resultid="3032" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1220" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2607" />
                    <RANKING order="2" place="2" resultid="2057" />
                    <RANKING order="3" place="3" resultid="2394" />
                    <RANKING order="4" place="4" resultid="1821" />
                    <RANKING order="5" place="5" resultid="3106" />
                    <RANKING order="6" place="6" resultid="2697" />
                    <RANKING order="7" place="7" resultid="1829" />
                    <RANKING order="8" place="8" resultid="2751" />
                    <RANKING order="9" place="9" resultid="3080" />
                    <RANKING order="10" place="10" resultid="2359" />
                    <RANKING order="11" place="11" resultid="1722" />
                    <RANKING order="12" place="12" resultid="1634" />
                    <RANKING order="13" place="13" resultid="1695" />
                    <RANKING order="14" place="14" resultid="3050" />
                    <RANKING order="15" place="15" resultid="1461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1221" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1797" />
                    <RANKING order="2" place="2" resultid="3071" />
                    <RANKING order="3" place="3" resultid="2843" />
                    <RANKING order="4" place="4" resultid="2973" />
                    <RANKING order="5" place="5" resultid="2787" />
                    <RANKING order="6" place="6" resultid="3007" />
                    <RANKING order="7" place="7" resultid="2793" />
                    <RANKING order="8" place="8" resultid="3042" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1222" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3614" />
                    <RANKING order="2" place="2" resultid="1771" />
                    <RANKING order="3" place="3" resultid="1529" />
                    <RANKING order="4" place="4" resultid="2898" />
                    <RANKING order="5" place="5" resultid="3164" />
                    <RANKING order="6" place="6" resultid="1364" />
                    <RANKING order="7" place="7" resultid="1540" />
                    <RANKING order="8" place="8" resultid="1701" />
                    <RANKING order="9" place="9" resultid="1674" />
                    <RANKING order="10" place="10" resultid="2829" />
                    <RANKING order="11" place="11" resultid="2747" />
                    <RANKING order="12" place="12" resultid="1418" />
                    <RANKING order="13" place="13" resultid="1810" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1223" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2404" />
                    <RANKING order="2" place="2" resultid="1532" />
                    <RANKING order="3" place="3" resultid="1551" />
                    <RANKING order="4" place="4" resultid="2908" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3540" daytime="18:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3541" daytime="18:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3542" daytime="18:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3543" daytime="18:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3544" daytime="18:22" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3545" daytime="18:24" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="3546" daytime="18:26" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="3547" daytime="18:28" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="3548" daytime="18:28" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="3549" daytime="18:30" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="3550" daytime="18:32" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-03-03" daytime="08:40" endtime="12:46" name="4ª Etapa (Infantil/Sênior)" number="4" officialmeeting="08:00" warmupfrom="07:30" warmupuntil="08:30">
          <EVENTS>
            <EVENT eventid="1224" daytime="08:40" gender="F" number="41" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1225" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2196" />
                    <RANKING order="2" place="2" resultid="2032" />
                    <RANKING order="3" place="3" resultid="1984" />
                    <RANKING order="4" place="4" resultid="2603" />
                    <RANKING order="5" place="5" resultid="2014" />
                    <RANKING order="6" place="6" resultid="2186" />
                    <RANKING order="7" place="7" resultid="2008" />
                    <RANKING order="8" place="8" resultid="2598" />
                    <RANKING order="9" place="9" resultid="1995" />
                    <RANKING order="10" place="-1" resultid="2804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1226" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1937" />
                    <RANKING order="2" place="2" resultid="1783" />
                    <RANKING order="3" place="3" resultid="2400" />
                    <RANKING order="4" place="4" resultid="1889" />
                    <RANKING order="5" place="5" resultid="2894" />
                    <RANKING order="6" place="6" resultid="1895" />
                    <RANKING order="7" place="7" resultid="2046" />
                    <RANKING order="8" place="7" resultid="2712" />
                    <RANKING order="9" place="9" resultid="1926" />
                    <RANKING order="10" place="10" resultid="1949" />
                    <RANKING order="11" place="-1" resultid="3219" />
                    <RANKING order="12" place="-1" resultid="2179" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1227" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1853" />
                    <RANKING order="2" place="2" resultid="1731" />
                    <RANKING order="3" place="3" resultid="1844" />
                    <RANKING order="4" place="4" resultid="1840" />
                    <RANKING order="5" place="5" resultid="1577" />
                    <RANKING order="6" place="-1" resultid="2777" />
                    <RANKING order="7" place="-1" resultid="1353" />
                    <RANKING order="8" place="-1" resultid="1787" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1228" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1727" />
                    <RANKING order="2" place="2" resultid="2611" />
                    <RANKING order="3" place="3" resultid="2838" />
                    <RANKING order="4" place="-1" resultid="1447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1229" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1767" />
                    <RANKING order="2" place="2" resultid="2811" />
                    <RANKING order="3" place="3" resultid="1612" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2624" />
                    <RANKING order="2" place="2" resultid="1339" />
                    <RANKING order="3" place="3" resultid="2875" />
                    <RANKING order="4" place="4" resultid="2884" />
                    <RANKING order="5" place="-1" resultid="2932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1231" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="2592" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3551" daytime="08:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3552" daytime="08:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3553" daytime="08:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3554" daytime="08:54" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3555" daytime="08:58" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3556" daytime="09:02" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1232" daytime="09:06" gender="M" number="42" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1233" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2037" />
                    <RANKING order="2" place="2" resultid="2019" />
                    <RANKING order="3" place="3" resultid="1959" />
                    <RANKING order="4" place="4" resultid="2001" />
                    <RANKING order="5" place="5" resultid="2026" />
                    <RANKING order="6" place="6" resultid="1989" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1234" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1567" />
                    <RANKING order="2" place="2" resultid="1908" />
                    <RANKING order="3" place="3" resultid="2411" />
                    <RANKING order="4" place="4" resultid="1913" />
                    <RANKING order="5" place="5" resultid="1931" />
                    <RANKING order="6" place="6" resultid="1919" />
                    <RANKING order="7" place="7" resultid="1943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1235" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1526" />
                    <RANKING order="2" place="2" resultid="1330" />
                    <RANKING order="3" place="3" resultid="2849" />
                    <RANKING order="4" place="4" resultid="1836" />
                    <RANKING order="5" place="5" resultid="1848" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1236" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1863" />
                    <RANKING order="2" place="2" resultid="1818" />
                    <RANKING order="3" place="3" resultid="1813" />
                    <RANKING order="4" place="4" resultid="2247" />
                    <RANKING order="5" place="5" resultid="2889" />
                    <RANKING order="6" place="6" resultid="1452" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1237" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1801" />
                    <RANKING order="2" place="2" resultid="3089" />
                    <RANKING order="3" place="3" resultid="2918" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1238" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1772" />
                    <RANKING order="2" place="2" resultid="1745" />
                    <RANKING order="3" place="3" resultid="1675" />
                    <RANKING order="4" place="4" resultid="2937" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1239" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1867" />
                    <RANKING order="2" place="2" resultid="1533" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3557" daytime="09:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3558" daytime="09:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3559" daytime="09:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3560" daytime="09:18" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3561" daytime="09:22" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1240" daytime="09:26" gender="F" number="43" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1241" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2198" />
                    <RANKING order="2" place="2" resultid="2033" />
                    <RANKING order="3" place="3" resultid="2015" />
                    <RANKING order="4" place="4" resultid="2605" />
                    <RANKING order="5" place="5" resultid="1401" />
                    <RANKING order="6" place="6" resultid="1985" />
                    <RANKING order="7" place="7" resultid="2009" />
                    <RANKING order="8" place="8" resultid="1682" />
                    <RANKING order="9" place="9" resultid="2187" />
                    <RANKING order="10" place="10" resultid="2806" />
                    <RANKING order="11" place="11" resultid="2599" />
                    <RANKING order="12" place="12" resultid="2871" />
                    <RANKING order="13" place="13" resultid="1997" />
                    <RANKING order="14" place="14" resultid="1660" />
                    <RANKING order="15" place="15" resultid="1473" />
                    <RANKING order="16" place="16" resultid="1482" />
                    <RANKING order="17" place="17" resultid="3358" />
                    <RANKING order="18" place="-1" resultid="1513" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1242" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1458" />
                    <RANKING order="2" place="2" resultid="1784" />
                    <RANKING order="3" place="3" resultid="3369" />
                    <RANKING order="4" place="4" resultid="1897" />
                    <RANKING order="5" place="5" resultid="1891" />
                    <RANKING order="6" place="6" resultid="2401" />
                    <RANKING order="7" place="7" resultid="1903" />
                    <RANKING order="8" place="8" resultid="1939" />
                    <RANKING order="9" place="9" resultid="1885" />
                    <RANKING order="10" place="10" resultid="1927" />
                    <RANKING order="11" place="11" resultid="2048" />
                    <RANKING order="12" place="12" resultid="2713" />
                    <RANKING order="13" place="13" resultid="1438" />
                    <RANKING order="14" place="14" resultid="2181" />
                    <RANKING order="15" place="15" resultid="1951" />
                    <RANKING order="16" place="16" resultid="1383" />
                    <RANKING order="17" place="17" resultid="1372" />
                    <RANKING order="18" place="18" resultid="2955" />
                    <RANKING order="19" place="19" resultid="2949" />
                    <RANKING order="20" place="-1" resultid="3384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1243" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1741" />
                    <RANKING order="2" place="2" resultid="3063" />
                    <RANKING order="3" place="3" resultid="2779" />
                    <RANKING order="4" place="4" resultid="3178" />
                    <RANKING order="5" place="5" resultid="1854" />
                    <RANKING order="6" place="6" resultid="1345" />
                    <RANKING order="7" place="7" resultid="3111" />
                    <RANKING order="8" place="8" resultid="3103" />
                    <RANKING order="9" place="9" resultid="3125" />
                    <RANKING order="10" place="10" resultid="1583" />
                    <RANKING order="11" place="11" resultid="2990" />
                    <RANKING order="12" place="12" resultid="2757" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1244" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2192" />
                    <RANKING order="2" place="2" resultid="1443" />
                    <RANKING order="3" place="3" resultid="2981" />
                    <RANKING order="4" place="4" resultid="2914" />
                    <RANKING order="5" place="5" resultid="3085" />
                    <RANKING order="6" place="6" resultid="1639" />
                    <RANKING order="7" place="7" resultid="2960" />
                    <RANKING order="8" place="8" resultid="1468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1245" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1794" />
                    <RANKING order="2" place="2" resultid="1768" />
                    <RANKING order="3" place="3" resultid="1350" />
                    <RANKING order="4" place="4" resultid="1618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1433" />
                    <RANKING order="2" place="2" resultid="2745" />
                    <RANKING order="3" place="3" resultid="2933" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2943" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3562" daytime="09:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3563" daytime="09:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3564" daytime="09:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3565" daytime="09:34" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3566" daytime="09:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3567" daytime="09:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="3568" daytime="09:42" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="3569" daytime="09:44" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="3570" daytime="09:46" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1248" daytime="09:50" gender="M" number="44" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1249" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2155" />
                    <RANKING order="2" place="2" resultid="2021" />
                    <RANKING order="3" place="3" resultid="1973" />
                    <RANKING order="4" place="4" resultid="1967" />
                    <RANKING order="5" place="5" resultid="3175" />
                    <RANKING order="6" place="6" resultid="1687" />
                    <RANKING order="7" place="7" resultid="1495" />
                    <RANKING order="8" place="8" resultid="1378" />
                    <RANKING order="9" place="9" resultid="2039" />
                    <RANKING order="10" place="10" resultid="2367" />
                    <RANKING order="11" place="11" resultid="1979" />
                    <RANKING order="12" place="12" resultid="2306" />
                    <RANKING order="13" place="13" resultid="1991" />
                    <RANKING order="14" place="14" resultid="3015" />
                    <RANKING order="15" place="15" resultid="1562" />
                    <RANKING order="16" place="16" resultid="1622" />
                    <RANKING order="17" place="17" resultid="2819" />
                    <RANKING order="18" place="18" resultid="2970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1250" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2412" />
                    <RANKING order="2" place="2" resultid="2054" />
                    <RANKING order="3" place="3" resultid="1874" />
                    <RANKING order="4" place="4" resultid="1915" />
                    <RANKING order="5" place="5" resultid="1933" />
                    <RANKING order="6" place="6" resultid="1945" />
                    <RANKING order="7" place="7" resultid="1880" />
                    <RANKING order="8" place="8" resultid="1631" />
                    <RANKING order="9" place="9" resultid="3026" />
                    <RANKING order="10" place="10" resultid="2764" />
                    <RANKING order="11" place="11" resultid="2860" />
                    <RANKING order="12" place="-1" resultid="1598" />
                    <RANKING order="13" place="-1" resultid="3284" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1251" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1326" />
                    <RANKING order="2" place="2" resultid="1527" />
                    <RANKING order="3" place="3" resultid="1757" />
                    <RANKING order="4" place="4" resultid="1791" />
                    <RANKING order="5" place="5" resultid="1837" />
                    <RANKING order="6" place="6" resultid="1573" />
                    <RANKING order="7" place="7" resultid="3099" />
                    <RANKING order="8" place="8" resultid="3095" />
                    <RANKING order="9" place="9" resultid="3115" />
                    <RANKING order="10" place="10" resultid="1557" />
                    <RANKING order="11" place="11" resultid="1627" />
                    <RANKING order="12" place="12" resultid="3373" />
                    <RANKING order="13" place="13" resultid="1706" />
                    <RANKING order="14" place="14" resultid="3034" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1252" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2059" />
                    <RANKING order="2" place="2" resultid="1761" />
                    <RANKING order="3" place="3" resultid="2609" />
                    <RANKING order="4" place="4" resultid="2395" />
                    <RANKING order="5" place="5" resultid="3107" />
                    <RANKING order="6" place="6" resultid="1749" />
                    <RANKING order="7" place="7" resultid="1864" />
                    <RANKING order="8" place="8" resultid="2753" />
                    <RANKING order="9" place="9" resultid="3081" />
                    <RANKING order="10" place="10" resultid="2361" />
                    <RANKING order="11" place="11" resultid="1652" />
                    <RANKING order="12" place="12" resultid="1723" />
                    <RANKING order="13" place="13" resultid="3053" />
                    <RANKING order="14" place="14" resultid="1698" />
                    <RANKING order="15" place="15" resultid="1463" />
                    <RANKING order="16" place="-1" resultid="1636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1253" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1798" />
                    <RANKING order="2" place="2" resultid="3073" />
                    <RANKING order="3" place="3" resultid="2693" />
                    <RANKING order="4" place="4" resultid="2845" />
                    <RANKING order="5" place="5" resultid="2975" />
                    <RANKING order="6" place="6" resultid="2790" />
                    <RANKING order="7" place="7" resultid="3376" />
                    <RANKING order="8" place="8" resultid="3010" />
                    <RANKING order="9" place="9" resultid="3044" />
                    <RANKING order="10" place="10" resultid="2796" />
                    <RANKING order="11" place="11" resultid="1709" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1254" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2629" />
                    <RANKING order="2" place="2" resultid="3121" />
                    <RANKING order="3" place="3" resultid="1955" />
                    <RANKING order="4" place="4" resultid="2900" />
                    <RANKING order="5" place="5" resultid="3166" />
                    <RANKING order="6" place="6" resultid="3161" />
                    <RANKING order="7" place="7" resultid="1541" />
                    <RANKING order="8" place="8" resultid="1702" />
                    <RANKING order="9" place="9" resultid="2748" />
                    <RANKING order="10" place="10" resultid="2831" />
                    <RANKING order="11" place="11" resultid="2938" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1255" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1806" />
                    <RANKING order="2" place="2" resultid="2042" />
                    <RANKING order="3" place="3" resultid="2406" />
                    <RANKING order="4" place="4" resultid="1537" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3571" daytime="09:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3572" daytime="09:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3573" daytime="09:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3574" daytime="09:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3575" daytime="10:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3576" daytime="10:04" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="3577" daytime="10:06" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="3578" daytime="10:08" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="3579" daytime="10:10" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="3580" daytime="10:12" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="3581" daytime="10:14" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1256" daytime="10:16" gender="F" number="45" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1257" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1258" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1896" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1778" />
                    <RANKING order="2" place="2" resultid="3177" />
                    <RANKING order="3" place="3" resultid="3102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1260" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1261" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2812" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1262" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2200" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2415" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3582" daytime="10:16" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1264" daytime="10:36" gender="M" number="46" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1265" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1966" />
                    <RANKING order="2" place="2" resultid="1978" />
                    <RANKING order="3" place="3" resultid="1961" />
                    <RANKING order="4" place="4" resultid="2020" />
                    <RANKING order="5" place="5" resultid="1972" />
                    <RANKING order="6" place="6" resultid="2003" />
                    <RANKING order="7" place="7" resultid="2928" />
                    <RANKING order="8" place="8" resultid="3185" />
                    <RANKING order="9" place="9" resultid="2366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1921" />
                    <RANKING order="2" place="2" resultid="1879" />
                    <RANKING order="3" place="3" resultid="2856" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1267" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2851" />
                    <RANKING order="2" place="2" resultid="2866" />
                    <RANKING order="3" place="3" resultid="1860" />
                    <RANKING order="4" place="4" resultid="1361" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1268" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1269" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2974" />
                    <RANKING order="2" place="2" resultid="2920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1270" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1775" />
                    <RANKING order="2" place="2" resultid="2632" />
                    <RANKING order="3" place="3" resultid="2834" />
                    <RANKING order="4" place="4" resultid="1366" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1271" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2910" />
                    <RANKING order="2" place="2" resultid="1545" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3583" daytime="10:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3584" daytime="10:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3585" daytime="11:16" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1272" daytime="11:38" gender="F" number="47" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1273" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1400" />
                    <RANKING order="2" place="2" resultid="2870" />
                    <RANKING order="3" place="3" resultid="1659" />
                    <RANKING order="4" place="4" resultid="1681" />
                    <RANKING order="5" place="5" resultid="1512" />
                    <RANKING order="6" place="-1" resultid="2993" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1274" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1437" />
                    <RANKING order="2" place="2" resultid="1371" />
                    <RANKING order="3" place="3" resultid="3380" />
                    <RANKING order="4" place="4" resultid="2948" />
                    <RANKING order="5" place="5" resultid="1506" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1275" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1522" />
                    <RANKING order="2" place="2" resultid="1344" />
                    <RANKING order="3" place="3" resultid="1740" />
                    <RANKING order="4" place="4" resultid="3110" />
                    <RANKING order="5" place="5" resultid="3124" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1276" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2612" />
                    <RANKING order="2" place="2" resultid="1736" />
                    <RANKING order="3" place="3" resultid="3153" />
                    <RANKING order="4" place="4" resultid="2840" />
                    <RANKING order="5" place="5" resultid="1467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1277" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3068" />
                    <RANKING order="2" place="2" resultid="1349" />
                    <RANKING order="3" place="3" resultid="1617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1278" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1432" />
                    <RANKING order="2" place="2" resultid="2885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1279" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2942" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3586" daytime="11:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3587" daytime="11:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3588" daytime="11:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3589" daytime="11:46" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1280" daytime="11:48" gender="M" number="48" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1281" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1494" />
                    <RANKING order="2" place="2" resultid="3133" />
                    <RANKING order="3" place="3" resultid="2927" />
                    <RANKING order="4" place="4" resultid="2818" />
                    <RANKING order="5" place="5" resultid="1621" />
                    <RANKING order="6" place="-1" resultid="1377" />
                    <RANKING order="7" place="-1" resultid="2969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1282" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1914" />
                    <RANKING order="2" place="2" resultid="1878" />
                    <RANKING order="3" place="3" resultid="1630" />
                    <RANKING order="4" place="4" resultid="1692" />
                    <RANKING order="5" place="5" resultid="2859" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1283" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1325" />
                    <RANKING order="2" place="2" resultid="2865" />
                    <RANKING order="3" place="3" resultid="1572" />
                    <RANKING order="4" place="4" resultid="1332" />
                    <RANKING order="5" place="5" resultid="1626" />
                    <RANKING order="6" place="6" resultid="1705" />
                    <RANKING order="7" place="7" resultid="3033" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1284" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1831" />
                    <RANKING order="2" place="2" resultid="1814" />
                    <RANKING order="3" place="3" resultid="2752" />
                    <RANKING order="4" place="4" resultid="1697" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2692" />
                    <RANKING order="2" place="2" resultid="2789" />
                    <RANKING order="3" place="3" resultid="3009" />
                    <RANKING order="4" place="4" resultid="2795" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1286" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3120" />
                    <RANKING order="2" place="2" resultid="1677" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1287" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2041" />
                    <RANKING order="2" place="2" resultid="2405" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3590" daytime="11:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3591" daytime="11:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3592" daytime="11:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3593" daytime="11:56" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1288" daytime="11:58" gender="F" number="49" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1289" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2197" />
                    <RANKING order="2" place="2" resultid="2604" />
                    <RANKING order="3" place="3" resultid="1472" />
                    <RANKING order="4" place="4" resultid="1996" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1290" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3157" />
                    <RANKING order="2" place="2" resultid="1938" />
                    <RANKING order="3" place="3" resultid="1950" />
                    <RANKING order="4" place="4" resultid="1890" />
                    <RANKING order="5" place="5" resultid="2047" />
                    <RANKING order="6" place="6" resultid="2895" />
                    <RANKING order="7" place="7" resultid="1902" />
                    <RANKING order="8" place="8" resultid="2180" />
                    <RANKING order="9" place="9" resultid="2954" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1291" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3062" />
                    <RANKING order="2" place="2" resultid="2778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1735" />
                    <RANKING order="2" place="2" resultid="1442" />
                    <RANKING order="3" place="3" resultid="2980" />
                    <RANKING order="4" place="4" resultid="1638" />
                    <RANKING order="5" place="5" resultid="2839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1293" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1294" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3077" />
                    <RANKING order="2" place="2" resultid="2876" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1295" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2593" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3594" daytime="11:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3595" daytime="12:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3596" daytime="12:04" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1296" daytime="12:06" gender="M" number="50" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1297" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2154" />
                    <RANKING order="2" place="2" resultid="1965" />
                    <RANKING order="3" place="3" resultid="2002" />
                    <RANKING order="4" place="4" resultid="1960" />
                    <RANKING order="5" place="5" resultid="2038" />
                    <RANKING order="6" place="6" resultid="2305" />
                    <RANKING order="7" place="7" resultid="2027" />
                    <RANKING order="8" place="8" resultid="1990" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1298" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1568" />
                    <RANKING order="2" place="2" resultid="2053" />
                    <RANKING order="3" place="3" resultid="3149" />
                    <RANKING order="4" place="4" resultid="1909" />
                    <RANKING order="5" place="5" resultid="1932" />
                    <RANKING order="6" place="6" resultid="1944" />
                    <RANKING order="7" place="7" resultid="1920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1299" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2621" />
                    <RANKING order="2" place="2" resultid="3094" />
                    <RANKING order="3" place="3" resultid="1324" />
                    <RANKING order="4" place="4" resultid="2850" />
                    <RANKING order="5" place="5" resultid="1857" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1300" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1760" />
                    <RANKING order="2" place="2" resultid="2058" />
                    <RANKING order="3" place="3" resultid="1748" />
                    <RANKING order="4" place="4" resultid="1753" />
                    <RANKING order="5" place="5" resultid="2418" />
                    <RANKING order="6" place="6" resultid="1453" />
                    <RANKING order="7" place="7" resultid="1651" />
                    <RANKING order="8" place="8" resultid="3052" />
                    <RANKING order="9" place="-1" resultid="1822" />
                    <RANKING order="10" place="-1" resultid="1635" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1301" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1802" />
                    <RANKING order="2" place="2" resultid="3072" />
                    <RANKING order="3" place="3" resultid="2844" />
                    <RANKING order="4" place="4" resultid="3043" />
                    <RANKING order="5" place="-1" resultid="2794" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1302" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1954" />
                    <RANKING order="2" place="2" resultid="2628" />
                    <RANKING order="3" place="3" resultid="3165" />
                    <RANKING order="4" place="4" resultid="2899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1303" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1552" />
                    <RANKING order="2" place="2" resultid="1536" />
                    <RANKING order="3" place="3" resultid="2909" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3597" daytime="12:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3598" daytime="12:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3599" daytime="12:12" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3600" daytime="12:14" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3601" daytime="12:16" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3602" daytime="12:20" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1304" daytime="12:22" gender="F" number="51" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1305" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2805" />
                    <RANKING order="2" place="2" resultid="3182" />
                    <RANKING order="3" place="3" resultid="1680" />
                    <RANKING order="4" place="4" resultid="2761" />
                    <RANKING order="5" place="5" resultid="1481" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1306" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3199" />
                    <RANKING order="2" place="2" resultid="3220" />
                    <RANKING order="3" place="3" resultid="1457" />
                    <RANKING order="4" place="4" resultid="1382" />
                    <RANKING order="5" place="5" resultid="1370" />
                    <RANKING order="6" place="6" resultid="2767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1307" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1578" />
                    <RANKING order="2" place="2" resultid="1841" />
                    <RANKING order="3" place="3" resultid="1845" />
                    <RANKING order="4" place="4" resultid="1354" />
                    <RANKING order="5" place="5" resultid="1671" />
                    <RANKING order="6" place="6" resultid="1582" />
                    <RANKING order="7" place="7" resultid="2756" />
                    <RANKING order="8" place="-1" resultid="1788" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1308" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1728" />
                    <RANKING order="2" place="2" resultid="2191" />
                    <RANKING order="3" place="3" resultid="1448" />
                    <RANKING order="4" place="4" resultid="2913" />
                    <RANKING order="5" place="5" resultid="2959" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1309" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3067" />
                    <RANKING order="2" place="2" resultid="1613" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1310" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2625" />
                    <RANKING order="2" place="2" resultid="1340" />
                    <RANKING order="3" place="3" resultid="2744" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1311" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3603" daytime="12:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3604" daytime="12:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3605" daytime="12:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3606" daytime="12:28" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1312" daytime="12:30" gender="M" number="52" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1313" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3141" />
                    <RANKING order="2" place="2" resultid="1376" />
                    <RANKING order="3" place="3" resultid="3014" />
                    <RANKING order="4" place="4" resultid="1607" />
                    <RANKING order="5" place="5" resultid="1712" />
                    <RANKING order="6" place="6" resultid="2926" />
                    <RANKING order="7" place="-1" resultid="1561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1314" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1873" />
                    <RANKING order="2" place="2" resultid="3025" />
                    <RANKING order="3" place="3" resultid="2763" />
                    <RANKING order="4" place="4" resultid="1691" />
                    <RANKING order="5" place="-1" resultid="2855" />
                    <RANKING order="6" place="-1" resultid="2858" />
                    <RANKING order="7" place="-1" resultid="1597" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1315" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1331" />
                    <RANKING order="2" place="2" resultid="2864" />
                    <RANKING order="3" place="3" resultid="1571" />
                    <RANKING order="4" place="4" resultid="1849" />
                    <RANKING order="5" place="5" resultid="1556" />
                    <RANKING order="6" place="6" resultid="1704" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1316" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2608" />
                    <RANKING order="2" place="2" resultid="1764" />
                    <RANKING order="3" place="3" resultid="2360" />
                    <RANKING order="4" place="4" resultid="1826" />
                    <RANKING order="5" place="5" resultid="2890" />
                    <RANKING order="6" place="6" resultid="2740" />
                    <RANKING order="7" place="7" resultid="1830" />
                    <RANKING order="8" place="8" resultid="1696" />
                    <RANKING order="9" place="9" resultid="3051" />
                    <RANKING order="10" place="10" resultid="1462" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1317" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3090" />
                    <RANKING order="2" place="2" resultid="2919" />
                    <RANKING order="3" place="-1" resultid="2788" />
                    <RANKING order="4" place="-1" resultid="3008" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1318" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1530" />
                    <RANKING order="2" place="2" resultid="3160" />
                    <RANKING order="3" place="3" resultid="1365" />
                    <RANKING order="4" place="4" resultid="2830" />
                    <RANKING order="5" place="5" resultid="1676" />
                    <RANKING order="6" place="6" resultid="1419" />
                    <RANKING order="7" place="-1" resultid="1773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1319" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1805" />
                    <RANKING order="2" place="2" resultid="1868" />
                    <RANKING order="3" place="3" resultid="1335" />
                    <RANKING order="4" place="4" resultid="1548" />
                    <RANKING order="5" place="-1" resultid="3617" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="3607" daytime="12:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="3608" daytime="12:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="3609" daytime="12:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="3610" daytime="12:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="3611" daytime="12:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="3612" daytime="12:40" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="263" nation="BRA" region="PR" clubid="1724" swrid="75436" name="Clube Curitibano" shortname="Curitibano">
          <ATHLETES>
            <ATHLETE firstname="Betina" lastname="Vieira Pellanda" birthdate="2014-02-16" gender="F" nation="BRA" license="391041" swrid="5602589" athleteid="2486" externalid="391041">
              <RESULTS>
                <RESULT eventid="1092" points="124" swimtime="00:01:40.58" resultid="2487" heatid="3438" lane="6" entrytime="00:01:36.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="136" swimtime="00:00:49.00" resultid="2488" heatid="3419" lane="7" entrytime="00:00:52.40" entrycourse="SCM" />
                <RESULT eventid="1108" points="60" swimtime="00:01:01.99" resultid="2489" heatid="3455" lane="7" entrytime="00:01:00.01" entrycourse="SCM" />
                <RESULT eventid="1128" points="157" swimtime="00:00:42.42" resultid="2490" heatid="3469" lane="7" entrytime="00:00:44.77" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gael" lastname="Stramandinoli Zanicotti" birthdate="2015-03-21" gender="M" nation="BRA" license="406954" athleteid="2719" externalid="406954">
              <RESULTS>
                <RESULT eventid="1095" points="17" swimtime="00:02:52.13" resultid="2720" heatid="3441" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:19.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="35" swimtime="00:01:07.50" resultid="2721" heatid="3421" lane="8" />
                <RESULT eventid="1111" points="13" swimtime="00:01:31.38" resultid="2722" heatid="3457" lane="2" />
                <RESULT eventid="1131" points="28" swimtime="00:01:05.66" resultid="2723" heatid="3470" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="De Albuquerque" birthdate="2010-06-08" gender="F" nation="BRA" license="356249" swrid="5600145" athleteid="1881" externalid="356249">
              <RESULTS>
                <RESULT eventid="1144" points="344" swimtime="00:05:30.01" resultid="1882" heatid="3491" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:15.33" />
                    <SPLIT distance="150" swimtime="00:01:57.44" />
                    <SPLIT distance="200" swimtime="00:02:39.66" />
                    <SPLIT distance="250" swimtime="00:03:21.88" />
                    <SPLIT distance="300" swimtime="00:04:05.10" />
                    <SPLIT distance="350" swimtime="00:04:48.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="354" swimtime="00:01:17.58" resultid="1883" heatid="3527" lane="8" entrytime="00:01:14.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="257" swimtime="00:01:38.08" resultid="1884" heatid="3503" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="382" swimtime="00:01:09.23" resultid="1885" heatid="3562" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Cavalca Petraglia" birthdate="2015-08-06" gender="M" nation="BRA" license="397275" swrid="5641757" athleteid="2555" externalid="397275">
              <RESULTS>
                <RESULT eventid="1083" points="53" swimtime="00:00:58.56" resultid="2556" heatid="3422" lane="7" />
                <RESULT eventid="1071" points="57" swimtime="00:01:04.65" resultid="2557" heatid="3403" lane="3" entrytime="00:01:09.02" entrycourse="SCM" />
                <RESULT eventid="1111" points="58" swimtime="00:00:55.88" resultid="2558" heatid="3458" lane="3" entrytime="00:01:14.29" entrycourse="SCM" />
                <RESULT eventid="1131" points="52" swimtime="00:00:53.86" resultid="2559" heatid="3472" lane="6" entrytime="00:00:55.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Prosdocimo" birthdate="2012-11-30" gender="M" nation="BRA" license="369272" swrid="5602575" athleteid="2105" externalid="369272">
              <RESULTS>
                <RESULT eventid="1089" points="252" swimtime="00:02:37.19" resultid="2106" heatid="3434" lane="7" entrytime="00:02:43.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.30" />
                    <SPLIT distance="100" swimtime="00:01:16.91" />
                    <SPLIT distance="150" swimtime="00:01:57.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="195" reactiontime="+72" swimtime="00:00:38.07" resultid="2107" heatid="3415" lane="7" entrytime="00:00:40.51" entrycourse="SCM" />
                <RESULT eventid="1105" points="180" swimtime="00:01:27.22" resultid="2108" heatid="3448" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="219" swimtime="00:00:33.44" resultid="2109" heatid="3487" lane="8" entrytime="00:00:34.63" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorena" lastname="Mascarenhas" birthdate="2011-08-31" gender="F" nation="BRA" license="370581" swrid="5602558" athleteid="2182" externalid="370581">
              <RESULTS>
                <RESULT eventid="1144" points="324" swimtime="00:05:36.53" resultid="2183" heatid="3492" lane="4" entrytime="00:05:46.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.38" />
                    <SPLIT distance="100" swimtime="00:01:15.38" />
                    <SPLIT distance="150" swimtime="00:01:57.49" />
                    <SPLIT distance="200" swimtime="00:02:41.76" />
                    <SPLIT distance="250" swimtime="00:03:25.81" />
                    <SPLIT distance="300" swimtime="00:04:09.72" />
                    <SPLIT distance="350" swimtime="00:04:53.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="333" swimtime="00:01:19.14" resultid="2184" heatid="3525" lane="5" entrytime="00:01:23.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="312" swimtime="00:01:31.93" resultid="2185" heatid="3503" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="327" swimtime="00:02:56.82" resultid="2186" heatid="3554" lane="7" entrytime="00:03:05.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:24.41" />
                    <SPLIT distance="150" swimtime="00:02:15.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="349" swimtime="00:01:11.36" resultid="2187" heatid="3567" lane="8" entrytime="00:01:12.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Cabrini Vieira" birthdate="2012-02-11" gender="F" nation="BRA" license="376961" swrid="5588571" athleteid="2211" externalid="376961">
              <RESULTS>
                <RESULT eventid="1086" points="388" swimtime="00:02:31.16" resultid="2212" heatid="3428" lane="6" entrytime="00:02:40.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:14.67" />
                    <SPLIT distance="150" swimtime="00:01:52.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="330" swimtime="00:00:36.53" resultid="2213" heatid="3410" lane="5" entrytime="00:00:37.73" entrycourse="SCM" />
                <RESULT eventid="1102" points="308" swimtime="00:01:23.61" resultid="2214" heatid="3445" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="372" swimtime="00:00:31.88" resultid="2215" heatid="3481" lane="5" entrytime="00:00:32.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Trevisan" birthdate="2000-11-28" gender="M" nation="BRA" license="346847" swrid="5600266" athleteid="2402" externalid="346847">
              <RESULTS>
                <RESULT eventid="1184" points="574" swimtime="00:00:26.16" resultid="2403" heatid="3518" lane="1" />
                <RESULT eventid="1216" points="582" swimtime="00:00:24.14" resultid="2404" heatid="3550" lane="4" entrytime="00:00:23.93" entrycourse="SCM" />
                <RESULT eventid="1280" points="484" reactiontime="+58" swimtime="00:00:28.15" resultid="2405" heatid="3593" lane="3" entrytime="00:00:27.70" entrycourse="SCM" />
                <RESULT eventid="1248" points="591" swimtime="00:00:53.43" resultid="2406" heatid="3581" lane="2" entrytime="00:00:53.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diego" lastname="Rafael Navarchi Faria Vellozo" birthdate="2008-02-21" gender="M" nation="BRA" license="342231" swrid="5600239" athleteid="1827" externalid="342231">
              <RESULTS>
                <RESULT eventid="1200" points="415" reactiontime="+72" swimtime="00:01:04.79" resultid="1828" heatid="3532" lane="7" entrytime="00:01:07.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="409" swimtime="00:00:27.14" resultid="1829" heatid="3548" lane="5" entrytime="00:00:27.03" entrycourse="SCM" />
                <RESULT eventid="1312" points="308" swimtime="00:00:36.92" resultid="1830" heatid="3609" lane="1" />
                <RESULT eventid="1280" points="397" reactiontime="+52" swimtime="00:00:30.06" resultid="1831" heatid="3590" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Toscani Kim" birthdate="2015-10-02" gender="F" nation="BRA" license="397276" swrid="5641778" athleteid="2560" externalid="397276">
              <RESULTS>
                <RESULT eventid="1092" points="99" swimtime="00:01:48.33" resultid="2561" heatid="3436" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="122" swimtime="00:00:50.90" resultid="2562" heatid="3418" lane="7" />
                <RESULT eventid="1108" points="99" swimtime="00:00:52.60" resultid="2563" heatid="3452" lane="3" />
                <RESULT eventid="1128" points="114" swimtime="00:00:47.18" resultid="2564" heatid="3468" lane="8" entrytime="00:00:52.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Puppi Cardoso" birthdate="2015-03-30" gender="F" nation="BRA" license="406741" athleteid="2638" externalid="406741">
              <RESULTS>
                <RESULT eventid="1092" points="58" swimtime="00:02:09.78" resultid="2639" heatid="3435" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="90" reactiontime="+94" swimtime="00:00:56.23" resultid="2640" heatid="3416" lane="5" />
                <RESULT eventid="1108" points="39" swimtime="00:01:11.34" resultid="2641" heatid="3453" lane="2" />
                <RESULT eventid="1128" points="61" swimtime="00:00:58.19" resultid="2642" heatid="3467" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olavo" lastname="Valduga Artigas" birthdate="2012-06-26" gender="M" nation="BRA" license="369270" swrid="5588941" athleteid="2095" externalid="369270">
              <RESULTS>
                <RESULT eventid="1089" points="163" swimtime="00:03:01.81" resultid="2096" heatid="3432" lane="8" entrytime="00:03:10.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                    <SPLIT distance="100" swimtime="00:01:27.96" />
                    <SPLIT distance="150" swimtime="00:02:15.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="144" swimtime="00:01:45.29" resultid="2097" heatid="3398" lane="2" entrytime="00:01:42.05" entrycourse="SCM" />
                <RESULT eventid="1105" points="138" swimtime="00:01:35.23" resultid="2098" heatid="3449" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="171" swimtime="00:00:36.31" resultid="2099" heatid="3485" lane="4" entrytime="00:00:36.74" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Cristina Ferreira" birthdate="2011-08-24" gender="F" nation="BRA" license="358334" swrid="5588611" athleteid="2193" externalid="358334">
              <RESULTS>
                <RESULT eventid="1144" points="548" swimtime="00:04:42.63" resultid="2194" heatid="3494" lane="6" entrytime="00:04:40.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                    <SPLIT distance="100" swimtime="00:01:06.75" />
                    <SPLIT distance="150" swimtime="00:01:42.61" />
                    <SPLIT distance="200" swimtime="00:02:18.17" />
                    <SPLIT distance="250" swimtime="00:02:54.68" />
                    <SPLIT distance="300" swimtime="00:03:31.10" />
                    <SPLIT distance="350" swimtime="00:04:07.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="487" swimtime="00:01:19.22" resultid="2195" heatid="3506" lane="2" entrytime="00:01:21.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="510" swimtime="00:02:32.44" resultid="2196" heatid="3556" lane="5" entrytime="00:02:32.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="100" swimtime="00:01:12.51" />
                    <SPLIT distance="150" swimtime="00:01:58.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="594" swimtime="00:01:04.27" resultid="2197" heatid="3596" lane="4" entrytime="00:01:05.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="581" swimtime="00:01:00.19" resultid="2198" heatid="3563" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Fernandes Tramujas" birthdate="2015-01-15" gender="F" nation="BRA" license="406750" athleteid="2680" externalid="406750">
              <RESULTS>
                <RESULT eventid="1092" points="36" swimtime="00:02:31.88" resultid="2681" heatid="3436" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="57" swimtime="00:01:13.59" resultid="2682" heatid="3399" lane="3" />
                <RESULT eventid="1108" points="29" swimtime="00:01:18.61" resultid="2683" heatid="3453" lane="5" />
                <RESULT eventid="1128" status="DNS" swimtime="00:00:00.00" resultid="2684" heatid="3466" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Baptistella" birthdate="2013-01-23" gender="M" nation="BRA" license="391152" swrid="5602545" athleteid="2491" externalid="391152">
              <RESULTS>
                <RESULT eventid="1089" points="142" swimtime="00:03:10.42" resultid="2492" heatid="3432" lane="1" entrytime="00:03:08.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:01:29.96" />
                    <SPLIT distance="150" swimtime="00:02:21.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="140" reactiontime="+76" swimtime="00:00:42.53" resultid="2493" heatid="3414" lane="3" entrytime="00:00:41.56" entrycourse="SCM" />
                <RESULT eventid="1105" points="140" swimtime="00:01:34.88" resultid="2494" heatid="3451" lane="8" entrytime="00:01:43.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="160" swimtime="00:00:37.09" resultid="2495" heatid="3485" lane="5" entrytime="00:00:37.25" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Muxfeldt" birthdate="2011-05-13" gender="F" nation="BRA" license="366903" swrid="5602563" athleteid="2004" externalid="366903">
              <RESULTS>
                <RESULT eventid="1144" points="358" swimtime="00:05:25.53" resultid="2005" heatid="3492" lane="5" entrytime="00:06:03.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:14.38" />
                    <SPLIT distance="150" swimtime="00:01:56.11" />
                    <SPLIT distance="200" swimtime="00:02:38.08" />
                    <SPLIT distance="250" swimtime="00:03:20.32" />
                    <SPLIT distance="300" swimtime="00:04:03.34" />
                    <SPLIT distance="350" swimtime="00:04:46.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="276" reactiontime="+86" swimtime="00:01:24.22" resultid="2006" heatid="3524" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="340" swimtime="00:01:29.32" resultid="2007" heatid="3504" lane="6" entrytime="00:01:34.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="316" swimtime="00:02:58.75" resultid="2008" heatid="3552" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                    <SPLIT distance="100" swimtime="00:01:28.68" />
                    <SPLIT distance="150" swimtime="00:02:20.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="377" swimtime="00:01:09.53" resultid="2009" heatid="3566" lane="3" entrytime="00:01:14.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Iglesias Vargas" birthdate="2009-01-11" gender="M" nation="BRA" license="324792" swrid="5600189" athleteid="1789" externalid="324792">
              <RESULTS>
                <RESULT eventid="1152" points="502" swimtime="00:04:26.92" resultid="1790" heatid="3501" lane="2" entrytime="00:04:34.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.85" />
                    <SPLIT distance="100" swimtime="00:01:04.77" />
                    <SPLIT distance="150" swimtime="00:01:38.05" />
                    <SPLIT distance="200" swimtime="00:02:11.80" />
                    <SPLIT distance="250" swimtime="00:02:45.17" />
                    <SPLIT distance="300" swimtime="00:03:19.56" />
                    <SPLIT distance="350" swimtime="00:03:53.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="501" swimtime="00:00:56.45" resultid="1791" heatid="3572" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Felipe Paes Feres" birthdate="2008-07-28" gender="M" nation="BRA" license="307676" swrid="5600156" athleteid="1815" externalid="307676">
              <RESULTS>
                <RESULT eventid="1200" points="396" reactiontime="+62" swimtime="00:01:05.81" resultid="1816" heatid="3532" lane="2" entrytime="00:01:06.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="343" swimtime="00:01:18.90" resultid="1817" heatid="3509" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="412" swimtime="00:02:27.25" resultid="1818" heatid="3560" lane="4" entrytime="00:02:29.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                    <SPLIT distance="100" swimtime="00:01:09.66" />
                    <SPLIT distance="150" swimtime="00:01:54.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Kremer De Aguiar" birthdate="2009-12-22" gender="F" nation="BRA" license="338987" swrid="5600196" athleteid="1842" externalid="338987">
              <RESULTS>
                <RESULT eventid="1160" points="433" swimtime="00:01:22.41" resultid="1843" heatid="3505" lane="7" entrytime="00:01:28.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="393" swimtime="00:02:46.28" resultid="1844" heatid="3555" lane="2" entrytime="00:02:55.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="100" swimtime="00:01:21.52" />
                    <SPLIT distance="150" swimtime="00:02:08.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="421" swimtime="00:00:37.85" resultid="1845" heatid="3606" lane="1" entrytime="00:00:40.78" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nina" lastname="Rocha Ribeiro Da Silva" birthdate="2010-09-22" gender="F" nation="BRA" license="367216" swrid="5588884" athleteid="2396" externalid="367216">
              <RESULTS>
                <RESULT eventid="1208" points="414" swimtime="00:00:30.76" resultid="2397" heatid="3537" lane="4" entrytime="00:00:31.76" entrycourse="SCM" />
                <RESULT eventid="1192" points="271" reactiontime="+76" swimtime="00:01:24.82" resultid="2398" heatid="3524" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="472" swimtime="00:01:20.09" resultid="2399" heatid="3505" lane="2" entrytime="00:01:27.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="352" swimtime="00:02:52.45" resultid="2400" heatid="3554" lane="8" entrytime="00:03:06.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:23.58" />
                    <SPLIT distance="150" swimtime="00:02:10.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="414" swimtime="00:01:07.39" resultid="2401" heatid="3567" lane="6" entrytime="00:01:11.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Pacheco" birthdate="2012-10-13" gender="F" nation="BRA" license="376981" swrid="5602566" athleteid="2276" externalid="376981">
              <RESULTS>
                <RESULT eventid="1062" points="180" swimtime="00:01:50.44" resultid="2277" heatid="3394" lane="7" entrytime="00:02:02.94" entrycourse="SCM" />
                <RESULT eventid="1074" points="179" reactiontime="+77" swimtime="00:00:44.78" resultid="2278" heatid="3409" lane="1" entrytime="00:00:48.90" entrycourse="SCM" />
                <RESULT eventid="1102" points="162" swimtime="00:01:43.52" resultid="2279" heatid="3444" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="212" swimtime="00:00:38.44" resultid="2280" heatid="3479" lane="6" entrytime="00:00:41.08" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Simioni Albuquerque" birthdate="2014-12-23" gender="F" nation="BRA" license="401980" swrid="5661355" athleteid="2585" externalid="401980">
              <RESULTS>
                <RESULT eventid="1092" points="131" swimtime="00:01:38.92" resultid="2586" heatid="3437" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="114" reactiontime="+98" swimtime="00:00:51.93" resultid="2587" heatid="3418" lane="1" />
                <RESULT eventid="1108" points="119" swimtime="00:00:49.56" resultid="2588" heatid="3454" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Braun Prado" birthdate="2008-04-07" gender="M" nation="BRA" license="307663" swrid="5484324" athleteid="1861" externalid="307663">
              <RESULTS>
                <RESULT eventid="1200" points="472" reactiontime="+62" swimtime="00:01:02.06" resultid="1862" heatid="3532" lane="6" entrytime="00:01:03.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="439" swimtime="00:02:24.15" resultid="1863" heatid="3557" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                    <SPLIT distance="100" swimtime="00:01:06.32" />
                    <SPLIT distance="150" swimtime="00:01:50.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="469" swimtime="00:00:57.69" resultid="1864" heatid="3574" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Ribas Omar" birthdate="2014-11-28" gender="M" nation="BRA" license="406746" athleteid="2661" externalid="406746">
              <RESULTS>
                <RESULT eventid="1095" points="43" swimtime="00:02:07.50" resultid="2662" heatid="3440" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="60" swimtime="00:00:56.36" resultid="2663" heatid="3422" lane="8" />
                <RESULT eventid="1131" points="58" swimtime="00:00:51.97" resultid="2664" heatid="3471" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Alice Silva Gomes Xavier" birthdate="2013-02-25" gender="F" nation="BRA" license="371040" athleteid="2714" externalid="371040">
              <RESULTS>
                <RESULT eventid="1062" points="239" swimtime="00:01:40.35" resultid="2715" heatid="3393" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1086" points="284" swimtime="00:02:47.75" resultid="2716" heatid="3428" lane="8" entrytime="00:02:46.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:01:18.98" />
                    <SPLIT distance="150" swimtime="00:02:03.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1118" points="161" swimtime="00:01:39.23" resultid="2717" heatid="3462" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="299" swimtime="00:00:34.26" resultid="2718" heatid="3481" lane="8" entrytime="00:00:34.47" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Fontana" birthdate="2011-12-29" gender="M" nation="BRA" license="366897" swrid="5602539" athleteid="1986" externalid="366897">
              <RESULTS>
                <RESULT eventid="1200" points="160" swimtime="00:01:28.97" resultid="1987" heatid="3528" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="190" swimtime="00:01:36.06" resultid="1988" heatid="3510" lane="8" entrytime="00:01:47.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="192" swimtime="00:03:09.85" resultid="1989" heatid="3558" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.88" />
                    <SPLIT distance="100" swimtime="00:01:34.28" />
                    <SPLIT distance="150" swimtime="00:02:28.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="117" swimtime="00:01:37.58" resultid="1990" heatid="3598" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="206" swimtime="00:01:15.91" resultid="1991" heatid="3575" lane="5" entrytime="00:01:19.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Brandt De Macedo" birthdate="2006-04-22" gender="M" nation="BRA" license="296648" swrid="5622265" athleteid="1774" externalid="296648">
              <RESULTS>
                <RESULT eventid="1264" points="763" swimtime="00:15:26.71" resultid="1775" heatid="3583" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.74" />
                    <SPLIT distance="100" swimtime="00:00:57.85" />
                    <SPLIT distance="150" swimtime="00:01:28.51" />
                    <SPLIT distance="200" swimtime="00:01:59.09" />
                    <SPLIT distance="250" swimtime="00:02:30.02" />
                    <SPLIT distance="300" swimtime="00:03:00.84" />
                    <SPLIT distance="350" swimtime="00:03:31.91" />
                    <SPLIT distance="400" swimtime="00:04:02.93" />
                    <SPLIT distance="450" swimtime="00:04:33.99" />
                    <SPLIT distance="500" swimtime="00:05:05.08" />
                    <SPLIT distance="550" swimtime="00:05:35.55" />
                    <SPLIT distance="600" swimtime="00:06:06.54" />
                    <SPLIT distance="650" swimtime="00:06:37.65" />
                    <SPLIT distance="700" swimtime="00:07:09.01" />
                    <SPLIT distance="750" swimtime="00:07:40.45" />
                    <SPLIT distance="800" swimtime="00:08:11.56" />
                    <SPLIT distance="850" swimtime="00:08:42.75" />
                    <SPLIT distance="900" swimtime="00:09:14.23" />
                    <SPLIT distance="950" swimtime="00:09:45.83" />
                    <SPLIT distance="1000" swimtime="00:10:17.20" />
                    <SPLIT distance="1050" swimtime="00:10:48.08" />
                    <SPLIT distance="1100" swimtime="00:11:19.43" />
                    <SPLIT distance="1150" swimtime="00:11:50.87" />
                    <SPLIT distance="1200" swimtime="00:12:22.49" />
                    <SPLIT distance="1250" swimtime="00:12:53.77" />
                    <SPLIT distance="1300" swimtime="00:13:24.61" />
                    <SPLIT distance="1350" swimtime="00:13:56.05" />
                    <SPLIT distance="1400" swimtime="00:14:27.00" />
                    <SPLIT distance="1450" swimtime="00:14:57.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Hallage Papp" birthdate="2012-07-02" gender="M" nation="BRA" license="377042" swrid="5588736" athleteid="2312" externalid="377042">
              <RESULTS>
                <RESULT eventid="1077" points="121" swimtime="00:00:44.65" resultid="2313" heatid="3414" lane="8" entrytime="00:00:47.64" entrycourse="SCM" />
                <RESULT eventid="1065" points="120" swimtime="00:01:51.80" resultid="2314" heatid="3398" lane="1" entrytime="00:01:57.95" entrycourse="SCM" />
                <RESULT eventid="1105" points="119" swimtime="00:01:40.06" resultid="2315" heatid="3449" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="158" swimtime="00:00:37.26" resultid="2316" heatid="3485" lane="7" entrytime="00:00:38.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Fontoura" birthdate="2010-08-26" gender="M" nation="BRA" license="338922" swrid="5600167" athleteid="1940" externalid="338922">
              <RESULTS>
                <RESULT eventid="1184" points="256" swimtime="00:00:34.23" resultid="1941" heatid="3520" lane="8" />
                <RESULT eventid="1152" points="329" swimtime="00:05:07.25" resultid="1942" heatid="3498" lane="3" entrytime="00:05:39.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:12.09" />
                    <SPLIT distance="150" swimtime="00:01:51.24" />
                    <SPLIT distance="200" swimtime="00:02:31.00" />
                    <SPLIT distance="250" swimtime="00:03:09.94" />
                    <SPLIT distance="300" swimtime="00:03:49.85" />
                    <SPLIT distance="350" swimtime="00:04:29.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="277" swimtime="00:02:48.07" resultid="1943" heatid="3558" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="100" swimtime="00:01:22.45" />
                    <SPLIT distance="150" swimtime="00:02:10.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="238" swimtime="00:01:17.06" resultid="1944" heatid="3598" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="332" swimtime="00:01:04.71" resultid="1945" heatid="3576" lane="7" entrytime="00:01:13.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Poletto Abrahao" birthdate="2014-10-20" gender="M" nation="BRA" license="382128" swrid="5602571" athleteid="2388" externalid="382128">
              <RESULTS>
                <RESULT eventid="1095" points="150" swimtime="00:01:24.33" resultid="2389" heatid="3442" lane="6" entrytime="00:01:34.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="161" swimtime="00:00:45.79" resultid="2390" heatid="3404" lane="4" entrytime="00:00:46.30" entrycourse="SCM" />
                <RESULT eventid="1111" points="129" swimtime="00:00:42.97" resultid="2391" heatid="3459" lane="5" entrytime="00:00:44.53" entrycourse="SCM" />
                <RESULT eventid="1131" points="169" swimtime="00:00:36.40" resultid="2392" heatid="3474" lane="3" entrytime="00:00:39.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Estevao" lastname="Valduga Artigas" birthdate="2009-06-01" gender="M" nation="BRA" license="339556" swrid="5600267" athleteid="1832" externalid="339556" />
            <ATHLETE firstname="Gael" lastname="Gluck" birthdate="2011-01-28" gender="M" nation="BRA" license="366891" swrid="5588726" athleteid="1968" externalid="366891">
              <RESULTS>
                <RESULT eventid="1200" points="196" reactiontime="+76" swimtime="00:01:23.20" resultid="1969" heatid="3529" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="298" swimtime="00:01:22.74" resultid="1970" heatid="3511" lane="7" entrytime="00:01:25.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="297" swimtime="00:00:30.19" resultid="1971" heatid="3545" lane="4" entrytime="00:00:30.57" entrycourse="SCM" />
                <RESULT eventid="1264" points="339" swimtime="00:20:13.53" resultid="1972" heatid="3583" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.85" />
                    <SPLIT distance="100" swimtime="00:01:15.13" />
                    <SPLIT distance="150" swimtime="00:01:55.09" />
                    <SPLIT distance="200" swimtime="00:02:35.67" />
                    <SPLIT distance="250" swimtime="00:03:16.43" />
                    <SPLIT distance="300" swimtime="00:03:56.98" />
                    <SPLIT distance="350" swimtime="00:04:37.58" />
                    <SPLIT distance="400" swimtime="00:05:19.13" />
                    <SPLIT distance="450" swimtime="00:06:00.54" />
                    <SPLIT distance="500" swimtime="00:06:41.66" />
                    <SPLIT distance="550" swimtime="00:07:22.43" />
                    <SPLIT distance="600" swimtime="00:08:03.06" />
                    <SPLIT distance="650" swimtime="00:08:43.80" />
                    <SPLIT distance="700" swimtime="00:09:24.33" />
                    <SPLIT distance="750" swimtime="00:10:05.08" />
                    <SPLIT distance="800" swimtime="00:10:45.12" />
                    <SPLIT distance="850" swimtime="00:11:25.16" />
                    <SPLIT distance="900" swimtime="00:12:05.56" />
                    <SPLIT distance="950" swimtime="00:12:46.26" />
                    <SPLIT distance="1000" swimtime="00:13:26.80" />
                    <SPLIT distance="1050" swimtime="00:14:07.38" />
                    <SPLIT distance="1100" swimtime="00:14:48.49" />
                    <SPLIT distance="1150" swimtime="00:15:29.52" />
                    <SPLIT distance="1200" swimtime="00:16:09.98" />
                    <SPLIT distance="1250" swimtime="00:16:50.81" />
                    <SPLIT distance="1300" swimtime="00:17:31.77" />
                    <SPLIT distance="1350" swimtime="00:18:12.69" />
                    <SPLIT distance="1400" swimtime="00:18:54.09" />
                    <SPLIT distance="1450" swimtime="00:19:35.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="331" swimtime="00:01:04.76" resultid="1973" heatid="3577" lane="7" entrytime="00:01:08.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Schiavo Vianna" birthdate="2013-04-27" gender="F" nation="BRA" license="391005" swrid="5602582" athleteid="2419" externalid="391005">
              <RESULTS>
                <RESULT eventid="1062" status="DSQ" swimtime="00:03:33.49" resultid="2420" heatid="3392" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1086" points="137" swimtime="00:03:33.54" resultid="2421" heatid="3425" lane="3" entrytime="00:03:51.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.16" />
                    <SPLIT distance="100" swimtime="00:01:46.02" />
                    <SPLIT distance="150" swimtime="00:02:41.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="138" swimtime="00:01:49.19" resultid="2422" heatid="3446" lane="2" entrytime="00:02:12.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="170" swimtime="00:00:41.32" resultid="2423" heatid="3478" lane="7" entrytime="00:00:47.12" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Albuquerque" birthdate="2008-03-14" gender="F" nation="BRA" license="324787" swrid="5315259" athleteid="1725" externalid="324787">
              <RESULTS>
                <RESULT eventid="1160" points="561" swimtime="00:01:15.57" resultid="1726" heatid="3506" lane="3" entrytime="00:01:17.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="481" swimtime="00:02:35.52" resultid="1727" heatid="3552" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="100" swimtime="00:01:17.10" />
                    <SPLIT distance="150" swimtime="00:02:00.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="502" swimtime="00:00:35.68" resultid="1728" heatid="3604" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Massimo" lastname="Puppi Cardoso" birthdate="2015-03-30" gender="M" nation="BRA" license="406742" athleteid="2643" externalid="406742">
              <RESULTS>
                <RESULT eventid="1083" points="47" reactiontime="+67" swimtime="00:01:00.99" resultid="2644" heatid="3421" lane="3" />
                <RESULT eventid="1071" points="45" swimtime="00:01:09.85" resultid="2645" heatid="3402" lane="1" />
                <RESULT eventid="1111" points="25" swimtime="00:01:13.69" resultid="2646" heatid="3456" lane="5" />
                <RESULT eventid="1131" points="49" swimtime="00:00:55.00" resultid="2647" heatid="3472" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Xavier Jardim" birthdate="2012-01-23" gender="M" nation="BRA" license="369259" swrid="5641781" athleteid="2065" externalid="369259">
              <RESULTS>
                <RESULT eventid="1089" points="247" swimtime="00:02:38.17" resultid="2066" heatid="3434" lane="5" entrytime="00:02:39.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:16.28" />
                    <SPLIT distance="150" swimtime="00:01:58.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="186" reactiontime="+80" swimtime="00:00:38.73" resultid="2067" heatid="3415" lane="6" entrytime="00:00:39.21" entrycourse="SCM" />
                <RESULT eventid="1121" points="148" swimtime="00:01:30.22" resultid="2068" heatid="3464" lane="2" entrytime="00:01:37.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="241" swimtime="00:00:32.37" resultid="2069" heatid="3488" lane="7" entrytime="00:00:32.37" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariana" lastname="Stoberl" birthdate="2010-07-09" gender="F" nation="BRA" license="356250" swrid="5600265" athleteid="1886" externalid="356250">
              <RESULTS>
                <RESULT eventid="1144" points="444" swimtime="00:05:03.18" resultid="1887" heatid="3490" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.43" />
                    <SPLIT distance="100" swimtime="00:01:12.57" />
                    <SPLIT distance="150" swimtime="00:01:50.56" />
                    <SPLIT distance="200" swimtime="00:02:29.07" />
                    <SPLIT distance="250" swimtime="00:03:08.07" />
                    <SPLIT distance="300" swimtime="00:03:47.24" />
                    <SPLIT distance="350" swimtime="00:04:26.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="456" swimtime="00:00:29.79" resultid="1888" heatid="3539" lane="7" entrytime="00:00:30.16" entrycourse="SCM" />
                <RESULT eventid="1224" points="348" swimtime="00:02:53.17" resultid="1889" heatid="3551" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:01:21.96" />
                    <SPLIT distance="150" swimtime="00:02:15.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="261" swimtime="00:01:24.51" resultid="1890" heatid="3595" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="419" swimtime="00:01:07.10" resultid="1891" heatid="3570" lane="7" entrytime="00:01:04.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Rossi Mattioli" birthdate="2013-05-08" gender="F" nation="BRA" license="376988" swrid="5588892" athleteid="2332" externalid="376988">
              <RESULTS>
                <RESULT eventid="1062" points="225" swimtime="00:01:42.50" resultid="2333" heatid="3394" lane="1" />
                <RESULT eventid="1086" points="257" swimtime="00:02:53.28" resultid="2334" heatid="3427" lane="1" entrytime="00:02:59.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                    <SPLIT distance="100" swimtime="00:01:25.95" />
                    <SPLIT distance="150" swimtime="00:02:11.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="250" swimtime="00:01:29.64" resultid="2335" heatid="3447" lane="2" entrytime="00:01:39.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="297" swimtime="00:00:34.36" resultid="2336" heatid="3480" lane="2" entrytime="00:00:36.21" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rene" lastname="Osternack Erbe" birthdate="2011-04-03" gender="M" nation="BRA" license="366907" swrid="5588842" athleteid="2022" externalid="366907">
              <RESULTS>
                <RESULT eventid="1200" points="220" reactiontime="+78" swimtime="00:01:20.02" resultid="2023" heatid="3530" lane="6" entrytime="00:01:22.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="310" swimtime="00:05:13.55" resultid="2024" heatid="3499" lane="6" entrytime="00:05:27.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:14.73" />
                    <SPLIT distance="150" swimtime="00:01:55.02" />
                    <SPLIT distance="200" swimtime="00:02:36.23" />
                    <SPLIT distance="250" swimtime="00:03:15.55" />
                    <SPLIT distance="300" swimtime="00:03:56.79" />
                    <SPLIT distance="350" swimtime="00:04:35.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="271" swimtime="00:00:31.14" resultid="2025" heatid="3545" lane="2" entrytime="00:00:31.30" entrycourse="SCM" />
                <RESULT eventid="1232" points="224" swimtime="00:03:00.40" resultid="2026" heatid="3559" lane="7" entrytime="00:03:02.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                    <SPLIT distance="100" swimtime="00:01:25.21" />
                    <SPLIT distance="150" swimtime="00:02:22.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="153" swimtime="00:01:29.17" resultid="2027" heatid="3600" lane="7" entrytime="00:01:36.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Godino" birthdate="2010-04-27" gender="F" nation="BRA" license="356355" swrid="5600176" athleteid="1922" externalid="356355">
              <RESULTS>
                <RESULT eventid="1144" points="411" swimtime="00:05:11.09" resultid="1923" heatid="3493" lane="8" entrytime="00:05:32.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                    <SPLIT distance="100" swimtime="00:01:14.21" />
                    <SPLIT distance="150" swimtime="00:01:54.03" />
                    <SPLIT distance="200" swimtime="00:02:33.66" />
                    <SPLIT distance="250" swimtime="00:03:13.12" />
                    <SPLIT distance="300" swimtime="00:03:52.80" />
                    <SPLIT distance="350" swimtime="00:04:32.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="341" swimtime="00:00:32.81" resultid="1924" heatid="3537" lane="1" entrytime="00:00:32.81" entrycourse="SCM" />
                <RESULT eventid="1192" points="279" reactiontime="+87" swimtime="00:01:23.98" resultid="1925" heatid="3524" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="294" swimtime="00:03:03.15" resultid="1926" heatid="3551" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.33" />
                    <SPLIT distance="100" swimtime="00:01:29.20" />
                    <SPLIT distance="150" swimtime="00:02:25.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="360" swimtime="00:01:10.61" resultid="1927" heatid="3567" lane="2" entrytime="00:01:12.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Mayer Paludetto" birthdate="2012-10-30" gender="F" nation="BRA" license="369264" swrid="5588811" athleteid="2080" externalid="369264">
              <RESULTS>
                <RESULT eventid="1062" points="277" swimtime="00:01:35.63" resultid="2081" heatid="3394" lane="3" entrytime="00:01:36.95" entrycourse="SCM" />
                <RESULT eventid="1074" points="322" swimtime="00:00:36.82" resultid="2082" heatid="3410" lane="3" entrytime="00:00:38.11" entrycourse="SCM" />
                <RESULT eventid="1102" points="341" swimtime="00:01:20.88" resultid="2083" heatid="3445" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1118" points="219" swimtime="00:01:29.57" resultid="2084" heatid="3462" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Fortes Traub" birthdate="2012-04-26" gender="M" nation="BRA" license="369532" swrid="5588707" athleteid="2156" externalid="369532">
              <RESULTS>
                <RESULT eventid="1089" points="187" swimtime="00:02:53.50" resultid="2157" heatid="3432" lane="6" entrytime="00:03:01.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:01:25.13" />
                    <SPLIT distance="150" swimtime="00:02:10.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="132" reactiontime="+72" swimtime="00:00:43.32" resultid="2158" heatid="3412" lane="6" />
                <RESULT eventid="1105" status="DSQ" swimtime="00:01:37.19" resultid="2159" heatid="3450" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="164" swimtime="00:00:36.81" resultid="2160" heatid="3486" lane="8" entrytime="00:00:36.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Tallao Benke" birthdate="2012-01-02" gender="F" nation="BRA" license="376984" swrid="5588931" athleteid="2291" externalid="376984">
              <RESULTS>
                <RESULT eventid="1086" points="445" swimtime="00:02:24.44" resultid="2292" heatid="3427" lane="4" entrytime="00:02:48.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.36" />
                    <SPLIT distance="100" swimtime="00:01:09.74" />
                    <SPLIT distance="150" swimtime="00:01:47.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="401" swimtime="00:00:34.22" resultid="2293" heatid="3410" lane="4" entrytime="00:00:37.68" entrycourse="SCM" />
                <RESULT eventid="1118" points="408" swimtime="00:01:12.85" resultid="2294" heatid="3462" lane="4" entrytime="00:01:21.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="451" swimtime="00:00:29.88" resultid="2295" heatid="3481" lane="4" entrytime="00:00:32.23" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="De Czarnecki" birthdate="2008-06-24" gender="M" nation="BRA" license="329641" swrid="5600146" athleteid="1746" externalid="329641">
              <RESULTS>
                <RESULT eventid="1200" points="511" reactiontime="+67" swimtime="00:01:00.44" resultid="1747" heatid="3528" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="443" swimtime="00:01:02.67" resultid="1748" heatid="3599" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="506" swimtime="00:00:56.26" resultid="1749" heatid="3574" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Pellanda" birthdate="2010-11-12" gender="M" nation="BRA" license="356352" swrid="5600233" athleteid="1904" externalid="356352">
              <RESULTS>
                <RESULT eventid="1168" points="316" swimtime="00:01:21.12" resultid="1905" heatid="3510" lane="4" entrytime="00:01:26.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="535" swimtime="00:04:21.43" resultid="1906" heatid="3500" lane="8" entrytime="00:05:01.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.96" />
                    <SPLIT distance="100" swimtime="00:01:02.33" />
                    <SPLIT distance="150" swimtime="00:01:35.50" />
                    <SPLIT distance="200" swimtime="00:02:09.06" />
                    <SPLIT distance="250" swimtime="00:02:42.47" />
                    <SPLIT distance="300" swimtime="00:03:15.40" />
                    <SPLIT distance="350" swimtime="00:03:48.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="368" swimtime="00:00:28.13" resultid="1907" heatid="3546" lane="3" entrytime="00:00:29.02" entrycourse="SCM" />
                <RESULT eventid="1232" points="399" swimtime="00:02:28.86" resultid="1908" heatid="3560" lane="7" entrytime="00:02:42.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                    <SPLIT distance="100" swimtime="00:01:10.01" />
                    <SPLIT distance="150" swimtime="00:01:56.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="296" swimtime="00:01:11.62" resultid="1909" heatid="3599" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Pens Correa" birthdate="2015-11-27" gender="M" nation="BRA" license="393262" swrid="5616449" athleteid="2520" externalid="393262">
              <RESULTS>
                <RESULT eventid="1095" points="135" swimtime="00:01:27.24" resultid="2521" heatid="3439" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="138" swimtime="00:00:42.75" resultid="2522" heatid="3423" lane="2" entrytime="00:00:48.79" entrycourse="SCM" />
                <RESULT eventid="1111" points="144" swimtime="00:00:41.42" resultid="2523" heatid="3459" lane="8" entrytime="00:00:57.16" entrycourse="SCM" />
                <RESULT eventid="1131" points="153" swimtime="00:00:37.64" resultid="2524" heatid="3474" lane="1" entrytime="00:00:42.42" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Jardim" birthdate="2010-03-23" gender="F" nation="BRA" license="368006" swrid="5600192" athleteid="2043" externalid="368006">
              <RESULTS>
                <RESULT eventid="1144" points="342" swimtime="00:05:30.74" resultid="2044" heatid="3489" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                    <SPLIT distance="100" swimtime="00:01:16.51" />
                    <SPLIT distance="150" swimtime="00:01:58.84" />
                    <SPLIT distance="200" swimtime="00:02:41.50" />
                    <SPLIT distance="250" swimtime="00:03:24.84" />
                    <SPLIT distance="300" swimtime="00:04:08.45" />
                    <SPLIT distance="350" swimtime="00:04:51.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="367" swimtime="00:00:32.00" resultid="2045" heatid="3537" lane="7" entrytime="00:00:32.30" entrycourse="SCM" />
                <RESULT eventid="1224" points="302" swimtime="00:03:01.49" resultid="2046" heatid="3552" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.34" />
                    <SPLIT distance="100" swimtime="00:01:25.95" />
                    <SPLIT distance="150" swimtime="00:02:22.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="260" swimtime="00:01:24.61" resultid="2047" heatid="3595" lane="3" entrytime="00:01:25.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="355" swimtime="00:01:10.92" resultid="2048" heatid="3568" lane="8" entrytime="00:01:10.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucca" lastname="Cruz Tonin" birthdate="2004-03-19" gender="M" nation="BRA" license="270821" swrid="5622272" athleteid="2040" externalid="270821" level="FUNDESPORT">
              <RESULTS>
                <RESULT eventid="1280" points="631" reactiontime="+46" swimtime="00:00:25.77" resultid="2041" heatid="3593" lane="4" entrytime="00:00:25.71" entrycourse="SCM" />
                <RESULT eventid="1248" points="612" swimtime="00:00:52.79" resultid="2042" heatid="3573" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Ramos Marcon" birthdate="2008-01-12" gender="M" nation="BRA" license="372281" swrid="5600240" athleteid="2393" externalid="372281">
              <RESULTS>
                <RESULT eventid="1216" points="492" swimtime="00:00:25.52" resultid="2394" heatid="3549" lane="6" entrytime="00:00:26.11" entrycourse="SCM" />
                <RESULT eventid="1248" points="519" swimtime="00:00:55.78" resultid="2395" heatid="3580" lane="2" entrytime="00:00:56.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Severo" lastname="Berger Leal" birthdate="2008-08-05" gender="M" nation="BRA" license="330073" swrid="5449277" athleteid="1823" externalid="330073">
              <RESULTS>
                <RESULT eventid="1184" points="350" swimtime="00:00:30.86" resultid="1824" heatid="3518" lane="6" />
                <RESULT eventid="1168" points="407" swimtime="00:01:14.57" resultid="1825" heatid="3512" lane="3" entrytime="00:01:14.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="375" swimtime="00:00:34.57" resultid="1826" heatid="3608" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Estevao" lastname="Sarmento Ribas" birthdate="2012-11-19" gender="M" nation="BRA" license="369273" swrid="5588898" athleteid="2110" externalid="369273">
              <RESULTS>
                <RESULT eventid="1089" points="301" swimtime="00:02:28.13" resultid="2111" heatid="3434" lane="4" entrytime="00:02:34.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:11.76" />
                    <SPLIT distance="150" swimtime="00:01:50.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="185" reactiontime="+83" swimtime="00:00:38.76" resultid="2112" heatid="3412" lane="5" />
                <RESULT eventid="1121" points="176" swimtime="00:01:25.25" resultid="2113" heatid="3464" lane="6" entrytime="00:01:32.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="265" swimtime="00:00:31.37" resultid="2114" heatid="3488" lane="5" entrytime="00:00:31.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marco" lastname="Antonio Barichello" birthdate="2013-01-14" gender="M" nation="BRA" license="376969" swrid="5588526" athleteid="2235" externalid="376969">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="2236" heatid="3431" lane="1" entrytime="00:03:39.13" entrycourse="SCM" />
                <RESULT eventid="1065" status="DNS" swimtime="00:00:00.00" resultid="2237" heatid="3397" lane="8" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="2238" heatid="3449" lane="4" />
                <RESULT eventid="1141" status="DNS" swimtime="00:00:00.00" resultid="2239" heatid="3483" lane="4" entrytime="00:00:45.42" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Vitoria Kuzmann Cercal" birthdate="2009-04-10" gender="F" nation="BRA" license="339082" swrid="5600274" athleteid="1850" externalid="339082">
              <RESULTS>
                <RESULT eventid="1144" points="489" swimtime="00:04:53.44" resultid="1851" heatid="3490" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                    <SPLIT distance="100" swimtime="00:01:08.74" />
                    <SPLIT distance="150" swimtime="00:01:45.53" />
                    <SPLIT distance="200" swimtime="00:02:22.92" />
                    <SPLIT distance="250" swimtime="00:03:00.49" />
                    <SPLIT distance="300" swimtime="00:03:38.62" />
                    <SPLIT distance="350" swimtime="00:04:17.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="392" reactiontime="+84" swimtime="00:01:14.98" resultid="1852" heatid="3524" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="431" swimtime="00:02:41.27" resultid="1853" heatid="3555" lane="5" entrytime="00:02:49.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                    <SPLIT distance="100" swimtime="00:01:14.79" />
                    <SPLIT distance="150" swimtime="00:02:04.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="475" swimtime="00:01:04.40" resultid="1854" heatid="3569" lane="5" entrytime="00:01:06.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelo" lastname="Vanhazebrouck" birthdate="2010-01-09" gender="M" nation="BRA" license="339043" swrid="5600269" athleteid="1869" externalid="339043">
              <RESULTS>
                <RESULT eventid="1168" points="330" swimtime="00:01:19.92" resultid="1870" heatid="3508" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="436" swimtime="00:04:39.79" resultid="1871" heatid="3500" lane="4" entrytime="00:04:46.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                    <SPLIT distance="100" swimtime="00:01:04.30" />
                    <SPLIT distance="150" swimtime="00:01:38.91" />
                    <SPLIT distance="200" swimtime="00:02:14.25" />
                    <SPLIT distance="250" swimtime="00:02:50.14" />
                    <SPLIT distance="300" swimtime="00:03:26.31" />
                    <SPLIT distance="350" swimtime="00:04:03.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="404" swimtime="00:00:27.26" resultid="1872" heatid="3547" lane="2" entrytime="00:00:28.65" entrycourse="SCM" />
                <RESULT eventid="1312" points="358" swimtime="00:00:35.11" resultid="1873" heatid="3611" lane="2" entrytime="00:00:37.67" entrycourse="SCM" />
                <RESULT eventid="1248" points="429" swimtime="00:00:59.45" resultid="1874" heatid="3578" lane="3" entrytime="00:01:01.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Vieira Motta" birthdate="2009-09-19" gender="M" nation="BRA" license="339064" swrid="5600271" athleteid="1858" externalid="339064">
              <RESULTS>
                <RESULT eventid="1200" points="364" swimtime="00:01:07.64" resultid="1859" heatid="3531" lane="8" entrytime="00:01:16.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="461" swimtime="00:18:15.80" resultid="1860" heatid="3584" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:10.27" />
                    <SPLIT distance="150" swimtime="00:01:46.65" />
                    <SPLIT distance="200" swimtime="00:02:23.15" />
                    <SPLIT distance="250" swimtime="00:02:59.77" />
                    <SPLIT distance="300" swimtime="00:03:36.20" />
                    <SPLIT distance="350" swimtime="00:04:12.89" />
                    <SPLIT distance="400" swimtime="00:04:50.14" />
                    <SPLIT distance="450" swimtime="00:05:27.52" />
                    <SPLIT distance="500" swimtime="00:06:04.23" />
                    <SPLIT distance="550" swimtime="00:06:41.92" />
                    <SPLIT distance="600" swimtime="00:07:19.09" />
                    <SPLIT distance="650" swimtime="00:07:56.07" />
                    <SPLIT distance="700" swimtime="00:08:33.07" />
                    <SPLIT distance="750" swimtime="00:09:09.66" />
                    <SPLIT distance="800" swimtime="00:09:46.16" />
                    <SPLIT distance="850" swimtime="00:10:23.15" />
                    <SPLIT distance="900" swimtime="00:11:00.15" />
                    <SPLIT distance="950" swimtime="00:11:37.04" />
                    <SPLIT distance="1000" swimtime="00:12:13.40" />
                    <SPLIT distance="1050" swimtime="00:12:50.23" />
                    <SPLIT distance="1100" swimtime="00:13:27.31" />
                    <SPLIT distance="1150" swimtime="00:14:04.36" />
                    <SPLIT distance="1200" swimtime="00:14:41.23" />
                    <SPLIT distance="1250" swimtime="00:15:18.04" />
                    <SPLIT distance="1300" swimtime="00:15:54.23" />
                    <SPLIT distance="1350" swimtime="00:16:30.00" />
                    <SPLIT distance="1400" swimtime="00:17:06.29" />
                    <SPLIT distance="1450" swimtime="00:17:41.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Steven" lastname="Matheussi Viana E Silva" birthdate="2012-05-03" gender="M" nation="BRA" license="376986" swrid="5588810" athleteid="2337" externalid="376986">
              <RESULTS>
                <RESULT eventid="1089" points="210" swimtime="00:02:47.12" resultid="2338" heatid="3433" lane="8" entrytime="00:02:56.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="100" swimtime="00:01:20.45" />
                    <SPLIT distance="150" swimtime="00:02:03.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="181" swimtime="00:01:37.58" resultid="2339" heatid="3398" lane="7" entrytime="00:01:45.26" entrycourse="SCM" />
                <RESULT eventid="1121" points="160" swimtime="00:01:28.01" resultid="2340" heatid="3464" lane="7" entrytime="00:01:38.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="193" swimtime="00:00:34.84" resultid="2341" heatid="3485" lane="1" entrytime="00:00:38.17" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Vian" birthdate="2014-03-25" gender="F" nation="BRA" license="393919" swrid="5641779" athleteid="2540" externalid="393919">
              <RESULTS>
                <RESULT eventid="1092" points="119" swimtime="00:01:42.04" resultid="2541" heatid="3437" lane="4" entrytime="00:01:55.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="125" swimtime="00:00:50.47" resultid="2542" heatid="3419" lane="6" entrytime="00:00:51.10" entrycourse="SCM" />
                <RESULT eventid="1108" points="83" swimtime="00:00:55.88" resultid="2543" heatid="3454" lane="4" entrytime="00:01:03.01" entrycourse="SCM" />
                <RESULT eventid="1128" points="154" swimtime="00:00:42.69" resultid="2544" heatid="3468" lane="4" entrytime="00:00:45.31" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia" lastname="Salesi Chicon" birthdate="2002-04-16" gender="F" nation="BRA" license="250865" swrid="5600255" athleteid="2413" externalid="250865">
              <RESULTS>
                <RESULT eventid="1144" points="757" swimtime="00:04:13.76" resultid="2414" heatid="3494" lane="4" entrytime="00:04:14.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.07" />
                    <SPLIT distance="100" swimtime="00:01:00.24" />
                    <SPLIT distance="150" swimtime="00:01:32.07" />
                    <SPLIT distance="200" swimtime="00:02:04.43" />
                    <SPLIT distance="250" swimtime="00:02:36.78" />
                    <SPLIT distance="300" swimtime="00:03:09.17" />
                    <SPLIT distance="350" swimtime="00:03:41.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="717" swimtime="00:16:54.63" resultid="2415" heatid="3582" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="100" swimtime="00:01:04.43" />
                    <SPLIT distance="150" swimtime="00:01:37.87" />
                    <SPLIT distance="200" swimtime="00:02:11.65" />
                    <SPLIT distance="250" swimtime="00:02:45.50" />
                    <SPLIT distance="300" swimtime="00:03:19.33" />
                    <SPLIT distance="350" swimtime="00:03:53.06" />
                    <SPLIT distance="400" swimtime="00:04:26.81" />
                    <SPLIT distance="450" swimtime="00:05:00.55" />
                    <SPLIT distance="500" swimtime="00:05:34.28" />
                    <SPLIT distance="550" swimtime="00:06:07.96" />
                    <SPLIT distance="600" swimtime="00:06:41.65" />
                    <SPLIT distance="650" swimtime="00:07:15.03" />
                    <SPLIT distance="700" swimtime="00:07:48.57" />
                    <SPLIT distance="750" swimtime="00:08:22.64" />
                    <SPLIT distance="800" swimtime="00:08:56.25" />
                    <SPLIT distance="850" swimtime="00:09:30.46" />
                    <SPLIT distance="900" swimtime="00:10:04.89" />
                    <SPLIT distance="950" swimtime="00:10:38.74" />
                    <SPLIT distance="1000" swimtime="00:11:12.94" />
                    <SPLIT distance="1050" swimtime="00:11:46.69" />
                    <SPLIT distance="1100" swimtime="00:12:20.66" />
                    <SPLIT distance="1150" swimtime="00:12:54.36" />
                    <SPLIT distance="1200" swimtime="00:13:28.62" />
                    <SPLIT distance="1250" swimtime="00:14:03.10" />
                    <SPLIT distance="1300" swimtime="00:14:37.58" />
                    <SPLIT distance="1350" swimtime="00:15:11.85" />
                    <SPLIT distance="1400" swimtime="00:15:46.48" />
                    <SPLIT distance="1450" swimtime="00:16:20.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luigi" lastname="Antoniuk Paganini" birthdate="2014-11-13" gender="M" nation="BRA" license="382127" swrid="5602509" athleteid="2383" externalid="382127">
              <RESULTS>
                <RESULT eventid="1083" points="100" swimtime="00:00:47.63" resultid="2384" heatid="3423" lane="7" entrytime="00:00:50.50" entrycourse="SCM" />
                <RESULT eventid="1071" points="72" swimtime="00:00:59.72" resultid="2385" heatid="3404" lane="1" entrytime="00:01:01.72" entrycourse="SCM" />
                <RESULT eventid="1111" points="81" swimtime="00:00:50.20" resultid="2386" heatid="3459" lane="2" entrytime="00:00:49.47" entrycourse="SCM" />
                <RESULT eventid="1131" points="104" swimtime="00:00:42.84" resultid="2387" heatid="3474" lane="8" entrytime="00:00:42.83" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Emili Da Silva Gomes Xavier" birthdate="2010-09-08" gender="F" nation="BRA" license="372519" athleteid="2708" externalid="372519">
              <RESULTS>
                <RESULT eventid="1144" points="339" swimtime="00:05:31.60" resultid="2709" heatid="3489" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.64" />
                    <SPLIT distance="100" swimtime="00:01:18.53" />
                    <SPLIT distance="150" swimtime="00:02:00.78" />
                    <SPLIT distance="200" swimtime="00:02:43.22" />
                    <SPLIT distance="250" swimtime="00:03:26.26" />
                    <SPLIT distance="300" swimtime="00:04:09.56" />
                    <SPLIT distance="350" swimtime="00:04:52.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="287" reactiontime="+73" swimtime="00:01:23.16" resultid="2710" heatid="3524" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="334" swimtime="00:01:29.87" resultid="2711" heatid="3503" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="302" swimtime="00:03:01.49" resultid="2712" heatid="3553" lane="4" entrytime="00:03:08.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                    <SPLIT distance="100" swimtime="00:01:26.49" />
                    <SPLIT distance="150" swimtime="00:02:19.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="348" swimtime="00:01:11.40" resultid="2713" heatid="3567" lane="3" entrytime="00:01:11.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Zaroni" birthdate="2010-03-03" gender="F" nation="BRA" license="356345" swrid="5600282" athleteid="1779" externalid="356345">
              <RESULTS>
                <RESULT eventid="1144" points="399" swimtime="00:05:14.18" resultid="1780" heatid="3490" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                    <SPLIT distance="100" swimtime="00:01:14.69" />
                    <SPLIT distance="150" swimtime="00:01:55.06" />
                    <SPLIT distance="200" swimtime="00:02:35.62" />
                    <SPLIT distance="250" swimtime="00:03:15.92" />
                    <SPLIT distance="300" swimtime="00:03:56.44" />
                    <SPLIT distance="350" swimtime="00:04:37.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="409" swimtime="00:00:30.88" resultid="1781" heatid="3537" lane="2" entrytime="00:00:32.29" entrycourse="SCM" />
                <RESULT eventid="1160" points="424" swimtime="00:01:22.95" resultid="1782" heatid="3506" lane="1" entrytime="00:01:21.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="383" swimtime="00:02:47.69" resultid="1783" heatid="3556" lane="1" entrytime="00:02:46.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                    <SPLIT distance="100" swimtime="00:01:22.71" />
                    <SPLIT distance="150" swimtime="00:02:09.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="432" swimtime="00:01:06.44" resultid="1784" heatid="3568" lane="7" entrytime="00:01:09.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maya" lastname="Assahida Moreria" birthdate="2014-02-24" gender="F" nation="BRA" license="391020" swrid="5602512" athleteid="2456" externalid="391020">
              <RESULTS>
                <RESULT eventid="1092" points="142" swimtime="00:01:36.19" resultid="2457" heatid="3438" lane="3" entrytime="00:01:33.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="98" swimtime="00:00:54.61" resultid="2458" heatid="3419" lane="8" entrytime="00:00:56.82" entrycourse="SCM" />
                <RESULT eventid="1108" points="99" swimtime="00:00:52.65" resultid="2459" heatid="3455" lane="3" entrytime="00:00:51.30" entrycourse="SCM" />
                <RESULT eventid="1128" points="154" swimtime="00:00:42.75" resultid="2460" heatid="3469" lane="6" entrytime="00:00:42.49" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Toscani Kim" birthdate="2013-02-15" gender="F" nation="BRA" license="372683" swrid="5588939" athleteid="2171" externalid="372683">
              <RESULTS>
                <RESULT eventid="1062" points="299" swimtime="00:01:33.19" resultid="2172" heatid="3393" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1086" points="286" swimtime="00:02:47.30" resultid="2173" heatid="3427" lane="3" entrytime="00:02:51.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                    <SPLIT distance="100" swimtime="00:01:21.83" />
                    <SPLIT distance="150" swimtime="00:02:05.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="282" swimtime="00:01:26.13" resultid="2174" heatid="3447" lane="6" entrytime="00:01:35.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1118" points="184" swimtime="00:01:34.90" resultid="2175" heatid="3461" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Galvao" birthdate="2011-03-11" gender="M" nation="BRA" license="381989" swrid="5602541" athleteid="2362" externalid="381989">
              <RESULTS>
                <RESULT eventid="1200" points="157" reactiontime="+73" swimtime="00:01:29.49" resultid="2363" heatid="3530" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="276" swimtime="00:05:25.67" resultid="2364" heatid="3498" lane="5" entrytime="00:05:34.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                    <SPLIT distance="100" swimtime="00:01:17.45" />
                    <SPLIT distance="150" swimtime="00:01:59.50" />
                    <SPLIT distance="200" swimtime="00:02:41.26" />
                    <SPLIT distance="250" swimtime="00:03:23.58" />
                    <SPLIT distance="300" swimtime="00:04:05.62" />
                    <SPLIT distance="350" swimtime="00:04:46.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="270" swimtime="00:00:31.17" resultid="2365" heatid="3545" lane="3" entrytime="00:00:31.14" entrycourse="SCM" />
                <RESULT eventid="1264" points="247" swimtime="00:22:28.55" resultid="2366" heatid="3583" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.08" />
                    <SPLIT distance="100" swimtime="00:01:25.99" />
                    <SPLIT distance="150" swimtime="00:02:11.61" />
                    <SPLIT distance="200" swimtime="00:02:57.81" />
                    <SPLIT distance="250" swimtime="00:03:42.81" />
                    <SPLIT distance="300" swimtime="00:04:28.32" />
                    <SPLIT distance="350" swimtime="00:05:13.99" />
                    <SPLIT distance="400" swimtime="00:05:59.59" />
                    <SPLIT distance="450" swimtime="00:06:45.24" />
                    <SPLIT distance="500" swimtime="00:07:31.58" />
                    <SPLIT distance="550" swimtime="00:08:17.49" />
                    <SPLIT distance="600" swimtime="00:09:02.25" />
                    <SPLIT distance="650" swimtime="00:09:47.84" />
                    <SPLIT distance="700" swimtime="00:10:33.04" />
                    <SPLIT distance="750" swimtime="00:11:18.14" />
                    <SPLIT distance="800" swimtime="00:12:03.88" />
                    <SPLIT distance="850" swimtime="00:12:49.29" />
                    <SPLIT distance="900" swimtime="00:13:34.18" />
                    <SPLIT distance="950" swimtime="00:14:19.59" />
                    <SPLIT distance="1000" swimtime="00:15:05.15" />
                    <SPLIT distance="1050" swimtime="00:15:51.62" />
                    <SPLIT distance="1100" swimtime="00:16:35.23" />
                    <SPLIT distance="1150" swimtime="00:17:19.97" />
                    <SPLIT distance="1200" swimtime="00:18:04.53" />
                    <SPLIT distance="1250" swimtime="00:18:49.62" />
                    <SPLIT distance="1300" swimtime="00:19:34.85" />
                    <SPLIT distance="1350" swimtime="00:20:19.87" />
                    <SPLIT distance="1400" swimtime="00:21:03.61" />
                    <SPLIT distance="1450" swimtime="00:21:47.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="269" swimtime="00:01:09.39" resultid="2367" heatid="3576" lane="5" entrytime="00:01:10.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Braga Amatuzzi" birthdate="2006-01-18" gender="M" nation="BRA" license="296650" swrid="5465902" athleteid="1769" externalid="296650">
              <RESULTS>
                <RESULT eventid="1168" points="686" swimtime="00:01:02.66" resultid="1770" heatid="3513" lane="4" entrytime="00:01:02.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="607" swimtime="00:00:23.80" resultid="1771" heatid="3542" lane="7" />
                <RESULT eventid="1232" points="634" swimtime="00:02:07.60" resultid="1772" heatid="3561" lane="5" entrytime="00:02:07.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.96" />
                    <SPLIT distance="100" swimtime="00:01:01.81" />
                    <SPLIT distance="150" swimtime="00:01:37.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" status="DNS" swimtime="00:00:00.00" resultid="1773" heatid="3612" lane="2" entrytime="00:00:31.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Lazzarotti Matias" birthdate="2012-03-19" gender="F" nation="BRA" license="391026" swrid="5602552" athleteid="2476" externalid="391026">
              <RESULTS>
                <RESULT eventid="1062" points="275" swimtime="00:01:35.88" resultid="2477" heatid="3393" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="340" swimtime="00:00:36.15" resultid="2478" heatid="3410" lane="2" entrytime="00:00:38.13" entrycourse="SCM" />
                <RESULT eventid="1102" points="305" swimtime="00:01:23.95" resultid="2479" heatid="3445" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="347" swimtime="00:00:32.63" resultid="2480" heatid="3481" lane="2" entrytime="00:00:33.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elisa" lastname="Osternack Almeida" birthdate="2015-04-14" gender="F" nation="BRA" license="406747" athleteid="2665" externalid="406747">
              <RESULTS>
                <RESULT eventid="1092" points="60" swimtime="00:02:07.84" resultid="2666" heatid="3435" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="80" reactiontime="+70" swimtime="00:00:58.37" resultid="2667" heatid="3417" lane="4" />
                <RESULT eventid="1108" points="48" swimtime="00:01:07.04" resultid="2668" heatid="3454" lane="2" />
                <RESULT eventid="1128" points="69" swimtime="00:00:55.82" resultid="2669" heatid="3466" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Correa Nascimento" birthdate="2009-01-19" gender="M" nation="BRA" license="342235" swrid="5600140" athleteid="1833" externalid="342235">
              <RESULTS>
                <RESULT eventid="1168" points="418" swimtime="00:01:13.90" resultid="1834" heatid="3511" lane="4" entrytime="00:01:21.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="446" swimtime="00:00:26.37" resultid="1835" heatid="3547" lane="5" entrytime="00:00:27.98" entrycourse="SCM" />
                <RESULT eventid="1232" points="387" swimtime="00:02:30.41" resultid="1836" heatid="3558" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                    <SPLIT distance="100" swimtime="00:01:10.62" />
                    <SPLIT distance="150" swimtime="00:01:56.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="492" swimtime="00:00:56.77" resultid="1837" heatid="3578" lane="5" entrytime="00:01:01.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enrico" lastname="Hallage Bianchini" birthdate="2014-02-27" gender="M" nation="BRA" license="397164" swrid="5661348" athleteid="2545" externalid="397164">
              <RESULTS>
                <RESULT eventid="1095" points="113" swimtime="00:01:32.72" resultid="2546" heatid="3439" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="93" reactiontime="+66" swimtime="00:00:48.67" resultid="2547" heatid="3422" lane="2" />
                <RESULT eventid="1111" points="89" swimtime="00:00:48.69" resultid="2548" heatid="3458" lane="7" />
                <RESULT eventid="1131" points="131" swimtime="00:00:39.66" resultid="2549" heatid="3470" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Karam Barbosa Lima" birthdate="2012-12-11" gender="F" nation="BRA" license="376956" swrid="5588758" athleteid="2201" externalid="376956">
              <RESULTS>
                <RESULT eventid="1086" points="332" swimtime="00:02:39.17" resultid="2202" heatid="3428" lane="2" entrytime="00:02:40.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                    <SPLIT distance="100" swimtime="00:01:16.66" />
                    <SPLIT distance="150" swimtime="00:01:58.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="299" swimtime="00:00:37.76" resultid="2203" heatid="3410" lane="6" entrytime="00:00:38.12" entrycourse="SCM" />
                <RESULT eventid="1102" points="277" swimtime="00:01:26.65" resultid="2204" heatid="3446" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="355" swimtime="00:00:32.38" resultid="2205" heatid="3481" lane="3" entrytime="00:00:32.75" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Spadari Soso" birthdate="2012-12-28" gender="F" nation="BRA" license="377313" swrid="5588921" athleteid="2685" externalid="377313">
              <RESULTS>
                <RESULT eventid="1062" status="DSQ" swimtime="00:01:41.43" resultid="2686" heatid="3393" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1086" points="260" swimtime="00:02:52.81" resultid="2687" heatid="3425" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.14" />
                    <SPLIT distance="100" swimtime="00:01:26.91" />
                    <SPLIT distance="150" swimtime="00:02:11.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="202" swimtime="00:01:36.18" resultid="2688" heatid="3445" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="306" swimtime="00:00:34.02" resultid="2689" heatid="3476" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joshua" lastname="Gomide Capraro" birthdate="2009-01-18" gender="M" nation="BRA" license="339030" swrid="5600177" athleteid="1754" externalid="339030">
              <RESULTS>
                <RESULT eventid="1152" points="509" swimtime="00:04:25.79" resultid="1755" heatid="3501" lane="6" entrytime="00:04:32.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                    <SPLIT distance="100" swimtime="00:01:02.54" />
                    <SPLIT distance="150" swimtime="00:01:35.97" />
                    <SPLIT distance="200" swimtime="00:02:09.99" />
                    <SPLIT distance="250" swimtime="00:02:44.24" />
                    <SPLIT distance="300" swimtime="00:03:18.57" />
                    <SPLIT distance="350" swimtime="00:03:52.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="527" swimtime="00:00:24.95" resultid="1756" heatid="3550" lane="1" entrytime="00:00:25.39" entrycourse="SCM" />
                <RESULT eventid="1248" points="539" swimtime="00:00:55.07" resultid="1757" heatid="3580" lane="5" entrytime="00:00:55.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Petraglia" birthdate="2012-03-28" gender="M" nation="BRA" license="369282" swrid="5602569" athleteid="2145" externalid="369282">
              <RESULTS>
                <RESULT eventid="1089" points="241" swimtime="00:02:39.55" resultid="2146" heatid="3434" lane="6" entrytime="00:02:42.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                    <SPLIT distance="100" swimtime="00:01:17.61" />
                    <SPLIT distance="150" swimtime="00:01:59.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="188" swimtime="00:01:36.36" resultid="2147" heatid="3398" lane="6" entrytime="00:01:39.29" entrycourse="SCM" />
                <RESULT eventid="1105" points="177" swimtime="00:01:27.67" resultid="2148" heatid="3451" lane="5" entrytime="00:01:29.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="221" swimtime="00:00:33.30" resultid="2149" heatid="3487" lane="1" entrytime="00:00:34.48" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Schmidt Wozniaki" birthdate="2012-07-07" gender="M" nation="BRA" license="376963" swrid="5588905" athleteid="2221" externalid="376963">
              <RESULTS>
                <RESULT eventid="1077" points="80" reactiontime="+69" swimtime="00:00:51.15" resultid="2222" heatid="3413" lane="4" entrytime="00:00:50.63" entrycourse="SCM" />
                <RESULT eventid="1065" points="124" swimtime="00:01:50.66" resultid="2223" heatid="3397" lane="4" entrytime="00:02:07.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" status="DSQ" swimtime="00:00:37.61" resultid="2224" heatid="3485" lane="6" entrytime="00:00:37.84" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Carcereri Navarro" birthdate="2013-12-19" gender="M" nation="BRA" license="376962" swrid="5588576" athleteid="2216" externalid="376962">
              <RESULTS>
                <RESULT eventid="1089" points="130" swimtime="00:03:16.08" resultid="2217" heatid="3432" lane="7" entrytime="00:03:07.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.20" />
                    <SPLIT distance="100" swimtime="00:01:34.16" />
                    <SPLIT distance="150" swimtime="00:02:27.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="146" swimtime="00:01:44.76" resultid="2218" heatid="3397" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="100" swimtime="00:01:42.72" resultid="2219" heatid="3464" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="166" swimtime="00:00:36.63" resultid="2220" heatid="3485" lane="3" entrytime="00:00:37.38" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia" lastname="Ziliotto Mehl" birthdate="2015-10-09" gender="F" nation="BRA" license="400122" swrid="5652905" athleteid="2580" externalid="400122">
              <RESULTS>
                <RESULT eventid="1092" points="82" swimtime="00:01:55.26" resultid="2581" heatid="3436" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="90" swimtime="00:01:03.12" resultid="2582" heatid="3399" lane="7" />
                <RESULT eventid="1108" points="49" swimtime="00:01:06.37" resultid="2583" heatid="3452" lane="7" />
                <RESULT eventid="1128" points="88" swimtime="00:00:51.36" resultid="2584" heatid="3465" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Guimaraes Mesquita" birthdate="2013-12-30" gender="F" nation="BRA" license="391027" swrid="5602544" athleteid="2481" externalid="391027">
              <RESULTS>
                <RESULT eventid="1062" points="134" swimtime="00:02:01.69" resultid="2482" heatid="3392" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1086" points="144" swimtime="00:03:30.16" resultid="2483" heatid="3426" lane="8" entrytime="00:03:31.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.59" />
                    <SPLIT distance="100" swimtime="00:01:43.54" />
                    <SPLIT distance="150" swimtime="00:02:37.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="141" swimtime="00:01:48.33" resultid="2484" heatid="3446" lane="3" entrytime="00:01:56.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="141" swimtime="00:00:43.97" resultid="2485" heatid="3478" lane="5" entrytime="00:00:43.95" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Salomao" birthdate="2012-05-07" gender="M" nation="BRA" license="369261" swrid="5602581" athleteid="2070" externalid="369261">
              <RESULTS>
                <RESULT eventid="1089" points="244" swimtime="00:02:38.99" resultid="2071" heatid="3434" lane="2" entrytime="00:02:42.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:01:16.82" />
                    <SPLIT distance="150" swimtime="00:01:58.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="171" reactiontime="+69" swimtime="00:00:39.80" resultid="2072" heatid="3414" lane="4" entrytime="00:00:41.14" entrycourse="SCM" />
                <RESULT eventid="1121" points="148" swimtime="00:01:30.26" resultid="2073" heatid="3464" lane="3" entrytime="00:01:28.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="223" swimtime="00:00:33.24" resultid="2074" heatid="3488" lane="8" entrytime="00:00:32.98" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Leao" birthdate="2011-09-18" gender="M" nation="BRA" license="366880" swrid="5602553" athleteid="1956" externalid="366880">
              <RESULTS>
                <RESULT eventid="1200" points="198" reactiontime="+76" swimtime="00:01:22.79" resultid="1957" heatid="3529" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="346" swimtime="00:05:02.33" resultid="1958" heatid="3499" lane="3" entrytime="00:05:16.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.90" />
                    <SPLIT distance="100" swimtime="00:01:11.69" />
                    <SPLIT distance="150" swimtime="00:01:50.36" />
                    <SPLIT distance="200" swimtime="00:02:29.44" />
                    <SPLIT distance="250" swimtime="00:03:08.78" />
                    <SPLIT distance="300" swimtime="00:03:47.79" />
                    <SPLIT distance="350" swimtime="00:04:26.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="248" swimtime="00:02:54.42" resultid="1959" heatid="3559" lane="2" entrytime="00:03:01.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                    <SPLIT distance="100" swimtime="00:01:22.50" />
                    <SPLIT distance="150" swimtime="00:02:16.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="192" swimtime="00:01:22.73" resultid="1960" heatid="3600" lane="2" entrytime="00:01:24.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="353" swimtime="00:19:57.66" resultid="1961" heatid="3584" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                    <SPLIT distance="100" swimtime="00:01:15.03" />
                    <SPLIT distance="150" swimtime="00:01:54.84" />
                    <SPLIT distance="200" swimtime="00:02:34.41" />
                    <SPLIT distance="250" swimtime="00:03:13.72" />
                    <SPLIT distance="300" swimtime="00:03:53.52" />
                    <SPLIT distance="350" swimtime="00:04:32.57" />
                    <SPLIT distance="400" swimtime="00:05:12.17" />
                    <SPLIT distance="450" swimtime="00:05:52.23" />
                    <SPLIT distance="500" swimtime="00:06:32.03" />
                    <SPLIT distance="550" swimtime="00:07:11.81" />
                    <SPLIT distance="600" swimtime="00:07:51.95" />
                    <SPLIT distance="650" swimtime="00:08:31.84" />
                    <SPLIT distance="700" swimtime="00:09:12.15" />
                    <SPLIT distance="750" swimtime="00:09:52.14" />
                    <SPLIT distance="800" swimtime="00:10:32.49" />
                    <SPLIT distance="850" swimtime="00:11:12.99" />
                    <SPLIT distance="900" swimtime="00:11:52.47" />
                    <SPLIT distance="950" swimtime="00:12:33.70" />
                    <SPLIT distance="1000" swimtime="00:13:15.01" />
                    <SPLIT distance="1050" swimtime="00:13:54.37" />
                    <SPLIT distance="1100" swimtime="00:14:35.20" />
                    <SPLIT distance="1150" swimtime="00:15:15.52" />
                    <SPLIT distance="1200" swimtime="00:15:56.29" />
                    <SPLIT distance="1250" swimtime="00:16:37.31" />
                    <SPLIT distance="1300" swimtime="00:17:18.09" />
                    <SPLIT distance="1350" swimtime="00:17:58.84" />
                    <SPLIT distance="1400" swimtime="00:18:39.42" />
                    <SPLIT distance="1450" swimtime="00:19:20.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Livia Bittencourt" birthdate="2015-11-23" gender="F" nation="BRA" license="393260" swrid="5616446" athleteid="2510" externalid="393260">
              <RESULTS>
                <RESULT eventid="1092" points="41" swimtime="00:02:25.55" resultid="2511" heatid="3437" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:09.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="52" swimtime="00:01:15.59" resultid="2512" heatid="3400" lane="5" entrytime="00:01:12.03" entrycourse="SCM" />
                <RESULT eventid="1108" points="39" swimtime="00:01:11.43" resultid="2513" heatid="3452" lane="5" />
                <RESULT eventid="1128" points="52" swimtime="00:01:01.13" resultid="2514" heatid="3467" lane="2" entrytime="00:01:08.10" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Kraemer Geremia" birthdate="2013-08-16" gender="M" nation="BRA" license="377041" swrid="5588762" athleteid="2307" externalid="377041">
              <RESULTS>
                <RESULT eventid="1089" points="199" swimtime="00:02:50.10" resultid="2308" heatid="3433" lane="3" entrytime="00:02:51.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                    <SPLIT distance="100" swimtime="00:01:20.74" />
                    <SPLIT distance="150" swimtime="00:02:05.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="161" swimtime="00:01:41.43" resultid="2309" heatid="3396" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="177" swimtime="00:01:27.62" resultid="2310" heatid="3451" lane="3" entrytime="00:01:30.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="235" swimtime="00:00:32.64" resultid="2311" heatid="3487" lane="6" entrytime="00:00:33.70" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="LIV" lastname="Carvalho" birthdate="2011-09-13" gender="F" nation="BRA" license="366899" swrid="5602524" athleteid="1992" externalid="366899">
              <RESULTS>
                <RESULT eventid="1144" points="282" swimtime="00:05:52.36" resultid="1993" heatid="3492" lane="2" entrytime="00:06:42.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="100" swimtime="00:01:20.81" />
                    <SPLIT distance="150" swimtime="00:02:06.07" />
                    <SPLIT distance="200" swimtime="00:02:51.78" />
                    <SPLIT distance="250" swimtime="00:03:36.99" />
                    <SPLIT distance="300" swimtime="00:04:22.32" />
                    <SPLIT distance="350" swimtime="00:05:07.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="266" swimtime="00:01:36.88" resultid="1994" heatid="3502" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="225" swimtime="00:03:20.20" resultid="1995" heatid="3553" lane="6" entrytime="00:03:30.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.59" />
                    <SPLIT distance="100" swimtime="00:01:42.36" />
                    <SPLIT distance="150" swimtime="00:02:36.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="120" swimtime="00:01:49.45" resultid="1996" heatid="3594" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="269" swimtime="00:01:17.77" resultid="1997" heatid="3565" lane="5" entrytime="00:01:21.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Moreira Pasqual" birthdate="2014-07-09" gender="M" nation="BRA" license="382125" swrid="5602562" athleteid="2378" externalid="382125">
              <RESULTS>
                <RESULT eventid="1095" points="119" swimtime="00:01:31.14" resultid="2379" heatid="3442" lane="8" entrytime="00:01:52.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="108" swimtime="00:00:46.42" resultid="2380" heatid="3423" lane="3" entrytime="00:00:48.39" entrycourse="SCM" />
                <RESULT eventid="1111" points="118" swimtime="00:00:44.32" resultid="2381" heatid="3459" lane="3" entrytime="00:00:49.15" entrycourse="SCM" />
                <RESULT eventid="1131" points="139" swimtime="00:00:38.83" resultid="2382" heatid="3473" lane="3" entrytime="00:00:43.76" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="De Lima Cavalcanti" birthdate="2014-10-07" gender="M" nation="BRA" license="385884" swrid="5684550" athleteid="2613" externalid="385884">
              <RESULTS>
                <RESULT eventid="1095" points="99" swimtime="00:01:36.64" resultid="2614" heatid="3442" lane="5" entrytime="00:01:24.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="136" swimtime="00:00:42.97" resultid="2615" heatid="3423" lane="4" entrytime="00:00:41.45" entrycourse="SCM" />
                <RESULT eventid="1111" points="45" swimtime="00:01:00.74" resultid="2616" heatid="3459" lane="6" entrytime="00:00:49.23" entrycourse="SCM" />
                <RESULT eventid="1131" points="120" swimtime="00:00:40.86" resultid="2617" heatid="3474" lane="5" entrytime="00:00:38.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Filipa" lastname="Saboia Ruiz" birthdate="2013-04-05" gender="F" nation="BRA" license="376976" swrid="5588894" athleteid="2258" externalid="376976">
              <RESULTS>
                <RESULT eventid="1086" points="131" swimtime="00:03:36.75" resultid="2259" heatid="3425" lane="5" entrytime="00:03:36.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.83" />
                    <SPLIT distance="100" swimtime="00:01:47.48" />
                    <SPLIT distance="150" swimtime="00:02:45.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="144" swimtime="00:00:48.14" resultid="2260" heatid="3408" lane="3" entrytime="00:00:52.01" entrycourse="SCM" />
                <RESULT eventid="1102" status="DNS" swimtime="00:00:00.00" resultid="2261" heatid="3446" lane="6" entrytime="00:01:59.74" entrycourse="SCM" />
                <RESULT eventid="1138" status="DNS" swimtime="00:00:00.00" resultid="2262" heatid="3478" lane="6" entrytime="00:00:45.58" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Prosdocimo" birthdate="2010-11-23" gender="F" nation="BRA" license="356251" swrid="5600238" athleteid="1892" externalid="356251">
              <RESULTS>
                <RESULT eventid="1144" points="444" swimtime="00:05:03.13" resultid="1893" heatid="3494" lane="8" entrytime="00:05:15.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:10.69" />
                    <SPLIT distance="150" swimtime="00:01:49.27" />
                    <SPLIT distance="200" swimtime="00:02:28.50" />
                    <SPLIT distance="250" swimtime="00:03:07.62" />
                    <SPLIT distance="300" swimtime="00:03:46.93" />
                    <SPLIT distance="350" swimtime="00:04:25.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="362" reactiontime="+69" swimtime="00:01:16.98" resultid="1894" heatid="3526" lane="5" entrytime="00:01:18.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="313" swimtime="00:02:59.43" resultid="1895" heatid="3554" lane="5" entrytime="00:03:00.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.12" />
                    <SPLIT distance="100" swimtime="00:01:25.11" />
                    <SPLIT distance="150" swimtime="00:02:22.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="397" swimtime="00:20:35.38" resultid="1896" heatid="3582" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.79" />
                    <SPLIT distance="100" swimtime="00:01:17.56" />
                    <SPLIT distance="150" swimtime="00:01:58.31" />
                    <SPLIT distance="200" swimtime="00:02:39.62" />
                    <SPLIT distance="250" swimtime="00:03:21.09" />
                    <SPLIT distance="300" swimtime="00:04:02.50" />
                    <SPLIT distance="350" swimtime="00:04:44.40" />
                    <SPLIT distance="400" swimtime="00:05:25.42" />
                    <SPLIT distance="450" swimtime="00:06:06.83" />
                    <SPLIT distance="500" swimtime="00:06:48.40" />
                    <SPLIT distance="550" swimtime="00:07:29.71" />
                    <SPLIT distance="600" swimtime="00:08:10.89" />
                    <SPLIT distance="650" swimtime="00:08:51.64" />
                    <SPLIT distance="700" swimtime="00:09:32.67" />
                    <SPLIT distance="750" swimtime="00:10:13.90" />
                    <SPLIT distance="800" swimtime="00:10:55.32" />
                    <SPLIT distance="850" swimtime="00:11:36.88" />
                    <SPLIT distance="900" swimtime="00:12:18.13" />
                    <SPLIT distance="950" swimtime="00:12:59.47" />
                    <SPLIT distance="1000" swimtime="00:13:40.99" />
                    <SPLIT distance="1050" swimtime="00:14:22.77" />
                    <SPLIT distance="1100" swimtime="00:15:04.84" />
                    <SPLIT distance="1150" swimtime="00:15:46.65" />
                    <SPLIT distance="1200" swimtime="00:16:28.20" />
                    <SPLIT distance="1250" swimtime="00:17:09.81" />
                    <SPLIT distance="1300" swimtime="00:17:51.22" />
                    <SPLIT distance="1350" swimtime="00:18:32.53" />
                    <SPLIT distance="1400" swimtime="00:19:13.95" />
                    <SPLIT distance="1450" swimtime="00:19:55.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="421" swimtime="00:01:07.00" resultid="1897" heatid="3568" lane="4" entrytime="00:01:08.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joana" lastname="Asinelli Casagrande" birthdate="2013-10-26" gender="F" nation="BRA" license="376970" swrid="5588536" athleteid="2240" externalid="376970">
              <RESULTS>
                <RESULT eventid="1086" points="189" swimtime="00:03:12.18" resultid="2241" heatid="3426" lane="2" entrytime="00:03:17.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.18" />
                    <SPLIT distance="100" swimtime="00:01:33.66" />
                    <SPLIT distance="150" swimtime="00:02:24.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="222" reactiontime="+69" swimtime="00:00:41.64" resultid="2242" heatid="3409" lane="4" entrytime="00:00:43.60" entrycourse="SCM" />
                <RESULT eventid="1102" points="199" swimtime="00:01:36.66" resultid="2243" heatid="3447" lane="7" entrytime="00:01:42.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1118" points="125" swimtime="00:01:47.93" resultid="2244" heatid="3461" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Moreira Segadaes" birthdate="2008-05-15" gender="M" nation="BRA" license="331574" swrid="5600220" athleteid="1762" externalid="331574">
              <RESULTS>
                <RESULT eventid="1168" points="546" swimtime="00:01:07.60" resultid="1763" heatid="3513" lane="1" entrytime="00:01:09.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="531" swimtime="00:00:30.80" resultid="1764" heatid="3612" lane="7" entrytime="00:00:31.60" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Geremia" birthdate="2011-07-20" gender="F" nation="BRA" license="366908" swrid="5602543" athleteid="2028" externalid="366908">
              <RESULTS>
                <RESULT eventid="1144" points="450" swimtime="00:05:01.80" resultid="2029" heatid="3493" lane="4" entrytime="00:05:18.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                    <SPLIT distance="100" swimtime="00:01:11.16" />
                    <SPLIT distance="150" swimtime="00:01:49.55" />
                    <SPLIT distance="200" swimtime="00:02:28.82" />
                    <SPLIT distance="250" swimtime="00:03:07.79" />
                    <SPLIT distance="300" swimtime="00:03:46.32" />
                    <SPLIT distance="350" swimtime="00:04:24.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="379" reactiontime="+68" swimtime="00:01:15.83" resultid="2030" heatid="3526" lane="7" entrytime="00:01:20.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="291" swimtime="00:01:34.00" resultid="2031" heatid="3505" lane="8" entrytime="00:01:32.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="399" swimtime="00:02:45.47" resultid="2032" heatid="3555" lane="6" entrytime="00:02:53.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.38" />
                    <SPLIT distance="100" swimtime="00:01:21.71" />
                    <SPLIT distance="150" swimtime="00:02:09.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="438" swimtime="00:01:06.15" resultid="2033" heatid="3568" lane="3" entrytime="00:01:08.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Rocha Silva" birthdate="2007-10-10" gender="M" nation="BRA" license="372280" athleteid="1795" externalid="372280">
              <RESULTS>
                <RESULT eventid="1152" points="638" swimtime="00:04:06.45" resultid="1796" heatid="3497" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.88" />
                    <SPLIT distance="100" swimtime="00:00:58.68" />
                    <SPLIT distance="150" swimtime="00:01:29.44" />
                    <SPLIT distance="200" swimtime="00:02:00.89" />
                    <SPLIT distance="250" swimtime="00:02:32.05" />
                    <SPLIT distance="300" swimtime="00:03:04.49" />
                    <SPLIT distance="350" swimtime="00:03:36.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="622" swimtime="00:00:23.61" resultid="1797" heatid="3550" lane="5" entrytime="00:00:24.40" entrycourse="SCM" />
                <RESULT eventid="1248" points="692" swimtime="00:00:50.69" resultid="1798" heatid="3581" lane="6" entrytime="00:00:52.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Heloisa Souza" birthdate="2007-01-15" gender="F" nation="BRA" license="336615" swrid="5600184" athleteid="1792" externalid="336615">
              <RESULTS>
                <RESULT eventid="1144" points="610" swimtime="00:04:32.60" resultid="1793" heatid="3494" lane="1" entrytime="00:04:49.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:05.01" />
                    <SPLIT distance="150" swimtime="00:01:38.63" />
                    <SPLIT distance="200" swimtime="00:02:13.36" />
                    <SPLIT distance="250" swimtime="00:02:48.13" />
                    <SPLIT distance="300" swimtime="00:03:22.94" />
                    <SPLIT distance="350" swimtime="00:03:57.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="585" swimtime="00:01:00.05" resultid="1794" heatid="3570" lane="5" entrytime="00:01:00.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Morais Shibata" birthdate="2014-02-09" gender="M" nation="BRA" license="391018" swrid="5602561" athleteid="2446" externalid="391018">
              <RESULTS>
                <RESULT eventid="1095" points="99" swimtime="00:01:36.62" resultid="2447" heatid="3441" lane="2" entrytime="00:02:17.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" status="DNS" swimtime="00:00:00.00" resultid="2448" heatid="3423" lane="1" entrytime="00:00:54.55" entrycourse="SCM" />
                <RESULT eventid="1111" points="75" swimtime="00:00:51.40" resultid="2449" heatid="3459" lane="1" entrytime="00:00:56.99" entrycourse="SCM" />
                <RESULT eventid="1131" points="117" swimtime="00:00:41.20" resultid="2450" heatid="3473" lane="4" entrytime="00:00:43.13" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Wolff Contin" birthdate="2015-10-10" gender="M" nation="BRA" license="406745" athleteid="2656" externalid="406745">
              <RESULTS>
                <RESULT eventid="1083" points="34" reactiontime="+56" swimtime="00:01:07.72" resultid="2657" heatid="3421" lane="2" />
                <RESULT eventid="1071" points="22" swimtime="00:01:28.47" resultid="2658" heatid="3403" lane="8" />
                <RESULT eventid="1111" points="12" swimtime="00:01:33.37" resultid="2659" heatid="3457" lane="3" />
                <RESULT eventid="1131" points="33" swimtime="00:01:02.31" resultid="2660" heatid="3470" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Garcia" birthdate="2015-10-26" gender="M" nation="BRA" license="406967" athleteid="2732" externalid="406967">
              <RESULTS>
                <RESULT eventid="1083" points="25" reactiontime="+81" swimtime="00:01:15.52" resultid="2733" heatid="3420" lane="6" />
                <RESULT eventid="1071" points="18" swimtime="00:01:34.42" resultid="2734" heatid="3402" lane="3" />
                <RESULT eventid="1111" points="14" swimtime="00:01:29.25" resultid="2735" heatid="3456" lane="7" />
                <RESULT eventid="1131" points="18" swimtime="00:01:16.80" resultid="2736" heatid="3470" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Magalhaes Dos Reis" birthdate="2010-05-05" gender="M" nation="BRA" license="356361" swrid="5600207" athleteid="1928" externalid="356361">
              <RESULTS>
                <RESULT eventid="1168" points="341" swimtime="00:01:19.06" resultid="1929" heatid="3511" lane="6" entrytime="00:01:24.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="382" swimtime="00:00:27.78" resultid="1930" heatid="3542" lane="5" />
                <RESULT eventid="1232" points="325" swimtime="00:02:39.39" resultid="1931" heatid="3559" lane="4" entrytime="00:02:49.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                    <SPLIT distance="100" swimtime="00:01:15.61" />
                    <SPLIT distance="150" swimtime="00:02:04.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="251" swimtime="00:01:15.71" resultid="1932" heatid="3599" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="375" swimtime="00:01:02.14" resultid="1933" heatid="3571" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Peret Saboia" birthdate="2009-11-25" gender="F" nation="BRA" license="342238" swrid="5600234" athleteid="1838" externalid="342238">
              <RESULTS>
                <RESULT eventid="1160" points="434" swimtime="00:01:22.34" resultid="1839" heatid="3505" lane="5" entrytime="00:01:24.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="369" swimtime="00:02:49.78" resultid="1840" heatid="3555" lane="3" entrytime="00:02:51.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.96" />
                    <SPLIT distance="100" swimtime="00:01:23.83" />
                    <SPLIT distance="150" swimtime="00:02:10.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="426" swimtime="00:00:37.68" resultid="1841" heatid="3605" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Sieczkowski Pacheco" birthdate="2015-11-20" gender="F" nation="BRA" license="393261" swrid="5616450" athleteid="2515" externalid="393261">
              <RESULTS>
                <RESULT eventid="1092" points="81" swimtime="00:01:55.92" resultid="2516" heatid="3435" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="113" swimtime="00:00:58.63" resultid="2517" heatid="3401" lane="7" entrytime="00:01:01.66" entrycourse="SCM" />
                <RESULT eventid="1108" points="61" swimtime="00:01:01.63" resultid="2518" heatid="3454" lane="1" />
                <RESULT eventid="1128" points="90" swimtime="00:00:50.99" resultid="2519" heatid="3468" lane="1" entrytime="00:00:51.61" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Martynychen" birthdate="2011-12-19" gender="M" nation="BRA" license="366893" swrid="5602557" athleteid="1974" externalid="366893">
              <RESULTS>
                <RESULT eventid="1200" points="204" reactiontime="+104" swimtime="00:01:22.08" resultid="1975" heatid="3530" lane="2" entrytime="00:01:24.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="344" swimtime="00:05:02.67" resultid="1976" heatid="3499" lane="2" entrytime="00:05:27.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:11.74" />
                    <SPLIT distance="150" swimtime="00:01:50.42" />
                    <SPLIT distance="200" swimtime="00:02:28.97" />
                    <SPLIT distance="250" swimtime="00:03:07.88" />
                    <SPLIT distance="300" swimtime="00:03:46.00" />
                    <SPLIT distance="350" swimtime="00:04:25.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="225" swimtime="00:00:33.14" resultid="1977" heatid="3544" lane="4" entrytime="00:00:33.53" entrycourse="SCM" />
                <RESULT eventid="1264" points="368" swimtime="00:19:40.88" resultid="1978" heatid="3584" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:15.87" />
                    <SPLIT distance="150" swimtime="00:01:56.48" />
                    <SPLIT distance="200" swimtime="00:02:35.25" />
                    <SPLIT distance="250" swimtime="00:03:14.56" />
                    <SPLIT distance="300" swimtime="00:03:54.21" />
                    <SPLIT distance="350" swimtime="00:04:33.75" />
                    <SPLIT distance="400" swimtime="00:05:12.83" />
                    <SPLIT distance="450" swimtime="00:05:52.13" />
                    <SPLIT distance="500" swimtime="00:06:31.66" />
                    <SPLIT distance="550" swimtime="00:07:11.29" />
                    <SPLIT distance="600" swimtime="00:07:51.70" />
                    <SPLIT distance="650" swimtime="00:08:31.28" />
                    <SPLIT distance="700" swimtime="00:09:10.80" />
                    <SPLIT distance="750" swimtime="00:09:50.60" />
                    <SPLIT distance="800" swimtime="00:10:30.96" />
                    <SPLIT distance="850" swimtime="00:11:10.57" />
                    <SPLIT distance="900" swimtime="00:11:50.62" />
                    <SPLIT distance="950" swimtime="00:12:31.02" />
                    <SPLIT distance="1000" swimtime="00:13:10.60" />
                    <SPLIT distance="1050" swimtime="00:13:50.02" />
                    <SPLIT distance="1100" swimtime="00:14:29.31" />
                    <SPLIT distance="1150" swimtime="00:15:08.53" />
                    <SPLIT distance="1200" swimtime="00:15:49.00" />
                    <SPLIT distance="1250" swimtime="00:16:27.46" />
                    <SPLIT distance="1300" swimtime="00:17:06.70" />
                    <SPLIT distance="1350" swimtime="00:17:46.70" />
                    <SPLIT distance="1400" swimtime="00:18:26.90" />
                    <SPLIT distance="1450" swimtime="00:19:05.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="252" swimtime="00:01:10.91" resultid="1979" heatid="3576" lane="2" entrytime="00:01:12.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Rocha" birthdate="2011-08-25" gender="F" nation="BRA" license="366904" swrid="5602578" athleteid="2010" externalid="366904">
              <RESULTS>
                <RESULT eventid="1144" points="417" swimtime="00:05:09.44" resultid="2011" heatid="3493" lane="3" entrytime="00:05:20.59" entrycourse="SCM" />
                <RESULT eventid="1192" points="346" reactiontime="+69" swimtime="00:01:18.12" resultid="2012" heatid="3526" lane="3" entrytime="00:01:19.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="266" swimtime="00:01:36.95" resultid="2013" heatid="3504" lane="8" entrytime="00:01:43.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="335" swimtime="00:02:55.29" resultid="2014" heatid="3554" lane="2" entrytime="00:03:04.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                    <SPLIT distance="100" swimtime="00:01:23.95" />
                    <SPLIT distance="150" swimtime="00:02:17.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="395" swimtime="00:01:08.48" resultid="2015" heatid="3568" lane="6" entrytime="00:01:09.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Ribas Luz" birthdate="2015-02-05" gender="F" nation="BRA" license="406743" athleteid="2648" externalid="406743">
              <RESULTS>
                <RESULT eventid="1080" points="43" swimtime="00:01:11.89" resultid="2649" heatid="3417" lane="2" />
                <RESULT eventid="1068" points="30" swimtime="00:01:30.45" resultid="2650" heatid="3399" lane="2" />
                <RESULT eventid="1108" points="15" swimtime="00:01:37.59" resultid="2651" heatid="3453" lane="7" />
                <RESULT eventid="1128" points="42" swimtime="00:01:05.73" resultid="2652" heatid="3465" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Zagonel Krempel" birthdate="2015-07-27" gender="F" nation="BRA" license="406962" athleteid="2724" externalid="406962">
              <RESULTS>
                <RESULT eventid="1080" points="44" swimtime="00:01:11.43" resultid="2725" heatid="3417" lane="5" />
                <RESULT eventid="1068" points="55" swimtime="00:01:14.49" resultid="2726" heatid="3400" lane="6" />
                <RESULT eventid="1128" points="39" swimtime="00:01:07.49" resultid="2727" heatid="3466" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Cipriani Presiazniuk" birthdate="2012-07-03" gender="M" nation="BRA" license="369267" swrid="5588594" athleteid="2085" externalid="369267">
              <RESULTS>
                <RESULT eventid="1089" points="211" swimtime="00:02:46.77" resultid="2086" heatid="3429" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                    <SPLIT distance="100" swimtime="00:01:22.32" />
                    <SPLIT distance="150" swimtime="00:02:06.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="185" reactiontime="+80" swimtime="00:00:38.76" resultid="2087" heatid="3415" lane="3" entrytime="00:00:38.27" entrycourse="SCM" />
                <RESULT eventid="1105" points="176" swimtime="00:01:27.90" resultid="2088" heatid="3449" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="230" swimtime="00:00:32.90" resultid="2089" heatid="3487" lane="5" entrytime="00:00:33.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Araujo Barros" birthdate="2008-12-26" gender="M" nation="BRA" license="331713" swrid="5367497" athleteid="2055" externalid="331713">
              <RESULTS>
                <RESULT eventid="1152" points="600" swimtime="00:04:11.61" resultid="2056" heatid="3501" lane="3" entrytime="00:04:26.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                    <SPLIT distance="100" swimtime="00:01:00.35" />
                    <SPLIT distance="150" swimtime="00:01:32.65" />
                    <SPLIT distance="200" swimtime="00:02:03.92" />
                    <SPLIT distance="250" swimtime="00:02:36.22" />
                    <SPLIT distance="300" swimtime="00:03:08.36" />
                    <SPLIT distance="350" swimtime="00:03:40.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="494" swimtime="00:00:25.50" resultid="2057" heatid="3543" lane="7" />
                <RESULT eventid="1296" points="463" swimtime="00:01:01.75" resultid="2058" heatid="3599" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="578" swimtime="00:00:53.80" resultid="2059" heatid="3571" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Fantin Dias De Andrade" birthdate="2010-11-06" gender="F" nation="BRA" license="339262" swrid="5588684" athleteid="2176" externalid="339262">
              <RESULTS>
                <RESULT eventid="1192" points="233" reactiontime="+59" swimtime="00:01:29.16" resultid="2177" heatid="3524" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="301" swimtime="00:01:32.96" resultid="2178" heatid="3504" lane="2" entrytime="00:01:36.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" status="DSQ" swimtime="00:03:02.83" resultid="2179" heatid="3554" lane="3" entrytime="00:03:00.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                    <SPLIT distance="100" swimtime="00:01:29.46" />
                    <SPLIT distance="150" swimtime="00:02:23.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="202" swimtime="00:01:32.06" resultid="2180" heatid="3594" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="313" swimtime="00:01:13.94" resultid="2181" heatid="3566" lane="1" entrytime="00:01:15.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Albuquerque" birthdate="2012-08-17" gender="F" nation="BRA" license="369275" swrid="5602507" athleteid="2115" externalid="369275">
              <RESULTS>
                <RESULT eventid="1062" points="393" swimtime="00:01:25.13" resultid="2116" heatid="3394" lane="4" entrytime="00:01:32.18" entrycourse="SCM" />
                <RESULT eventid="1086" points="234" swimtime="00:02:58.83" resultid="2117" heatid="3426" lane="5" entrytime="00:03:05.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.66" />
                    <SPLIT distance="100" swimtime="00:01:24.81" />
                    <SPLIT distance="150" swimtime="00:02:11.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="273" swimtime="00:01:27.11" resultid="2118" heatid="3445" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="296" swimtime="00:00:34.37" resultid="2119" heatid="3480" lane="5" entrytime="00:00:35.49" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Lauand Lorenci" birthdate="2013-03-06" gender="M" nation="BRA" license="376982" swrid="5588764" athleteid="2281" externalid="376982">
              <RESULTS>
                <RESULT eventid="1089" points="178" swimtime="00:02:56.59" resultid="2282" heatid="3431" lane="3" entrytime="00:03:23.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                    <SPLIT distance="100" swimtime="00:01:27.32" />
                    <SPLIT distance="150" swimtime="00:02:13.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="191" swimtime="00:01:35.88" resultid="2283" heatid="3396" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="174" swimtime="00:01:28.15" resultid="2284" heatid="3451" lane="6" entrytime="00:01:33.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="195" swimtime="00:00:34.73" resultid="2285" heatid="3486" lane="1" entrytime="00:00:36.44" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Carneiro Silva" birthdate="2011-02-21" gender="F" nation="BRA" license="390924" swrid="5602522" athleteid="2594" externalid="390924">
              <RESULTS>
                <RESULT eventid="1144" points="334" swimtime="00:05:33.26" resultid="2595" heatid="3491" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.81" />
                    <SPLIT distance="100" swimtime="00:01:15.24" />
                    <SPLIT distance="150" swimtime="00:01:57.31" />
                    <SPLIT distance="200" swimtime="00:02:40.18" />
                    <SPLIT distance="250" swimtime="00:03:23.31" />
                    <SPLIT distance="300" swimtime="00:04:06.57" />
                    <SPLIT distance="350" swimtime="00:04:49.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="291" reactiontime="+89" swimtime="00:01:22.80" resultid="2596" heatid="3525" lane="4" entrytime="00:01:22.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="230" swimtime="00:01:41.67" resultid="2597" heatid="3502" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="276" swimtime="00:03:07.02" resultid="2598" heatid="3553" lane="3" entrytime="00:03:12.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.22" />
                    <SPLIT distance="100" swimtime="00:01:28.90" />
                    <SPLIT distance="150" swimtime="00:02:25.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="324" swimtime="00:01:13.16" resultid="2599" heatid="3567" lane="1" entrytime="00:01:12.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Taborda Ribas" birthdate="2015-12-30" gender="M" nation="BRA" license="406748" athleteid="2670" externalid="406748">
              <RESULTS>
                <RESULT eventid="1083" points="29" reactiontime="+70" swimtime="00:01:11.96" resultid="2671" heatid="3421" lane="6" />
                <RESULT eventid="1071" points="28" swimtime="00:01:21.49" resultid="2672" heatid="3402" lane="7" />
                <RESULT eventid="1111" points="15" swimtime="00:01:26.45" resultid="2673" heatid="3458" lane="2" />
                <RESULT eventid="1131" points="41" swimtime="00:00:58.00" resultid="2674" heatid="3470" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Szpak De Vasconcelos" birthdate="2012-06-29" gender="M" nation="BRA" license="369271" swrid="5588928" athleteid="2100" externalid="369271">
              <RESULTS>
                <RESULT eventid="1077" points="231" reactiontime="+69" swimtime="00:00:36.02" resultid="2101" heatid="3412" lane="4" />
                <RESULT eventid="1065" points="277" swimtime="00:01:24.75" resultid="2102" heatid="3398" lane="4" entrytime="00:01:26.42" entrycourse="SCM" />
                <RESULT eventid="1105" points="233" swimtime="00:01:20.01" resultid="2103" heatid="3451" lane="4" entrytime="00:01:20.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="293" swimtime="00:00:30.35" resultid="2104" heatid="3488" lane="4" entrytime="00:00:30.37" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Presiazniuk" birthdate="2010-10-14" gender="M" nation="BRA" license="356353" swrid="5600237" athleteid="1910" externalid="356353">
              <RESULTS>
                <RESULT eventid="1200" points="354" reactiontime="+67" swimtime="00:01:08.29" resultid="1911" heatid="3531" lane="1" entrytime="00:01:15.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="431" swimtime="00:04:40.81" resultid="1912" heatid="3497" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                    <SPLIT distance="100" swimtime="00:01:06.11" />
                    <SPLIT distance="150" swimtime="00:01:41.64" />
                    <SPLIT distance="200" swimtime="00:02:17.32" />
                    <SPLIT distance="250" swimtime="00:02:53.53" />
                    <SPLIT distance="300" swimtime="00:03:29.50" />
                    <SPLIT distance="350" swimtime="00:04:05.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="326" swimtime="00:02:39.19" resultid="1913" heatid="3559" lane="6" entrytime="00:02:57.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:01:15.76" />
                    <SPLIT distance="150" swimtime="00:02:05.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="332" swimtime="00:00:31.92" resultid="1914" heatid="3593" lane="8" entrytime="00:00:35.03" entrycourse="SCM" />
                <RESULT eventid="1248" points="417" swimtime="00:01:00.01" resultid="1915" heatid="3577" lane="4" entrytime="00:01:05.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Antunes Luzzi" birthdate="2014-02-14" gender="M" nation="BRA" license="391019" swrid="5602510" athleteid="2451" externalid="391019">
              <RESULTS>
                <RESULT eventid="1083" points="32" swimtime="00:01:09.06" resultid="2452" heatid="3422" lane="5" entrytime="00:01:05.37" entrycourse="SCM" />
                <RESULT eventid="1071" points="47" swimtime="00:01:08.68" resultid="2453" heatid="3403" lane="5" entrytime="00:01:08.73" entrycourse="SCM" />
                <RESULT eventid="1111" points="12" swimtime="00:01:34.31" resultid="2454" heatid="3456" lane="6" />
                <RESULT eventid="1131" points="26" swimtime="00:01:07.31" resultid="2455" heatid="3472" lane="1" entrytime="00:01:05.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Stramandinoli Zanicotti" birthdate="2013-06-18" gender="F" nation="BRA" license="376967" swrid="5588924" athleteid="2225" externalid="376967">
              <RESULTS>
                <RESULT eventid="1062" points="104" swimtime="00:02:12.33" resultid="2226" heatid="3392" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1086" points="103" swimtime="00:03:55.06" resultid="2227" heatid="3425" lane="2" entrytime="00:04:38.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.12" />
                    <SPLIT distance="100" swimtime="00:01:57.77" />
                    <SPLIT distance="150" swimtime="00:03:00.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="99" swimtime="00:02:01.88" resultid="2228" heatid="3444" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="122" swimtime="00:00:46.20" resultid="2229" heatid="3478" lane="1" entrytime="00:00:48.17" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Antunes Saboia" birthdate="2012-06-28" gender="M" nation="BRA" license="369278" swrid="5602511" athleteid="2130" externalid="369278">
              <RESULTS>
                <RESULT eventid="1077" points="152" reactiontime="+78" swimtime="00:00:41.34" resultid="2131" heatid="3412" lane="7" />
                <RESULT eventid="1065" points="229" swimtime="00:01:30.34" resultid="2132" heatid="3398" lane="3" entrytime="00:01:37.45" entrycourse="SCM" />
                <RESULT eventid="1105" points="187" swimtime="00:01:26.10" resultid="2133" heatid="3449" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="237" swimtime="00:00:32.56" resultid="2134" heatid="3487" lane="4" entrytime="00:00:33.12" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Artigas Pinheiro" birthdate="2011-08-25" gender="M" nation="BRA" license="377040" swrid="5588535" athleteid="2301" externalid="377040">
              <RESULTS>
                <RESULT eventid="1200" points="186" reactiontime="+86" swimtime="00:01:24.66" resultid="2302" heatid="3530" lane="7" entrytime="00:01:29.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="218" swimtime="00:01:31.76" resultid="2303" heatid="3510" lane="1" entrytime="00:01:38.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="291" swimtime="00:05:20.17" resultid="2304" heatid="3499" lane="7" entrytime="00:05:27.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.06" />
                    <SPLIT distance="100" swimtime="00:01:18.46" />
                    <SPLIT distance="150" swimtime="00:02:00.36" />
                    <SPLIT distance="200" swimtime="00:02:41.95" />
                    <SPLIT distance="250" swimtime="00:03:21.48" />
                    <SPLIT distance="300" swimtime="00:04:02.15" />
                    <SPLIT distance="350" swimtime="00:04:42.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="175" swimtime="00:01:25.42" resultid="2305" heatid="3598" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="245" swimtime="00:01:11.63" resultid="2306" heatid="3575" lane="4" entrytime="00:01:14.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Gonçalves Sperandio" birthdate="2013-05-22" gender="M" nation="BRA" license="376980" swrid="5588851" athleteid="2271" externalid="376980">
              <RESULTS>
                <RESULT eventid="1089" points="191" swimtime="00:02:52.51" resultid="2272" heatid="3433" lane="5" entrytime="00:02:50.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.69" />
                    <SPLIT distance="100" swimtime="00:01:24.79" />
                    <SPLIT distance="150" swimtime="00:02:09.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="148" swimtime="00:01:44.36" resultid="2273" heatid="3397" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="149" swimtime="00:01:32.93" resultid="2274" heatid="3451" lane="1" entrytime="00:01:41.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="194" swimtime="00:00:34.79" resultid="2275" heatid="3486" lane="2" entrytime="00:00:35.92" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Alzamora Calado" birthdate="2013-04-26" gender="F" nation="BRA" license="376960" swrid="5588522" athleteid="2206" externalid="376960">
              <RESULTS>
                <RESULT eventid="1062" points="163" swimtime="00:01:53.97" resultid="2207" heatid="3393" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1086" points="263" swimtime="00:02:52.11" resultid="2208" heatid="3427" lane="2" entrytime="00:02:54.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                    <SPLIT distance="100" swimtime="00:01:25.14" />
                    <SPLIT distance="150" swimtime="00:02:11.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="258" swimtime="00:01:28.68" resultid="2209" heatid="3447" lane="5" entrytime="00:01:34.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="315" swimtime="00:00:33.68" resultid="2210" heatid="3480" lane="3" entrytime="00:00:35.75" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo" lastname="Gabriel Nascimento" birthdate="2008-11-14" gender="M" nation="BRA" license="348028" swrid="5600171" athleteid="2416" externalid="348028" level="BIG BUM">
              <RESULTS>
                <RESULT eventid="1184" points="455" swimtime="00:00:28.27" resultid="2417" heatid="3522" lane="7" entrytime="00:00:29.27" entrycourse="SCM" />
                <RESULT eventid="1296" points="402" swimtime="00:01:04.71" resultid="2418" heatid="3601" lane="5" entrytime="00:01:04.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Saporiti Salvi" birthdate="2013-06-28" gender="M" nation="BRA" license="377032" swrid="5588896" athleteid="2296" externalid="377032">
              <RESULTS>
                <RESULT eventid="1089" points="187" swimtime="00:02:53.48" resultid="2297" heatid="3433" lane="6" entrytime="00:02:53.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.99" />
                    <SPLIT distance="100" swimtime="00:01:24.77" />
                    <SPLIT distance="150" swimtime="00:02:10.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="137" swimtime="00:01:47.13" resultid="2298" heatid="3396" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" status="DSQ" swimtime="00:01:37.98" resultid="2299" heatid="3463" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="188" swimtime="00:00:35.17" resultid="2300" heatid="3482" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Novak Bredt" birthdate="2009-09-08" gender="F" nation="BRA" license="338909" swrid="5622297" athleteid="1785" externalid="338909">
              <RESULTS>
                <RESULT eventid="1160" points="426" swimtime="00:01:22.87" resultid="1786" heatid="3505" lane="4" entrytime="00:01:22.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="1787" heatid="3556" lane="7" entrytime="00:02:43.49" entrycourse="SCM" />
                <RESULT eventid="1304" status="DNS" swimtime="00:00:00.00" resultid="1788" heatid="3604" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manoela" lastname="Andrade" birthdate="2010-03-10" gender="F" nation="BRA" license="339042" swrid="5363102" athleteid="1946" externalid="339042">
              <RESULTS>
                <RESULT eventid="1144" points="409" swimtime="00:05:11.41" resultid="1947" heatid="3493" lane="2" entrytime="00:05:24.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.77" />
                    <SPLIT distance="100" swimtime="00:01:13.00" />
                    <SPLIT distance="150" swimtime="00:01:52.16" />
                    <SPLIT distance="200" swimtime="00:02:31.66" />
                    <SPLIT distance="250" swimtime="00:03:12.12" />
                    <SPLIT distance="300" swimtime="00:03:51.92" />
                    <SPLIT distance="350" swimtime="00:04:32.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="231" swimtime="00:01:29.34" resultid="1948" heatid="3525" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="283" swimtime="00:03:05.52" resultid="1949" heatid="3554" lane="6" entrytime="00:03:03.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.89" />
                    <SPLIT distance="100" swimtime="00:01:27.42" />
                    <SPLIT distance="150" swimtime="00:02:25.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="275" swimtime="00:01:23.04" resultid="1950" heatid="3595" lane="4" entrytime="00:01:21.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="301" swimtime="00:01:14.91" resultid="1951" heatid="3564" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Cabrera Cirino" birthdate="2011-01-28" gender="M" nation="BRA" license="369531" swrid="5588569" athleteid="2150" externalid="369531">
              <RESULTS>
                <RESULT eventid="1200" points="318" reactiontime="+69" swimtime="00:01:10.77" resultid="2151" heatid="3531" lane="2" entrytime="00:01:12.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="377" swimtime="00:04:53.81" resultid="2152" heatid="3500" lane="1" entrytime="00:05:00.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.37" />
                    <SPLIT distance="100" swimtime="00:01:08.43" />
                    <SPLIT distance="150" swimtime="00:01:45.70" />
                    <SPLIT distance="200" swimtime="00:02:23.74" />
                    <SPLIT distance="250" swimtime="00:03:01.87" />
                    <SPLIT distance="300" swimtime="00:03:40.11" />
                    <SPLIT distance="350" swimtime="00:04:17.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="363" swimtime="00:00:28.24" resultid="2153" heatid="3547" lane="4" entrytime="00:00:27.95" entrycourse="SCM" />
                <RESULT eventid="1296" points="291" swimtime="00:01:12.04" resultid="2154" heatid="3600" lane="5" entrytime="00:01:19.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="378" swimtime="00:01:01.97" resultid="2155" heatid="3578" lane="6" entrytime="00:01:01.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Laurindo Netto" birthdate="2005-07-15" gender="M" nation="BRA" license="289995" swrid="5600198" athleteid="1742" externalid="289995">
              <RESULTS>
                <RESULT eventid="1200" points="484" reactiontime="+70" swimtime="00:01:01.53" resultid="1743" heatid="3528" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="533" swimtime="00:01:08.16" resultid="1744" heatid="3513" lane="6" entrytime="00:01:06.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="572" swimtime="00:02:12.01" resultid="1745" heatid="3561" lane="3" entrytime="00:02:07.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.25" />
                    <SPLIT distance="100" swimtime="00:01:01.90" />
                    <SPLIT distance="150" swimtime="00:01:39.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Yolanda Ferreira" birthdate="2008-03-17" gender="F" nation="BRA" license="358335" swrid="5600276" athleteid="2188" externalid="358335">
              <RESULTS>
                <RESULT eventid="1208" points="468" swimtime="00:00:29.53" resultid="2189" heatid="3533" lane="3" />
                <RESULT eventid="1160" points="479" swimtime="00:01:19.70" resultid="2190" heatid="3506" lane="6" entrytime="00:01:20.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="459" swimtime="00:00:36.77" resultid="2191" heatid="3606" lane="5" entrytime="00:00:37.48" entrycourse="SCM" />
                <RESULT eventid="1240" points="491" swimtime="00:01:03.67" resultid="2192" heatid="3569" lane="4" entrytime="00:01:05.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="David Cella" birthdate="2008-02-17" gender="M" nation="BRA" license="341107" swrid="5634581" athleteid="2606" externalid="341107">
              <RESULTS>
                <RESULT eventid="1216" points="553" swimtime="00:00:24.55" resultid="2607" heatid="3550" lane="6" entrytime="00:00:24.49" entrycourse="SCM" />
                <RESULT eventid="1312" points="549" swimtime="00:00:30.47" resultid="2608" heatid="3612" lane="6" entrytime="00:00:30.75" entrycourse="SCM" />
                <RESULT eventid="1248" points="548" swimtime="00:00:54.79" resultid="2609" heatid="3581" lane="8" entrytime="00:00:54.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Bernardi Pedrosa" birthdate="2013-03-09" gender="F" nation="BRA" license="376977" swrid="5588551" athleteid="2263" externalid="376977">
              <RESULTS>
                <RESULT eventid="1086" points="182" swimtime="00:03:14.57" resultid="2264" heatid="3426" lane="7" entrytime="00:03:26.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                    <SPLIT distance="100" swimtime="00:01:33.60" />
                    <SPLIT distance="150" swimtime="00:02:25.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="150" reactiontime="+70" swimtime="00:00:47.46" resultid="2265" heatid="3408" lane="2" entrytime="00:00:53.65" entrycourse="SCM" />
                <RESULT eventid="1102" points="172" swimtime="00:01:41.48" resultid="2266" heatid="3446" lane="5" entrytime="00:01:54.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="196" swimtime="00:00:39.41" resultid="2267" heatid="3478" lane="4" entrytime="00:00:43.87" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raphael" lastname="Rached Windmuller" birthdate="2003-05-19" gender="M" nation="BRA" license="249770" swrid="5302329" athleteid="1803" externalid="249770">
              <RESULTS>
                <RESULT eventid="1168" points="803" swimtime="00:00:59.47" resultid="1804" heatid="3508" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="714" swimtime="00:00:27.91" resultid="1805" heatid="3607" lane="6" />
                <RESULT eventid="1248" points="633" swimtime="00:00:52.22" resultid="1806" heatid="3572" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ferreira Motta" birthdate="2008-10-24" gender="M" nation="BRA" license="378068" swrid="5600160" athleteid="2357" externalid="378068">
              <RESULTS>
                <RESULT eventid="1168" points="442" swimtime="00:01:12.54" resultid="2358" heatid="3512" lane="1" entrytime="00:01:20.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="371" swimtime="00:00:28.04" resultid="2359" heatid="3546" lane="4" entrytime="00:00:28.88" entrycourse="SCM" />
                <RESULT eventid="1312" points="431" swimtime="00:00:33.03" resultid="2360" heatid="3607" lane="5" />
                <RESULT eventid="1248" points="407" swimtime="00:01:00.46" resultid="2361" heatid="3578" lane="2" entrytime="00:01:03.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Nishimura Ramina" birthdate="2013-11-25" gender="M" nation="BRA" license="376989" swrid="5588831" athleteid="2327" externalid="376989">
              <RESULTS>
                <RESULT eventid="1089" points="116" swimtime="00:03:23.57" resultid="2328" heatid="3431" lane="8" entrytime="00:03:48.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.87" />
                    <SPLIT distance="100" swimtime="00:01:36.38" />
                    <SPLIT distance="150" swimtime="00:02:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="91" swimtime="00:02:02.73" resultid="2329" heatid="3395" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="86" swimtime="00:01:51.33" resultid="2330" heatid="3450" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="107" swimtime="00:00:42.35" resultid="2331" heatid="3484" lane="1" entrytime="00:00:44.25" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Saboia" birthdate="2009-01-25" gender="M" nation="BRA" license="342252" swrid="5600253" athleteid="1846" externalid="342252">
              <RESULTS>
                <RESULT eventid="1168" points="406" swimtime="00:01:14.60" resultid="1847" heatid="3511" lane="2" entrytime="00:01:24.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="352" swimtime="00:02:35.22" resultid="1848" heatid="3560" lane="1" entrytime="00:02:44.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                    <SPLIT distance="100" swimtime="00:01:15.84" />
                    <SPLIT distance="150" swimtime="00:01:59.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="390" swimtime="00:00:34.14" resultid="1849" heatid="3608" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ravi" lastname="Osternack Erbe" birthdate="2013-08-10" gender="M" nation="BRA" license="372681" swrid="5588841" athleteid="2161" externalid="372681">
              <RESULTS>
                <RESULT eventid="1089" points="187" swimtime="00:02:53.57" resultid="2162" heatid="3433" lane="7" entrytime="00:02:54.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.94" />
                    <SPLIT distance="100" swimtime="00:01:23.06" />
                    <SPLIT distance="150" swimtime="00:02:06.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="163" swimtime="00:00:40.46" resultid="2163" heatid="3415" lane="8" entrytime="00:00:40.92" entrycourse="SCM" />
                <RESULT eventid="1121" points="122" swimtime="00:01:36.19" resultid="2164" heatid="3463" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="198" swimtime="00:00:34.54" resultid="2165" heatid="3486" lane="3" entrytime="00:00:35.59" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Artigas Pinheiro" birthdate="2013-07-31" gender="F" nation="BRA" license="377153" swrid="5588534" athleteid="2352" externalid="377153">
              <RESULTS>
                <RESULT eventid="1086" points="214" swimtime="00:03:04.41" resultid="2353" heatid="3426" lane="6" entrytime="00:03:15.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.65" />
                    <SPLIT distance="100" swimtime="00:01:28.91" />
                    <SPLIT distance="150" swimtime="00:02:17.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="195" reactiontime="+73" swimtime="00:00:43.50" resultid="2354" heatid="3409" lane="2" entrytime="00:00:47.07" entrycourse="SCM" />
                <RESULT eventid="1102" points="167" swimtime="00:01:42.61" resultid="2355" heatid="3444" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1118" points="117" swimtime="00:01:50.37" resultid="2356" heatid="3461" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Malucelli" birthdate="2014-06-06" gender="M" nation="BRA" license="392153" swrid="5616448" athleteid="2501" externalid="392153">
              <RESULTS>
                <RESULT eventid="1083" status="DNS" swimtime="00:00:00.00" resultid="2502" heatid="3422" lane="6" entrytime="00:01:13.34" entrycourse="SCM" />
                <RESULT eventid="1071" status="DNS" swimtime="00:00:00.00" resultid="2503" heatid="3403" lane="6" entrytime="00:01:24.83" entrycourse="SCM" />
                <RESULT eventid="1131" status="DNS" swimtime="00:00:00.00" resultid="2504" heatid="3472" lane="7" entrytime="00:01:05.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Liam" lastname="Batista Grise" birthdate="2014-03-27" gender="M" nation="BRA" license="391008" swrid="5602514" athleteid="2428" externalid="391008">
              <RESULTS>
                <RESULT eventid="1095" status="DNS" swimtime="00:00:00.00" resultid="2429" heatid="3441" lane="5" entrytime="00:01:53.82" entrycourse="SCM" />
                <RESULT eventid="1071" status="DNS" swimtime="00:00:00.00" resultid="2430" heatid="3404" lane="8" entrytime="00:01:01.90" entrycourse="SCM" />
                <RESULT eventid="1131" status="DNS" swimtime="00:00:00.00" resultid="2431" heatid="3474" lane="7" entrytime="00:00:42.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicole" lastname="Rosario Osternack" birthdate="2008-04-11" gender="F" nation="BRA" license="331584" swrid="5600248" athleteid="1732" externalid="331584">
              <RESULTS>
                <RESULT eventid="1192" points="470" reactiontime="+72" swimtime="00:01:10.55" resultid="1733" heatid="3527" lane="6" entrytime="00:01:09.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="509" swimtime="00:00:30.53" resultid="1734" heatid="3515" lane="5" />
                <RESULT eventid="1288" points="492" swimtime="00:01:08.45" resultid="1735" heatid="3596" lane="7" entrytime="00:01:14.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="491" swimtime="00:00:31.99" resultid="1736" heatid="3587" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Clara Fernandes Pereira" birthdate="2009-11-19" gender="F" nation="BRA" license="344340" swrid="5600137" athleteid="1729" externalid="344340">
              <RESULTS>
                <RESULT eventid="1144" points="560" swimtime="00:04:40.53" resultid="1730" heatid="3494" lane="7" entrytime="00:04:47.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                    <SPLIT distance="100" swimtime="00:01:06.20" />
                    <SPLIT distance="150" swimtime="00:01:41.29" />
                    <SPLIT distance="200" swimtime="00:02:16.77" />
                    <SPLIT distance="250" swimtime="00:02:52.64" />
                    <SPLIT distance="300" swimtime="00:03:28.69" />
                    <SPLIT distance="350" swimtime="00:04:04.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="430" swimtime="00:02:41.44" resultid="1731" heatid="3556" lane="2" entrytime="00:02:42.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="100" swimtime="00:01:16.06" />
                    <SPLIT distance="150" swimtime="00:02:05.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="De Fortes" birthdate="2015-06-01" gender="M" nation="BRA" license="399680" swrid="5652884" athleteid="2565" externalid="399680">
              <RESULTS>
                <RESULT eventid="1095" points="62" swimtime="00:01:53.21" resultid="2566" heatid="3441" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="59" reactiontime="+80" swimtime="00:00:56.53" resultid="2567" heatid="3420" lane="2" />
                <RESULT eventid="1111" points="53" swimtime="00:00:57.78" resultid="2568" heatid="3457" lane="7" />
                <RESULT eventid="1131" points="69" swimtime="00:00:49.13" resultid="2569" heatid="3471" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Martinez Diniz" birthdate="2008-11-22" gender="M" nation="BRA" license="339400" athleteid="2694" externalid="339400">
              <RESULTS>
                <RESULT eventid="1168" points="334" swimtime="00:01:19.67" resultid="2695" heatid="3509" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="431" swimtime="00:04:40.87" resultid="2696" heatid="3496" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.79" />
                    <SPLIT distance="100" swimtime="00:01:05.49" />
                    <SPLIT distance="150" swimtime="00:01:41.71" />
                    <SPLIT distance="200" swimtime="00:02:18.26" />
                    <SPLIT distance="250" swimtime="00:02:54.52" />
                    <SPLIT distance="300" swimtime="00:03:30.66" />
                    <SPLIT distance="350" swimtime="00:04:06.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="434" swimtime="00:00:26.62" resultid="2697" heatid="3541" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Saber" birthdate="2014-06-04" gender="F" nation="BRA" license="392141" swrid="5602554" athleteid="2496" externalid="392141">
              <RESULTS>
                <RESULT eventid="1092" points="126" swimtime="00:01:40.04" resultid="2497" heatid="3437" lane="3" entrytime="00:01:59.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="155" swimtime="00:00:52.71" resultid="2498" heatid="3401" lane="3" entrytime="00:00:55.14" entrycourse="SCM" />
                <RESULT eventid="1108" points="81" swimtime="00:00:56.24" resultid="2499" heatid="3453" lane="1" />
                <RESULT eventid="1128" points="126" swimtime="00:00:45.63" resultid="2500" heatid="3468" lane="3" entrytime="00:00:46.52" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thais" lastname="Mariany Bortolazzi" birthdate="2006-05-02" gender="F" nation="BRA" license="357048" swrid="5600210" athleteid="2199" externalid="357048">
              <RESULTS>
                <RESULT eventid="1256" points="620" swimtime="00:17:44.82" resultid="2200" heatid="3582" lane="4" entrytime="00:18:22.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                    <SPLIT distance="100" swimtime="00:01:06.16" />
                    <SPLIT distance="150" swimtime="00:01:41.16" />
                    <SPLIT distance="200" swimtime="00:02:16.78" />
                    <SPLIT distance="250" swimtime="00:02:52.43" />
                    <SPLIT distance="300" swimtime="00:03:28.08" />
                    <SPLIT distance="350" swimtime="00:04:03.71" />
                    <SPLIT distance="400" swimtime="00:04:39.27" />
                    <SPLIT distance="450" swimtime="00:05:14.95" />
                    <SPLIT distance="500" swimtime="00:05:50.54" />
                    <SPLIT distance="550" swimtime="00:06:26.30" />
                    <SPLIT distance="600" swimtime="00:07:01.99" />
                    <SPLIT distance="650" swimtime="00:07:37.69" />
                    <SPLIT distance="700" swimtime="00:08:13.39" />
                    <SPLIT distance="750" swimtime="00:08:49.13" />
                    <SPLIT distance="800" swimtime="00:09:25.03" />
                    <SPLIT distance="850" swimtime="00:10:00.90" />
                    <SPLIT distance="900" swimtime="00:10:36.65" />
                    <SPLIT distance="950" swimtime="00:11:12.38" />
                    <SPLIT distance="1000" swimtime="00:11:48.00" />
                    <SPLIT distance="1050" swimtime="00:12:23.68" />
                    <SPLIT distance="1100" swimtime="00:12:59.50" />
                    <SPLIT distance="1150" swimtime="00:13:35.14" />
                    <SPLIT distance="1200" swimtime="00:14:11.01" />
                    <SPLIT distance="1250" swimtime="00:14:46.81" />
                    <SPLIT distance="1300" swimtime="00:15:22.52" />
                    <SPLIT distance="1350" swimtime="00:15:58.38" />
                    <SPLIT distance="1400" swimtime="00:16:34.50" />
                    <SPLIT distance="1450" swimtime="00:17:10.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Fontolan Gomes" birthdate="2010-07-02" gender="M" nation="BRA" license="356245" swrid="5588705" athleteid="1875" externalid="356245">
              <RESULTS>
                <RESULT eventid="1200" points="316" reactiontime="+75" swimtime="00:01:10.92" resultid="1876" heatid="3530" lane="4" entrytime="00:01:18.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="216" swimtime="00:01:32.03" resultid="1877" heatid="3509" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="262" reactiontime="+54" swimtime="00:00:34.55" resultid="1878" heatid="3591" lane="1" />
                <RESULT eventid="1264" points="344" swimtime="00:20:07.76" resultid="1879" heatid="3585" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:11.92" />
                    <SPLIT distance="150" swimtime="00:01:50.53" />
                    <SPLIT distance="200" swimtime="00:02:29.51" />
                    <SPLIT distance="250" swimtime="00:03:08.71" />
                    <SPLIT distance="300" swimtime="00:03:48.43" />
                    <SPLIT distance="350" swimtime="00:04:28.63" />
                    <SPLIT distance="400" swimtime="00:05:08.38" />
                    <SPLIT distance="450" swimtime="00:05:48.73" />
                    <SPLIT distance="500" swimtime="00:06:29.35" />
                    <SPLIT distance="550" swimtime="00:07:09.83" />
                    <SPLIT distance="600" swimtime="00:07:50.53" />
                    <SPLIT distance="650" swimtime="00:08:31.12" />
                    <SPLIT distance="700" swimtime="00:09:12.12" />
                    <SPLIT distance="750" swimtime="00:09:53.13" />
                    <SPLIT distance="800" swimtime="00:10:34.06" />
                    <SPLIT distance="850" swimtime="00:11:14.81" />
                    <SPLIT distance="900" swimtime="00:11:56.05" />
                    <SPLIT distance="950" swimtime="00:12:37.57" />
                    <SPLIT distance="1000" swimtime="00:13:18.87" />
                    <SPLIT distance="1050" swimtime="00:14:00.08" />
                    <SPLIT distance="1100" swimtime="00:14:40.97" />
                    <SPLIT distance="1150" swimtime="00:15:22.19" />
                    <SPLIT distance="1200" swimtime="00:16:03.55" />
                    <SPLIT distance="1250" swimtime="00:16:45.01" />
                    <SPLIT distance="1300" swimtime="00:17:27.01" />
                    <SPLIT distance="1350" swimtime="00:18:07.98" />
                    <SPLIT distance="1400" swimtime="00:18:48.82" />
                    <SPLIT distance="1450" swimtime="00:19:29.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="313" swimtime="00:01:06.02" resultid="1880" heatid="3576" lane="4" entrytime="00:01:10.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Felipe Canalli" birthdate="2015-12-23" gender="M" nation="BRA" license="406749" athleteid="2675" externalid="406749">
              <RESULTS>
                <RESULT eventid="1095" points="34" swimtime="00:02:17.16" resultid="2676" heatid="3440" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="91" swimtime="00:00:55.35" resultid="2677" heatid="3403" lane="7" />
                <RESULT eventid="1111" points="33" swimtime="00:01:07.59" resultid="2678" heatid="3456" lane="3" />
                <RESULT eventid="1131" points="40" swimtime="00:00:58.75" resultid="2679" heatid="3471" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Bussmann" birthdate="2007-01-16" gender="F" nation="BRA" license="313781" swrid="5579983" athleteid="1765" externalid="313781">
              <RESULTS>
                <RESULT eventid="1160" points="599" swimtime="00:01:13.97" resultid="1766" heatid="3506" lane="5" entrytime="00:01:16.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="499" swimtime="00:02:33.56" resultid="1767" heatid="3553" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                    <SPLIT distance="100" swimtime="00:01:16.33" />
                    <SPLIT distance="150" swimtime="00:01:57.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="481" swimtime="00:01:04.09" resultid="1768" heatid="3562" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Della Villa Yang" birthdate="2015-02-27" gender="F" nation="BRA" license="393283" swrid="5616442" athleteid="2535" externalid="393283">
              <RESULTS>
                <RESULT eventid="1092" points="121" swimtime="00:01:41.59" resultid="2536" heatid="3436" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="91" swimtime="00:01:02.88" resultid="2537" heatid="3400" lane="3" entrytime="00:01:13.68" entrycourse="SCM" />
                <RESULT eventid="1108" points="85" swimtime="00:00:55.39" resultid="2538" heatid="3455" lane="1" entrytime="00:01:00.02" entrycourse="SCM" />
                <RESULT eventid="1128" points="124" swimtime="00:00:45.90" resultid="2539" heatid="3467" lane="3" entrytime="00:00:58.91" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Gomes Santos" birthdate="2006-05-09" gender="M" nation="BRA" license="342833" athleteid="2630" externalid="342833">
              <RESULTS>
                <RESULT eventid="1152" points="642" swimtime="00:04:06.03" resultid="2631" heatid="3496" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                    <SPLIT distance="100" swimtime="00:00:59.81" />
                    <SPLIT distance="150" swimtime="00:01:30.89" />
                    <SPLIT distance="200" swimtime="00:02:02.14" />
                    <SPLIT distance="250" swimtime="00:02:33.21" />
                    <SPLIT distance="300" swimtime="00:03:04.39" />
                    <SPLIT distance="350" swimtime="00:03:35.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="658" swimtime="00:16:13.35" resultid="2632" heatid="3583" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.49" />
                    <SPLIT distance="100" swimtime="00:01:02.61" />
                    <SPLIT distance="150" swimtime="00:01:35.53" />
                    <SPLIT distance="200" swimtime="00:02:07.73" />
                    <SPLIT distance="250" swimtime="00:02:40.36" />
                    <SPLIT distance="300" swimtime="00:03:12.80" />
                    <SPLIT distance="350" swimtime="00:03:45.59" />
                    <SPLIT distance="400" swimtime="00:04:18.25" />
                    <SPLIT distance="450" swimtime="00:04:50.93" />
                    <SPLIT distance="500" swimtime="00:05:23.62" />
                    <SPLIT distance="550" swimtime="00:05:56.06" />
                    <SPLIT distance="600" swimtime="00:06:28.79" />
                    <SPLIT distance="650" swimtime="00:07:01.47" />
                    <SPLIT distance="700" swimtime="00:07:34.06" />
                    <SPLIT distance="750" swimtime="00:08:06.71" />
                    <SPLIT distance="800" swimtime="00:08:39.31" />
                    <SPLIT distance="850" swimtime="00:09:11.96" />
                    <SPLIT distance="900" swimtime="00:09:44.30" />
                    <SPLIT distance="950" swimtime="00:10:17.05" />
                    <SPLIT distance="1000" swimtime="00:10:49.58" />
                    <SPLIT distance="1050" swimtime="00:11:22.39" />
                    <SPLIT distance="1100" swimtime="00:11:55.00" />
                    <SPLIT distance="1150" swimtime="00:12:27.60" />
                    <SPLIT distance="1200" swimtime="00:13:00.27" />
                    <SPLIT distance="1250" swimtime="00:13:32.75" />
                    <SPLIT distance="1300" swimtime="00:14:05.23" />
                    <SPLIT distance="1350" swimtime="00:14:37.84" />
                    <SPLIT distance="1400" swimtime="00:15:10.00" />
                    <SPLIT distance="1450" swimtime="00:15:42.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Francia Soares" birthdate="2014-06-01" gender="F" nation="BRA" license="391011" swrid="5602540" athleteid="2432" externalid="391011">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="2433" heatid="3438" lane="8" entrytime="00:01:54.37" entrycourse="SCM" />
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="2434" heatid="3418" lane="3" entrytime="00:01:10.31" entrycourse="SCM" />
                <RESULT eventid="1128" points="73" swimtime="00:00:54.66" resultid="2435" heatid="3467" lane="5" entrytime="00:00:55.84" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Jacob Brunetti" birthdate="2015-11-10" gender="M" nation="BRA" license="406837" athleteid="2703" externalid="406837">
              <RESULTS>
                <RESULT eventid="1095" status="DSQ" swimtime="00:02:52.15" resultid="2704" heatid="3439" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:51.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="22" swimtime="00:01:18.03" resultid="2705" heatid="3422" lane="1" />
                <RESULT eventid="1111" points="12" swimtime="00:01:34.76" resultid="2706" heatid="3456" lane="2" />
                <RESULT eventid="1131" points="21" swimtime="00:01:12.39" resultid="2707" heatid="3471" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Shwetz Clivatti" birthdate="2015-03-05" gender="M" nation="BRA" license="406963" athleteid="2728" externalid="406963">
              <RESULTS>
                <RESULT eventid="1083" points="23" swimtime="00:01:17.17" resultid="2729" heatid="3420" lane="3" />
                <RESULT eventid="1071" points="31" swimtime="00:01:18.59" resultid="2730" heatid="3402" lane="5" />
                <RESULT eventid="1131" points="28" swimtime="00:01:06.35" resultid="2731" heatid="3470" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Sabedotti" birthdate="2002-07-07" gender="M" nation="BRA" license="134704" swrid="5600252" athleteid="1865" externalid="134704" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1168" points="694" swimtime="00:01:02.41" resultid="1866" heatid="3513" lane="5" entrytime="00:01:03.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="681" swimtime="00:02:04.56" resultid="1867" heatid="3561" lane="4" entrytime="00:02:03.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.14" />
                    <SPLIT distance="100" swimtime="00:01:00.18" />
                    <SPLIT distance="150" swimtime="00:01:35.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="644" swimtime="00:00:28.89" resultid="1868" heatid="3612" lane="4" entrytime="00:00:28.35" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Vanzo Assumpcao" birthdate="2012-05-15" gender="M" nation="BRA" license="369258" swrid="5588942" athleteid="2060" externalid="369258">
              <RESULTS>
                <RESULT eventid="1089" points="259" swimtime="00:02:35.73" resultid="2061" heatid="3430" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:15.27" />
                    <SPLIT distance="150" swimtime="00:01:55.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="217" reactiontime="+71" swimtime="00:00:36.77" resultid="2062" heatid="3415" lane="5" entrytime="00:00:37.46" entrycourse="SCM" />
                <RESULT eventid="1121" points="192" swimtime="00:01:22.70" resultid="2063" heatid="3464" lane="4" entrytime="00:01:25.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="228" swimtime="00:00:32.99" resultid="2064" heatid="3488" lane="3" entrytime="00:00:31.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Fontes Bonardi" birthdate="2008-10-26" gender="M" nation="BRA" license="307662" swrid="5600164" athleteid="1750" externalid="307662">
              <RESULTS>
                <RESULT eventid="1200" points="400" reactiontime="+71" swimtime="00:01:05.56" resultid="1751" heatid="3529" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="477" swimtime="00:01:10.74" resultid="1752" heatid="3509" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="408" swimtime="00:01:04.40" resultid="1753" heatid="3600" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Fernandes  Dos Reis" birthdate="2012-09-18" gender="M" nation="BRA" license="369279" swrid="5588696" athleteid="2135" externalid="369279">
              <RESULTS>
                <RESULT eventid="1089" points="256" swimtime="00:02:36.47" resultid="2136" heatid="3434" lane="1" entrytime="00:02:45.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:12.26" />
                    <SPLIT distance="150" swimtime="00:01:53.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="170" reactiontime="+107" swimtime="00:00:39.91" resultid="2137" heatid="3411" lane="5" />
                <RESULT eventid="1121" points="204" swimtime="00:01:21.12" resultid="2138" heatid="3464" lane="5" entrytime="00:01:27.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="247" swimtime="00:00:32.13" resultid="2139" heatid="3483" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Fontolan Gomes" birthdate="2008-05-01" gender="M" nation="BRA" license="307667" swrid="5600166" athleteid="1811" externalid="307667">
              <RESULTS>
                <RESULT eventid="1200" points="368" reactiontime="+76" swimtime="00:01:07.41" resultid="1812" heatid="3531" lane="5" entrytime="00:01:09.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="400" swimtime="00:02:28.76" resultid="1813" heatid="3560" lane="6" entrytime="00:02:34.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:10.34" />
                    <SPLIT distance="150" swimtime="00:01:53.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="334" reactiontime="+63" swimtime="00:00:31.85" resultid="1814" heatid="3590" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Valduga Artigas" birthdate="2009-06-01" gender="M" nation="BRA" license="339569" swrid="5600268" athleteid="1855" externalid="339569">
              <RESULTS>
                <RESULT eventid="1184" points="299" swimtime="00:00:32.51" resultid="1856" heatid="3518" lane="3" />
                <RESULT eventid="1296" points="280" swimtime="00:01:12.95" resultid="1857" heatid="3600" lane="4" entrytime="00:01:16.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Dolberth Alcantara" birthdate="2014-09-26" gender="F" nation="BRA" license="382124" swrid="5602532" athleteid="2373" externalid="382124">
              <RESULTS>
                <RESULT eventid="1080" points="99" reactiontime="+107" swimtime="00:00:54.49" resultid="2374" heatid="3418" lane="5" entrytime="00:00:57.59" entrycourse="SCM" />
                <RESULT eventid="1068" points="106" swimtime="00:00:59.93" resultid="2375" heatid="3401" lane="8" entrytime="00:01:04.51" entrycourse="SCM" />
                <RESULT eventid="1108" points="79" swimtime="00:00:56.61" resultid="2376" heatid="3455" lane="6" entrytime="00:00:59.20" entrycourse="SCM" />
                <RESULT eventid="1128" points="125" swimtime="00:00:45.78" resultid="2377" heatid="3468" lane="5" entrytime="00:00:46.25" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Marie Silva" birthdate="2014-08-24" gender="F" nation="BRA" license="391025" swrid="5602556" athleteid="2471" externalid="391025">
              <RESULTS>
                <RESULT eventid="1092" points="140" swimtime="00:01:36.62" resultid="2472" heatid="3438" lane="2" entrytime="00:01:43.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="120" swimtime="00:00:57.39" resultid="2473" heatid="3401" lane="2" entrytime="00:01:00.79" entrycourse="SCM" />
                <RESULT eventid="1108" points="95" swimtime="00:00:53.26" resultid="2474" heatid="3453" lane="6" />
                <RESULT eventid="1128" points="166" swimtime="00:00:41.68" resultid="2475" heatid="3468" lane="2" entrytime="00:00:49.60" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo" lastname="De Lima Cavalcanti" birthdate="2009-12-17" gender="M" nation="BRA" license="380965" swrid="5634589" athleteid="2618" externalid="380965">
              <RESULTS>
                <RESULT eventid="1184" points="439" swimtime="00:00:28.60" resultid="2619" heatid="3522" lane="2" entrytime="00:00:29.20" entrycourse="SCM" />
                <RESULT eventid="1216" points="458" swimtime="00:00:26.14" resultid="2620" heatid="3549" lane="4" entrytime="00:00:25.95" entrycourse="SCM" />
                <RESULT eventid="1296" points="448" swimtime="00:01:02.44" resultid="2621" heatid="3602" lane="6" entrytime="00:01:01.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Da Cunha Souza" birthdate="2013-09-17" gender="M" nation="BRA" license="376975" swrid="5588618" athleteid="2253" externalid="376975">
              <RESULTS>
                <RESULT eventid="1089" points="130" swimtime="00:03:16.14" resultid="2254" heatid="3431" lane="4" entrytime="00:03:13.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.37" />
                    <SPLIT distance="100" swimtime="00:01:34.90" />
                    <SPLIT distance="150" swimtime="00:02:28.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="89" swimtime="00:02:03.47" resultid="2255" heatid="3397" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="70" swimtime="00:01:55.56" resultid="2256" heatid="3463" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="143" swimtime="00:00:38.55" resultid="2257" heatid="3485" lane="2" entrytime="00:00:38.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Gustavo Souza" birthdate="2011-08-24" gender="M" nation="BRA" license="366901" swrid="5588733" athleteid="1998" externalid="366901">
              <RESULTS>
                <RESULT eventid="1200" points="195" reactiontime="+86" swimtime="00:01:23.31" resultid="1999" heatid="3529" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="333" swimtime="00:05:05.93" resultid="2000" heatid="3499" lane="1" entrytime="00:05:30.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:01:16.01" />
                    <SPLIT distance="150" swimtime="00:01:55.15" />
                    <SPLIT distance="200" swimtime="00:02:34.33" />
                    <SPLIT distance="250" swimtime="00:03:12.79" />
                    <SPLIT distance="300" swimtime="00:03:52.15" />
                    <SPLIT distance="350" swimtime="00:04:30.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="245" swimtime="00:02:55.12" resultid="2001" heatid="3559" lane="1" entrytime="00:03:03.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                    <SPLIT distance="100" swimtime="00:01:23.88" />
                    <SPLIT distance="150" swimtime="00:02:18.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="231" swimtime="00:01:17.82" resultid="2002" heatid="3600" lane="6" entrytime="00:01:23.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="312" swimtime="00:20:47.55" resultid="2003" heatid="3584" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.23" />
                    <SPLIT distance="100" swimtime="00:01:21.65" />
                    <SPLIT distance="150" swimtime="00:02:03.61" />
                    <SPLIT distance="200" swimtime="00:02:45.68" />
                    <SPLIT distance="250" swimtime="00:03:27.92" />
                    <SPLIT distance="300" swimtime="00:04:10.61" />
                    <SPLIT distance="350" swimtime="00:04:52.82" />
                    <SPLIT distance="400" swimtime="00:05:34.84" />
                    <SPLIT distance="450" swimtime="00:06:17.54" />
                    <SPLIT distance="500" swimtime="00:07:00.19" />
                    <SPLIT distance="550" swimtime="00:07:42.94" />
                    <SPLIT distance="600" swimtime="00:08:25.31" />
                    <SPLIT distance="650" swimtime="00:09:07.33" />
                    <SPLIT distance="700" swimtime="00:09:50.38" />
                    <SPLIT distance="750" swimtime="00:10:32.59" />
                    <SPLIT distance="800" swimtime="00:11:14.21" />
                    <SPLIT distance="850" swimtime="00:11:56.39" />
                    <SPLIT distance="900" swimtime="00:12:38.40" />
                    <SPLIT distance="950" swimtime="00:13:20.38" />
                    <SPLIT distance="1000" swimtime="00:14:02.04" />
                    <SPLIT distance="1050" swimtime="00:14:43.83" />
                    <SPLIT distance="1100" swimtime="00:15:26.35" />
                    <SPLIT distance="1150" swimtime="00:16:07.91" />
                    <SPLIT distance="1200" swimtime="00:16:49.92" />
                    <SPLIT distance="1250" swimtime="00:17:30.93" />
                    <SPLIT distance="1300" swimtime="00:18:12.67" />
                    <SPLIT distance="1350" swimtime="00:18:51.59" />
                    <SPLIT distance="1400" swimtime="00:19:32.27" />
                    <SPLIT distance="1450" swimtime="00:20:11.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Portes Fabiane" birthdate="2012-12-28" gender="M" nation="BRA" license="376983" swrid="5588864" athleteid="2286" externalid="376983">
              <RESULTS>
                <RESULT eventid="1077" points="58" reactiontime="+79" swimtime="00:00:56.83" resultid="2287" heatid="3413" lane="2" entrytime="00:00:57.49" entrycourse="SCM" />
                <RESULT eventid="1065" points="85" swimtime="00:02:05.42" resultid="2288" heatid="3397" lane="5" entrytime="00:02:08.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="71" swimtime="00:01:58.66" resultid="2289" heatid="3449" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="79" swimtime="00:00:46.80" resultid="2290" heatid="3483" lane="6" entrytime="00:00:47.44" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Cury Abreu" birthdate="2013-05-17" gender="F" nation="BRA" license="376974" swrid="5588614" athleteid="2248" externalid="376974">
              <RESULTS>
                <RESULT eventid="1086" points="261" swimtime="00:02:52.45" resultid="2249" heatid="3426" lane="1" entrytime="00:03:31.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.06" />
                    <SPLIT distance="100" swimtime="00:01:24.18" />
                    <SPLIT distance="150" swimtime="00:02:11.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="249" reactiontime="+76" swimtime="00:00:40.12" resultid="2250" heatid="3407" lane="5" />
                <RESULT eventid="1102" status="DSQ" swimtime="00:01:33.38" resultid="2251" heatid="3447" lane="1" entrytime="00:01:47.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="303" swimtime="00:00:34.13" resultid="2252" heatid="3480" lane="1" entrytime="00:00:38.82" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietra" lastname="Ruschel Carvalho" birthdate="2009-03-21" gender="F" nation="BRA" license="324999" swrid="5600250" athleteid="1737" externalid="324999">
              <RESULTS>
                <RESULT eventid="1208" points="566" swimtime="00:00:27.71" resultid="1738" heatid="3539" lane="5" entrytime="00:00:28.19" entrycourse="SCM" />
                <RESULT eventid="1176" points="483" swimtime="00:00:31.07" resultid="1739" heatid="3516" lane="4" entrytime="00:00:32.32" entrycourse="SCM" />
                <RESULT eventid="1272" points="389" reactiontime="+57" swimtime="00:00:34.56" resultid="1740" heatid="3587" lane="1" />
                <RESULT eventid="1240" points="561" swimtime="00:01:00.92" resultid="1741" heatid="3570" lane="3" entrytime="00:01:01.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcela" lastname="Tallao Benke" birthdate="2014-10-07" gender="F" nation="BRA" license="382075" swrid="5602586" athleteid="2368" externalid="382075">
              <RESULTS>
                <RESULT eventid="1092" points="219" swimtime="00:01:23.36" resultid="2369" heatid="3438" lane="5" entrytime="00:01:26.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="208" swimtime="00:00:47.82" resultid="2370" heatid="3401" lane="5" entrytime="00:00:52.47" entrycourse="SCM" />
                <RESULT eventid="1108" points="215" swimtime="00:00:40.65" resultid="2371" heatid="3455" lane="5" entrytime="00:00:49.63" entrycourse="SCM" />
                <RESULT eventid="1128" points="239" swimtime="00:00:36.93" resultid="2372" heatid="3469" lane="5" entrytime="00:00:39.82" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Hadad" birthdate="2015-09-09" gender="M" nation="BRA" license="406740" athleteid="2633" externalid="406740">
              <RESULTS>
                <RESULT eventid="1083" points="30" swimtime="00:01:11.14" resultid="2634" heatid="3420" lane="4" />
                <RESULT eventid="1071" status="DSQ" swimtime="00:01:08.89" resultid="2635" heatid="3403" lane="2" />
                <RESULT eventid="1111" status="DSQ" swimtime="00:01:15.10" resultid="2636" heatid="3457" lane="1" />
                <RESULT eventid="1131" points="31" swimtime="00:01:03.84" resultid="2637" heatid="3471" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Azevedo Alanis" birthdate="2013-12-07" gender="M" nation="BRA" license="376991" swrid="5588540" athleteid="2317" externalid="376991">
              <RESULTS>
                <RESULT eventid="1089" points="102" swimtime="00:03:32.18" resultid="2318" heatid="3431" lane="7" entrytime="00:03:31.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.99" />
                    <SPLIT distance="100" swimtime="00:01:43.24" />
                    <SPLIT distance="150" swimtime="00:02:38.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="104" swimtime="00:01:57.27" resultid="2319" heatid="3395" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="101" swimtime="00:01:45.48" resultid="2320" heatid="3450" lane="4" entrytime="00:01:47.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="109" swimtime="00:00:42.16" resultid="2321" heatid="3484" lane="2" entrytime="00:00:42.46" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Henrique Tiboni Araujo" birthdate="2013-06-11" gender="M" nation="BRA" license="376968" swrid="5588747" athleteid="2230" externalid="376968">
              <RESULTS>
                <RESULT eventid="1089" points="121" swimtime="00:03:20.39" resultid="2231" heatid="3431" lane="6" entrytime="00:03:29.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.67" />
                    <SPLIT distance="100" swimtime="00:01:36.22" />
                    <SPLIT distance="150" swimtime="00:02:28.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="96" reactiontime="+55" swimtime="00:00:48.20" resultid="2232" heatid="3414" lane="7" entrytime="00:00:47.00" entrycourse="SCM" />
                <RESULT eventid="1105" points="103" swimtime="00:01:44.88" resultid="2233" heatid="3450" lane="5" entrytime="00:01:51.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="149" swimtime="00:00:37.98" resultid="2234" heatid="3484" lane="3" entrytime="00:00:39.63" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Luiz Garcia Franceschi" birthdate="2013-01-12" gender="M" nation="BRA" license="376979" swrid="5588781" athleteid="2268" externalid="376979">
              <RESULTS>
                <RESULT eventid="1089" points="93" swimtime="00:03:38.91" resultid="2269" heatid="3430" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.95" />
                    <SPLIT distance="100" swimtime="00:01:44.45" />
                    <SPLIT distance="150" swimtime="00:02:43.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="99" swimtime="00:01:59.17" resultid="2270" heatid="3396" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Mattioli" birthdate="2011-10-22" gender="F" nation="BRA" license="366896" swrid="5602559" athleteid="1980" externalid="366896">
              <RESULTS>
                <RESULT eventid="1144" points="409" swimtime="00:05:11.52" resultid="1981" heatid="3493" lane="6" entrytime="00:05:23.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:14.35" />
                    <SPLIT distance="150" swimtime="00:01:54.13" />
                    <SPLIT distance="200" swimtime="00:02:33.63" />
                    <SPLIT distance="250" swimtime="00:03:14.19" />
                    <SPLIT distance="300" swimtime="00:03:55.04" />
                    <SPLIT distance="350" swimtime="00:04:35.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="295" reactiontime="+92" swimtime="00:01:22.39" resultid="1982" heatid="3525" lane="6" entrytime="00:01:24.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="319" swimtime="00:01:31.22" resultid="1983" heatid="3505" lane="1" entrytime="00:01:31.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="361" swimtime="00:02:51.01" resultid="1984" heatid="3555" lane="8" entrytime="00:02:57.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                    <SPLIT distance="100" swimtime="00:01:23.31" />
                    <SPLIT distance="150" swimtime="00:02:13.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="382" swimtime="00:01:09.25" resultid="1985" heatid="3563" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Cabrera Cirino Dos Santos" birthdate="2013-03-30" gender="M" nation="BRA" license="376990" swrid="5588570" athleteid="2322" externalid="376990">
              <RESULTS>
                <RESULT eventid="1089" points="184" swimtime="00:02:54.59" resultid="2323" heatid="3433" lane="1" entrytime="00:02:54.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                    <SPLIT distance="100" swimtime="00:01:23.92" />
                    <SPLIT distance="150" swimtime="00:02:10.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="121" reactiontime="+79" swimtime="00:00:44.67" resultid="2324" heatid="3414" lane="2" entrytime="00:00:43.92" entrycourse="SCM" />
                <RESULT eventid="1105" points="144" swimtime="00:01:33.92" resultid="2325" heatid="3449" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="203" swimtime="00:00:34.29" resultid="2326" heatid="3487" lane="2" entrytime="00:00:34.37" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Krupacz" birthdate="2008-04-18" gender="F" nation="BRA" license="329187" swrid="5634611" athleteid="2610" externalid="329187">
              <RESULTS>
                <RESULT eventid="1224" points="477" swimtime="00:02:35.88" resultid="2611" heatid="3551" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                    <SPLIT distance="100" swimtime="00:01:10.85" />
                    <SPLIT distance="150" swimtime="00:01:59.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="556" reactiontime="+67" swimtime="00:00:30.70" resultid="2612" heatid="3589" lane="5" entrytime="00:00:31.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Cunha Moraes" birthdate="2012-11-26" gender="F" nation="BRA" license="406744" athleteid="2653" externalid="406744">
              <RESULTS>
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="2654" heatid="3406" lane="5" />
                <RESULT eventid="1138" status="DNS" swimtime="00:00:00.00" resultid="2655" heatid="3477" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Guimaraes E Souza" birthdate="2008-12-21" gender="M" nation="BRA" license="376972" swrid="5600182" athleteid="2245" externalid="376972">
              <RESULTS>
                <RESULT eventid="1168" points="440" swimtime="00:01:12.63" resultid="2246" heatid="3511" lane="3" entrytime="00:01:22.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="378" swimtime="00:02:31.56" resultid="2247" heatid="3560" lane="2" entrytime="00:02:39.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:15.04" />
                    <SPLIT distance="150" swimtime="00:01:59.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Clara Prado Biscaia" birthdate="2013-10-24" gender="F" nation="BRA" license="391015" swrid="5602526" athleteid="2436" externalid="391015">
              <RESULTS>
                <RESULT eventid="1086" points="161" swimtime="00:03:22.37" resultid="2437" heatid="3425" lane="4" entrytime="00:03:35.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.86" />
                    <SPLIT distance="100" swimtime="00:01:40.23" />
                    <SPLIT distance="150" swimtime="00:02:32.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="115" reactiontime="+94" swimtime="00:00:51.80" resultid="2438" heatid="3407" lane="7" />
                <RESULT eventid="1118" status="DSQ" swimtime="00:01:52.38" resultid="2439" heatid="3461" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="130" swimtime="00:00:45.18" resultid="2440" heatid="3479" lane="7" entrytime="00:00:43.21" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe Alves" lastname="Franca Silva" birthdate="1987-05-14" gender="M" nation="BRA" license="14360" swrid="4300572" athleteid="3615" externalid="14360">
              <RESULTS>
                <RESULT eventid="1168" points="685" swimtime="00:01:02.70" resultid="3616" heatid="3508" lane="8" late="yes">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" status="DNS" swimtime="00:00:00.00" resultid="3617" heatid="3607" lane="7" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fernandes" birthdate="2010-03-13" gender="M" nation="BRA" license="339266" swrid="5588695" athleteid="2407" externalid="339266">
              <RESULTS>
                <RESULT eventid="1200" points="389" swimtime="00:01:06.18" resultid="2408" heatid="3532" lane="8" entrytime="00:01:08.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="355" swimtime="00:01:18.02" resultid="2409" heatid="3509" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="444" swimtime="00:00:26.41" resultid="2410" heatid="3548" lane="4" entrytime="00:00:26.87" entrycourse="SCM" />
                <RESULT eventid="1232" points="385" swimtime="00:02:30.57" resultid="2411" heatid="3560" lane="5" entrytime="00:02:31.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                    <SPLIT distance="100" swimtime="00:01:11.02" />
                    <SPLIT distance="150" swimtime="00:01:57.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="457" swimtime="00:00:58.19" resultid="2412" heatid="3579" lane="2" entrytime="00:00:59.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="De Almeida Dias" birthdate="2012-02-18" gender="F" nation="BRA" license="369262" swrid="5588638" athleteid="2075" externalid="369262">
              <RESULTS>
                <RESULT eventid="1062" points="355" swimtime="00:01:28.05" resultid="2076" heatid="3394" lane="5" entrytime="00:01:35.59" entrycourse="SCM" />
                <RESULT eventid="1086" points="432" swimtime="00:02:25.83" resultid="2077" heatid="3428" lane="3" entrytime="00:02:38.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                    <SPLIT distance="100" swimtime="00:01:11.76" />
                    <SPLIT distance="150" swimtime="00:01:49.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="337" swimtime="00:01:21.17" resultid="2078" heatid="3444" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="373" swimtime="00:00:31.84" resultid="2079" heatid="3480" lane="4" entrytime="00:00:34.70" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolau" lastname="Neto" birthdate="2011-03-22" gender="M" nation="BRA" license="366906" swrid="5602565" athleteid="2016" externalid="366906">
              <RESULTS>
                <RESULT eventid="1168" points="306" swimtime="00:01:22.03" resultid="2017" heatid="3510" lane="3" entrytime="00:01:28.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="312" swimtime="00:00:29.70" resultid="2018" heatid="3546" lane="1" entrytime="00:00:30.34" entrycourse="SCM" />
                <RESULT eventid="1232" points="289" swimtime="00:02:45.70" resultid="2019" heatid="3559" lane="3" entrytime="00:02:55.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.26" />
                    <SPLIT distance="100" swimtime="00:01:26.21" />
                    <SPLIT distance="150" swimtime="00:02:10.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="343" swimtime="00:20:08.73" resultid="2020" heatid="3585" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:14.09" />
                    <SPLIT distance="150" swimtime="00:01:53.21" />
                    <SPLIT distance="200" swimtime="00:02:33.79" />
                    <SPLIT distance="250" swimtime="00:03:14.21" />
                    <SPLIT distance="300" swimtime="00:03:54.83" />
                    <SPLIT distance="350" swimtime="00:04:36.24" />
                    <SPLIT distance="400" swimtime="00:05:17.58" />
                    <SPLIT distance="450" swimtime="00:05:59.47" />
                    <SPLIT distance="500" swimtime="00:06:40.77" />
                    <SPLIT distance="550" swimtime="00:07:21.67" />
                    <SPLIT distance="600" swimtime="00:08:03.09" />
                    <SPLIT distance="650" swimtime="00:08:43.60" />
                    <SPLIT distance="700" swimtime="00:09:24.75" />
                    <SPLIT distance="750" swimtime="00:10:05.09" />
                    <SPLIT distance="800" swimtime="00:10:45.73" />
                    <SPLIT distance="850" swimtime="00:11:26.49" />
                    <SPLIT distance="900" swimtime="00:12:07.20" />
                    <SPLIT distance="950" swimtime="00:12:47.91" />
                    <SPLIT distance="1000" swimtime="00:13:28.67" />
                    <SPLIT distance="1050" swimtime="00:14:09.69" />
                    <SPLIT distance="1100" swimtime="00:14:50.64" />
                    <SPLIT distance="1150" swimtime="00:15:30.77" />
                    <SPLIT distance="1200" swimtime="00:16:11.11" />
                    <SPLIT distance="1250" swimtime="00:16:51.45" />
                    <SPLIT distance="1300" swimtime="00:17:32.33" />
                    <SPLIT distance="1350" swimtime="00:18:12.36" />
                    <SPLIT distance="1400" swimtime="00:18:52.40" />
                    <SPLIT distance="1450" swimtime="00:19:31.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="334" swimtime="00:01:04.59" resultid="2021" heatid="3576" lane="6" entrytime="00:01:12.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Kirchgassner" birthdate="2007-02-10" gender="M" nation="BRA" license="313535" swrid="5600230" athleteid="1799" externalid="313535">
              <RESULTS>
                <RESULT eventid="1168" points="605" swimtime="00:01:05.34" resultid="1800" heatid="3513" lane="2" entrytime="00:01:07.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="519" swimtime="00:02:16.39" resultid="1801" heatid="3561" lane="2" entrytime="00:02:19.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                    <SPLIT distance="100" swimtime="00:01:06.22" />
                    <SPLIT distance="150" swimtime="00:01:44.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="516" swimtime="00:00:59.56" resultid="1802" heatid="3599" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Szpak Zraik" birthdate="2015-04-10" gender="M" nation="BRA" license="393259" swrid="5616451" athleteid="2505" externalid="393259">
              <RESULTS>
                <RESULT eventid="1095" points="78" swimtime="00:01:44.79" resultid="2506" heatid="3440" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="102" swimtime="00:00:53.33" resultid="2507" heatid="3404" lane="7" entrytime="00:01:01.53" entrycourse="SCM" />
                <RESULT eventid="1111" points="31" swimtime="00:01:08.60" resultid="2508" heatid="3458" lane="6" />
                <RESULT eventid="1131" points="86" swimtime="00:00:45.52" resultid="2509" heatid="3472" lane="3" entrytime="00:00:52.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Pisani Ferreira" birthdate="2012-08-06" gender="F" nation="BRA" license="376985" swrid="5588862" athleteid="2342" externalid="376985">
              <RESULTS>
                <RESULT eventid="1062" points="186" swimtime="00:01:49.17" resultid="2343" heatid="3394" lane="2" entrytime="00:01:55.91" entrycourse="SCM" />
                <RESULT eventid="1074" points="122" swimtime="00:00:50.91" resultid="2344" heatid="3407" lane="8" />
                <RESULT eventid="1102" points="157" swimtime="00:01:44.61" resultid="2345" heatid="3446" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="198" swimtime="00:00:39.34" resultid="2346" heatid="3479" lane="1" entrytime="00:00:43.27" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Germer Munhoz" birthdate="2010-04-23" gender="F" nation="BRA" license="356632" swrid="5588722" athleteid="1934" externalid="356632">
              <RESULTS>
                <RESULT eventid="1144" points="495" swimtime="00:04:52.21" resultid="1935" heatid="3493" lane="5" entrytime="00:05:18.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:08.85" />
                    <SPLIT distance="150" swimtime="00:01:45.39" />
                    <SPLIT distance="200" swimtime="00:02:22.37" />
                    <SPLIT distance="250" swimtime="00:03:00.40" />
                    <SPLIT distance="300" swimtime="00:03:38.30" />
                    <SPLIT distance="350" swimtime="00:04:16.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" status="DSQ" swimtime="00:01:28.97" resultid="1936" heatid="3502" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="433" swimtime="00:02:41.06" resultid="1937" heatid="3556" lane="8" entrytime="00:02:47.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:18.67" />
                    <SPLIT distance="150" swimtime="00:02:06.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="346" swimtime="00:01:16.96" resultid="1938" heatid="3596" lane="1" entrytime="00:01:16.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="405" swimtime="00:01:07.90" resultid="1939" heatid="3569" lane="7" entrytime="00:01:07.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Da Cunha Souza" birthdate="2015-05-30" gender="F" nation="BRA" license="400016" swrid="5652883" athleteid="2575" externalid="400016">
              <RESULTS>
                <RESULT eventid="1092" points="94" swimtime="00:01:50.51" resultid="2576" heatid="3437" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="92" swimtime="00:01:02.80" resultid="2577" heatid="3400" lane="7" />
                <RESULT eventid="1108" points="61" swimtime="00:01:01.86" resultid="2578" heatid="3453" lane="3" />
                <RESULT eventid="1128" points="103" swimtime="00:00:48.76" resultid="2579" heatid="3465" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Almeida Jorge" birthdate="2015-05-27" gender="M" nation="BRA" license="406836" athleteid="2698" externalid="406836">
              <RESULTS>
                <RESULT eventid="1095" points="26" swimtime="00:02:30.60" resultid="2699" heatid="3439" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="45" swimtime="00:01:09.86" resultid="2700" heatid="3402" lane="6" />
                <RESULT eventid="1111" points="22" swimtime="00:01:17.22" resultid="2701" heatid="3458" lane="8" />
                <RESULT eventid="1131" points="27" swimtime="00:01:07.06" resultid="2702" heatid="3470" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Coelho" birthdate="2011-11-11" gender="M" nation="BRA" license="366889" swrid="5602527" athleteid="1962" externalid="366889">
              <RESULTS>
                <RESULT eventid="1200" points="216" swimtime="00:01:20.48" resultid="1963" heatid="3530" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="379" swimtime="00:04:53.26" resultid="1964" heatid="3499" lane="4" entrytime="00:05:08.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="100" swimtime="00:01:10.89" />
                    <SPLIT distance="150" swimtime="00:01:48.40" />
                    <SPLIT distance="200" swimtime="00:02:25.68" />
                    <SPLIT distance="250" swimtime="00:03:03.48" />
                    <SPLIT distance="300" swimtime="00:03:40.92" />
                    <SPLIT distance="350" swimtime="00:04:17.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="240" swimtime="00:01:16.81" resultid="1965" heatid="3600" lane="3" entrytime="00:01:19.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="376" swimtime="00:19:33.22" resultid="1966" heatid="3584" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                    <SPLIT distance="100" swimtime="00:01:19.18" />
                    <SPLIT distance="150" swimtime="00:01:59.67" />
                    <SPLIT distance="200" swimtime="00:02:40.20" />
                    <SPLIT distance="250" swimtime="00:03:20.11" />
                    <SPLIT distance="300" swimtime="00:04:00.38" />
                    <SPLIT distance="350" swimtime="00:04:40.45" />
                    <SPLIT distance="400" swimtime="00:05:20.81" />
                    <SPLIT distance="450" swimtime="00:06:00.36" />
                    <SPLIT distance="500" swimtime="00:06:40.51" />
                    <SPLIT distance="550" swimtime="00:07:19.98" />
                    <SPLIT distance="600" swimtime="00:08:00.10" />
                    <SPLIT distance="650" swimtime="00:08:39.99" />
                    <SPLIT distance="700" swimtime="00:09:19.86" />
                    <SPLIT distance="750" swimtime="00:09:59.69" />
                    <SPLIT distance="800" swimtime="00:10:39.08" />
                    <SPLIT distance="850" swimtime="00:11:18.69" />
                    <SPLIT distance="900" swimtime="00:11:57.69" />
                    <SPLIT distance="950" swimtime="00:12:36.96" />
                    <SPLIT distance="1000" swimtime="00:13:16.08" />
                    <SPLIT distance="1050" swimtime="00:13:55.35" />
                    <SPLIT distance="1100" swimtime="00:14:34.15" />
                    <SPLIT distance="1150" swimtime="00:15:12.20" />
                    <SPLIT distance="1200" swimtime="00:15:50.61" />
                    <SPLIT distance="1250" swimtime="00:16:28.53" />
                    <SPLIT distance="1300" swimtime="00:17:06.53" />
                    <SPLIT distance="1350" swimtime="00:17:43.93" />
                    <SPLIT distance="1400" swimtime="00:18:21.94" />
                    <SPLIT distance="1450" swimtime="00:18:58.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="331" swimtime="00:01:04.81" resultid="1967" heatid="3577" lane="5" entrytime="00:01:06.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Pereira Galle" birthdate="2011-08-02" gender="F" nation="BRA" license="369465" swrid="5627330" athleteid="2600" externalid="369465">
              <RESULTS>
                <RESULT eventid="1144" points="379" swimtime="00:05:19.59" resultid="2601" heatid="3493" lane="1" entrytime="00:05:30.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="100" swimtime="00:01:13.42" />
                    <SPLIT distance="150" swimtime="00:01:52.97" />
                    <SPLIT distance="200" swimtime="00:02:33.84" />
                    <SPLIT distance="250" swimtime="00:03:15.15" />
                    <SPLIT distance="300" swimtime="00:03:57.29" />
                    <SPLIT distance="350" swimtime="00:04:38.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="375" swimtime="00:01:26.43" resultid="2602" heatid="3505" lane="3" entrytime="00:01:24.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="353" swimtime="00:02:52.37" resultid="2603" heatid="3554" lane="4" entrytime="00:02:59.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.48" />
                    <SPLIT distance="100" swimtime="00:01:23.50" />
                    <SPLIT distance="150" swimtime="00:02:14.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="266" swimtime="00:01:23.97" resultid="2604" heatid="3594" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="394" swimtime="00:01:08.49" resultid="2605" heatid="3563" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Viera Correa" birthdate="2012-03-07" gender="M" nation="BRA" license="369269" swrid="5602590" athleteid="2090" externalid="369269">
              <RESULTS>
                <RESULT eventid="1089" points="245" swimtime="00:02:38.73" resultid="2091" heatid="3434" lane="3" entrytime="00:02:40.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:16.16" />
                    <SPLIT distance="150" swimtime="00:01:58.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="189" reactiontime="+84" swimtime="00:00:38.50" resultid="2092" heatid="3415" lane="2" entrytime="00:00:39.54" entrycourse="SCM" />
                <RESULT eventid="1105" points="206" swimtime="00:01:23.33" resultid="2093" heatid="3448" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="253" swimtime="00:00:31.84" resultid="2094" heatid="3488" lane="1" entrytime="00:00:32.79" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Bittencourt Ribas" birthdate="2013-02-01" gender="F" nation="BRA" license="372682" swrid="5588555" athleteid="2166" externalid="372682">
              <RESULTS>
                <RESULT eventid="1086" points="292" swimtime="00:02:46.11" resultid="2167" heatid="3427" lane="5" entrytime="00:02:48.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                    <SPLIT distance="100" swimtime="00:01:22.12" />
                    <SPLIT distance="150" swimtime="00:02:06.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="223" swimtime="00:00:41.60" resultid="2168" heatid="3410" lane="8" entrytime="00:00:41.65" entrycourse="SCM" />
                <RESULT eventid="1102" points="252" swimtime="00:01:29.43" resultid="2169" heatid="3447" lane="3" entrytime="00:01:34.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1118" status="DSQ" swimtime="00:01:36.17" resultid="2170" heatid="3461" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Fontes Hoshina" birthdate="2008-02-15" gender="M" nation="BRA" license="369445" swrid="5600165" athleteid="1758" externalid="369445">
              <RESULTS>
                <RESULT eventid="1184" points="565" swimtime="00:00:26.30" resultid="1759" heatid="3517" lane="6" />
                <RESULT eventid="1296" points="544" swimtime="00:00:58.51" resultid="1760" heatid="3598" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="561" swimtime="00:00:54.34" resultid="1761" heatid="3574" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Guimaraes Mesquita" birthdate="2015-10-05" gender="F" nation="BRA" license="393263" swrid="5616444" athleteid="2525" externalid="393263">
              <RESULTS>
                <RESULT eventid="1092" points="33" swimtime="00:02:35.77" resultid="2526" heatid="3436" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="54" swimtime="00:01:06.79" resultid="2527" heatid="3416" lane="4" />
                <RESULT eventid="1108" points="16" swimtime="00:01:35.32" resultid="2528" heatid="3452" lane="6" />
                <RESULT eventid="1128" points="28" swimtime="00:01:15.20" resultid="2529" heatid="3467" lane="7" entrytime="00:01:23.08" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Schiavon" birthdate="2010-05-03" gender="M" nation="BRA" license="356354" swrid="5600256" athleteid="1916" externalid="356354">
              <RESULTS>
                <RESULT eventid="1200" points="247" reactiontime="+80" swimtime="00:01:16.94" resultid="1917" heatid="3528" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="450" swimtime="00:04:36.80" resultid="1918" heatid="3499" lane="5" entrytime="00:05:11.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                    <SPLIT distance="100" swimtime="00:01:05.03" />
                    <SPLIT distance="150" swimtime="00:01:39.52" />
                    <SPLIT distance="200" swimtime="00:02:15.02" />
                    <SPLIT distance="250" swimtime="00:02:50.24" />
                    <SPLIT distance="300" swimtime="00:03:26.06" />
                    <SPLIT distance="350" swimtime="00:04:02.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="280" swimtime="00:02:47.49" resultid="1919" heatid="3559" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.59" />
                    <SPLIT distance="100" swimtime="00:01:20.15" />
                    <SPLIT distance="150" swimtime="00:02:10.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="171" swimtime="00:01:26.07" resultid="1920" heatid="3599" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="453" swimtime="00:18:22.11" resultid="1921" heatid="3584" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                    <SPLIT distance="100" swimtime="00:01:06.31" />
                    <SPLIT distance="150" swimtime="00:01:42.06" />
                    <SPLIT distance="200" swimtime="00:02:18.15" />
                    <SPLIT distance="250" swimtime="00:02:54.15" />
                    <SPLIT distance="300" swimtime="00:03:30.42" />
                    <SPLIT distance="350" swimtime="00:04:06.98" />
                    <SPLIT distance="400" swimtime="00:04:43.65" />
                    <SPLIT distance="450" swimtime="00:05:20.84" />
                    <SPLIT distance="500" swimtime="00:05:57.99" />
                    <SPLIT distance="550" swimtime="00:06:35.12" />
                    <SPLIT distance="600" swimtime="00:07:11.97" />
                    <SPLIT distance="650" swimtime="00:07:49.19" />
                    <SPLIT distance="700" swimtime="00:08:26.23" />
                    <SPLIT distance="750" swimtime="00:09:03.00" />
                    <SPLIT distance="800" swimtime="00:09:40.21" />
                    <SPLIT distance="850" swimtime="00:10:17.83" />
                    <SPLIT distance="900" swimtime="00:10:54.66" />
                    <SPLIT distance="950" swimtime="00:11:31.99" />
                    <SPLIT distance="1000" swimtime="00:12:09.53" />
                    <SPLIT distance="1050" swimtime="00:12:46.80" />
                    <SPLIT distance="1100" swimtime="00:13:23.97" />
                    <SPLIT distance="1150" swimtime="00:14:01.05" />
                    <SPLIT distance="1200" swimtime="00:14:38.58" />
                    <SPLIT distance="1250" swimtime="00:15:15.98" />
                    <SPLIT distance="1300" swimtime="00:15:54.03" />
                    <SPLIT distance="1350" swimtime="00:16:31.88" />
                    <SPLIT distance="1400" swimtime="00:17:09.65" />
                    <SPLIT distance="1450" swimtime="00:17:46.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivia" lastname="Jeger" birthdate="2004-12-19" gender="F" nation="BRA" license="325493" swrid="5600193" athleteid="2589" externalid="325493" level="UNIDOMBOSC">
              <RESULTS>
                <RESULT eventid="1144" points="647" swimtime="00:04:27.36" resultid="2590" heatid="3494" lane="5" entrytime="00:04:27.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="100" swimtime="00:01:04.07" />
                    <SPLIT distance="150" swimtime="00:01:37.96" />
                    <SPLIT distance="200" swimtime="00:02:11.92" />
                    <SPLIT distance="250" swimtime="00:02:45.88" />
                    <SPLIT distance="300" swimtime="00:03:20.07" />
                    <SPLIT distance="350" swimtime="00:03:54.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" status="DNS" swimtime="00:00:00.00" resultid="2591" heatid="3502" lane="7" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="2592" heatid="3556" lane="4" entrytime="00:02:25.78" entrycourse="SCM" />
                <RESULT eventid="1288" points="527" swimtime="00:01:06.89" resultid="2593" heatid="3596" lane="5" entrytime="00:01:06.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helen" lastname="Barato Bernardi" birthdate="2006-07-27" gender="F" nation="BRA" license="317031" athleteid="2622" externalid="317031">
              <RESULTS>
                <RESULT eventid="1160" points="624" swimtime="00:01:12.94" resultid="2623" heatid="3506" lane="4" entrytime="00:01:11.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="460" swimtime="00:02:37.80" resultid="2624" heatid="3556" lane="6" entrytime="00:02:41.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                    <SPLIT distance="100" swimtime="00:01:19.21" />
                    <SPLIT distance="150" swimtime="00:02:01.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="623" swimtime="00:00:33.20" resultid="2625" heatid="3606" lane="4" entrytime="00:00:32.53" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alan" lastname="Batista Grise" birthdate="2014-03-27" gender="M" nation="BRA" license="391007" swrid="5602513" athleteid="2424" externalid="391007">
              <RESULTS>
                <RESULT eventid="1095" status="DNS" swimtime="00:00:00.00" resultid="2425" heatid="3441" lane="6" entrytime="00:02:17.17" entrycourse="SCM" />
                <RESULT eventid="1071" status="DNS" swimtime="00:00:00.00" resultid="2426" heatid="3402" lane="4" entrytime="00:01:04.24" entrycourse="SCM" />
                <RESULT eventid="1131" status="DNS" swimtime="00:00:00.00" resultid="2427" heatid="3473" lane="8" entrytime="00:00:51.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Sachser Rocha" birthdate="2008-07-09" gender="M" nation="BRA" license="330072" swrid="5600254" athleteid="1819" externalid="330072">
              <RESULTS>
                <RESULT eventid="1184" points="525" swimtime="00:00:26.95" resultid="1820" heatid="3518" lane="2" />
                <RESULT eventid="1216" points="487" swimtime="00:00:25.62" resultid="1821" heatid="3541" lane="4" />
                <RESULT eventid="1296" status="DSQ" swimtime="00:01:01.78" resultid="1822" heatid="3601" lane="4" entrytime="00:01:04.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Afonso Fowler" birthdate="2014-01-22" gender="M" nation="BRA" license="393264" swrid="5661338" athleteid="2530" externalid="393264">
              <RESULTS>
                <RESULT eventid="1095" points="80" swimtime="00:01:43.99" resultid="2531" heatid="3440" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="71" reactiontime="+85" swimtime="00:00:53.27" resultid="2532" heatid="3421" lane="5" />
                <RESULT eventid="1111" points="41" swimtime="00:01:02.85" resultid="2533" heatid="3457" lane="4" />
                <RESULT eventid="1131" points="101" swimtime="00:00:43.27" resultid="2534" heatid="3471" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="De Krinski" birthdate="2007-07-20" gender="M" nation="BRA" license="334494" swrid="5600148" athleteid="2690" externalid="334494">
              <RESULTS>
                <RESULT eventid="1200" points="517" reactiontime="+65" swimtime="00:01:00.21" resultid="2691" heatid="3532" lane="4" entrytime="00:01:00.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="478" reactiontime="+56" swimtime="00:00:28.27" resultid="2692" heatid="3593" lane="6" entrytime="00:00:28.40" entrycourse="SCM" />
                <RESULT eventid="1248" points="550" swimtime="00:00:54.72" resultid="2693" heatid="3580" lane="6" entrytime="00:00:56.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Cury" birthdate="2005-09-28" gender="M" nation="BRA" license="329251" swrid="5600270" athleteid="1952" externalid="329251" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1184" points="608" swimtime="00:00:25.67" resultid="1953" heatid="3522" lane="4" entrytime="00:00:25.83" entrycourse="SCM" />
                <RESULT eventid="1296" points="629" swimtime="00:00:55.75" resultid="1954" heatid="3602" lane="4" entrytime="00:00:56.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="590" swimtime="00:00:53.45" resultid="1955" heatid="3581" lane="3" entrytime="00:00:52.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Clivatti" birthdate="2010-05-24" gender="M" nation="BRA" license="368007" swrid="5600139" athleteid="2049" externalid="368007">
              <RESULTS>
                <RESULT eventid="1184" points="300" swimtime="00:00:32.47" resultid="2050" heatid="3517" lane="4" />
                <RESULT eventid="1152" points="461" swimtime="00:04:34.68" resultid="2051" heatid="3500" lane="2" entrytime="00:04:54.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                    <SPLIT distance="100" swimtime="00:01:05.15" />
                    <SPLIT distance="150" swimtime="00:01:39.88" />
                    <SPLIT distance="200" swimtime="00:02:14.50" />
                    <SPLIT distance="250" swimtime="00:02:49.82" />
                    <SPLIT distance="300" swimtime="00:03:25.17" />
                    <SPLIT distance="350" swimtime="00:04:00.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="394" swimtime="00:00:27.48" resultid="2052" heatid="3546" lane="5" entrytime="00:00:28.92" entrycourse="SCM" />
                <RESULT eventid="1296" points="303" swimtime="00:01:11.06" resultid="2053" heatid="3597" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="436" swimtime="00:00:59.10" resultid="2054" heatid="3578" lane="7" entrytime="00:01:03.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Pisani Ferreira" birthdate="2014-01-26" gender="M" nation="BRA" license="391017" swrid="5602570" athleteid="2441" externalid="391017">
              <RESULTS>
                <RESULT eventid="1095" points="92" swimtime="00:01:39.12" resultid="2442" heatid="3441" lane="4" entrytime="00:01:53.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="90" swimtime="00:00:55.62" resultid="2443" heatid="3404" lane="3" entrytime="00:00:58.89" entrycourse="SCM" />
                <RESULT eventid="1111" points="62" swimtime="00:00:54.75" resultid="2444" heatid="3459" lane="7" entrytime="00:00:53.73" entrycourse="SCM" />
                <RESULT eventid="1131" points="103" swimtime="00:00:42.99" resultid="2445" heatid="3473" lane="2" entrytime="00:00:48.89" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Wolf Macedo" birthdate="2012-01-27" gender="F" nation="BRA" license="369277" swrid="5602592" athleteid="2125" externalid="369277">
              <RESULTS>
                <RESULT eventid="1086" points="357" swimtime="00:02:35.45" resultid="2126" heatid="3428" lane="5" entrytime="00:02:33.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:14.96" />
                    <SPLIT distance="150" swimtime="00:01:55.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="272" reactiontime="+75" swimtime="00:00:38.96" resultid="2127" heatid="3406" lane="3" />
                <RESULT eventid="1118" points="236" swimtime="00:01:27.42" resultid="2128" heatid="3462" lane="5" entrytime="00:01:25.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="371" swimtime="00:00:31.89" resultid="2129" heatid="3477" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Della Villa Yang" birthdate="2012-10-08" gender="F" nation="BRA" license="369276" swrid="5588653" athleteid="2120" externalid="369276">
              <RESULTS>
                <RESULT eventid="1086" points="373" swimtime="00:02:33.24" resultid="2121" heatid="3428" lane="4" entrytime="00:02:32.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                    <SPLIT distance="100" swimtime="00:01:13.44" />
                    <SPLIT distance="150" swimtime="00:01:53.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="244" reactiontime="+79" swimtime="00:00:40.39" resultid="2122" heatid="3406" lane="6" />
                <RESULT eventid="1102" points="309" swimtime="00:01:23.52" resultid="2123" heatid="3444" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="354" swimtime="00:00:32.40" resultid="2124" heatid="3481" lane="6" entrytime="00:00:32.88" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Estela" lastname="Albuquerque" birthdate="2010-11-23" gender="F" nation="BRA" license="356344" swrid="5653285" athleteid="1898" externalid="356344">
              <RESULTS>
                <RESULT eventid="1144" points="419" swimtime="00:05:08.97" resultid="1899" heatid="3489" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.76" />
                    <SPLIT distance="100" swimtime="00:01:15.91" />
                    <SPLIT distance="150" swimtime="00:01:55.92" />
                    <SPLIT distance="200" swimtime="00:02:36.01" />
                    <SPLIT distance="250" swimtime="00:03:16.22" />
                    <SPLIT distance="300" swimtime="00:03:54.84" />
                    <SPLIT distance="350" swimtime="00:04:32.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="396" swimtime="00:00:31.22" resultid="1900" heatid="3533" lane="8" />
                <RESULT eventid="1192" points="350" reactiontime="+72" swimtime="00:01:17.83" resultid="1901" heatid="3526" lane="2" entrytime="00:01:20.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="257" swimtime="00:01:24.95" resultid="1902" heatid="3594" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="411" swimtime="00:01:07.58" resultid="1903" heatid="3568" lane="2" entrytime="00:01:09.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giuliana" lastname="Sovierzoski Ferreira" birthdate="2015-01-20" gender="F" nation="BRA" license="397168" swrid="5641776" athleteid="2550" externalid="397168">
              <RESULTS>
                <RESULT eventid="1092" points="49" swimtime="00:02:16.76" resultid="2551" heatid="3436" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="120" swimtime="00:00:57.38" resultid="2552" heatid="3401" lane="1" entrytime="00:01:04.11" entrycourse="SCM" />
                <RESULT eventid="1108" points="28" swimtime="00:01:19.82" resultid="2553" heatid="3452" lane="1" />
                <RESULT eventid="1128" points="42" swimtime="00:01:05.71" resultid="2554" heatid="3467" lane="6" entrytime="00:01:04.25" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Trevisan De Paula" birthdate="2014-01-27" gender="M" nation="BRA" license="377152" swrid="5602568" athleteid="2347" externalid="377152">
              <RESULTS>
                <RESULT eventid="1095" points="160" swimtime="00:01:22.47" resultid="2348" heatid="3442" lane="4" entrytime="00:01:20.83" entrycourse="SCM" />
                <RESULT eventid="1083" points="160" swimtime="00:00:40.67" resultid="2349" heatid="3423" lane="5" entrytime="00:00:42.05" entrycourse="SCM" />
                <RESULT eventid="1111" points="182" swimtime="00:00:38.31" resultid="2350" heatid="3459" lane="4" entrytime="00:00:39.08" entrycourse="SCM" />
                <RESULT eventid="1131" points="169" swimtime="00:00:36.41" resultid="2351" heatid="3474" lane="4" entrytime="00:00:35.93" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabelly" lastname="Sinnott" birthdate="2009-03-14" gender="F" nation="BRA" license="367255" swrid="5600258" athleteid="1776" externalid="367255">
              <RESULTS>
                <RESULT eventid="1144" points="540" swimtime="00:04:43.98" resultid="1777" heatid="3494" lane="3" entrytime="00:04:40.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="250" swimtime="00:02:54.56" />
                    <SPLIT distance="300" swimtime="00:03:30.93" />
                    <SPLIT distance="350" swimtime="00:04:07.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="541" swimtime="00:18:34.44" resultid="1778" heatid="3582" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.34" />
                    <SPLIT distance="100" swimtime="00:01:09.47" />
                    <SPLIT distance="150" swimtime="00:01:46.32" />
                    <SPLIT distance="200" swimtime="00:02:23.38" />
                    <SPLIT distance="250" swimtime="00:03:00.22" />
                    <SPLIT distance="300" swimtime="00:03:37.03" />
                    <SPLIT distance="350" swimtime="00:04:14.06" />
                    <SPLIT distance="400" swimtime="00:04:51.24" />
                    <SPLIT distance="450" swimtime="00:05:28.40" />
                    <SPLIT distance="500" swimtime="00:06:05.62" />
                    <SPLIT distance="550" swimtime="00:06:42.82" />
                    <SPLIT distance="600" swimtime="00:07:20.10" />
                    <SPLIT distance="650" swimtime="00:07:58.00" />
                    <SPLIT distance="700" swimtime="00:08:35.82" />
                    <SPLIT distance="750" swimtime="00:09:13.41" />
                    <SPLIT distance="800" swimtime="00:09:51.01" />
                    <SPLIT distance="850" swimtime="00:10:28.30" />
                    <SPLIT distance="900" swimtime="00:11:05.89" />
                    <SPLIT distance="950" swimtime="00:11:43.62" />
                    <SPLIT distance="1000" swimtime="00:12:21.10" />
                    <SPLIT distance="1050" swimtime="00:12:58.58" />
                    <SPLIT distance="1100" swimtime="00:13:36.16" />
                    <SPLIT distance="1150" swimtime="00:14:13.88" />
                    <SPLIT distance="1200" swimtime="00:14:51.74" />
                    <SPLIT distance="1250" swimtime="00:15:29.36" />
                    <SPLIT distance="1300" swimtime="00:16:07.28" />
                    <SPLIT distance="1350" swimtime="00:16:44.56" />
                    <SPLIT distance="1400" swimtime="00:17:21.45" />
                    <SPLIT distance="1450" swimtime="00:17:58.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Lacerda" birthdate="2011-05-09" gender="M" nation="BRA" license="366909" swrid="5602550" athleteid="2034" externalid="366909">
              <RESULTS>
                <RESULT eventid="1168" points="262" swimtime="00:01:26.34" resultid="2035" heatid="3510" lane="2" entrytime="00:01:30.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="338" swimtime="00:05:04.57" resultid="2036" heatid="3495" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                    <SPLIT distance="100" swimtime="00:01:14.45" />
                    <SPLIT distance="150" swimtime="00:01:53.96" />
                    <SPLIT distance="200" swimtime="00:02:33.63" />
                    <SPLIT distance="250" swimtime="00:03:13.20" />
                    <SPLIT distance="300" swimtime="00:03:51.50" />
                    <SPLIT distance="350" swimtime="00:04:30.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="291" swimtime="00:02:45.29" resultid="2037" heatid="3559" lane="5" entrytime="00:02:52.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:22.23" />
                    <SPLIT distance="150" swimtime="00:02:11.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="188" swimtime="00:01:23.40" resultid="2038" heatid="3598" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="281" swimtime="00:01:08.43" resultid="2039" heatid="3577" lane="2" entrytime="00:01:07.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cecilia Carvalho" birthdate="2014-10-30" gender="F" nation="BRA" license="391021" swrid="5602525" athleteid="2461" externalid="391021">
              <RESULTS>
                <RESULT eventid="1092" points="96" swimtime="00:01:49.60" resultid="2462" heatid="3437" lane="5" entrytime="00:01:57.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="95" reactiontime="+77" swimtime="00:00:55.17" resultid="2463" heatid="3418" lane="4" entrytime="00:00:57.44" entrycourse="SCM" />
                <RESULT eventid="1108" points="74" swimtime="00:00:58.05" resultid="2464" heatid="3455" lane="2" entrytime="00:00:59.77" entrycourse="SCM" />
                <RESULT eventid="1128" points="126" swimtime="00:00:45.63" resultid="2465" heatid="3468" lane="7" entrytime="00:00:50.75" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Albuquerque" birthdate="2012-11-16" gender="F" nation="BRA" license="369281" swrid="5602506" athleteid="2140" externalid="369281">
              <RESULTS>
                <RESULT eventid="1062" points="270" swimtime="00:01:36.38" resultid="2141" heatid="3394" lane="6" entrytime="00:01:41.44" entrycourse="SCM" />
                <RESULT eventid="1074" points="230" reactiontime="+73" swimtime="00:00:41.18" resultid="2142" heatid="3407" lane="2" />
                <RESULT eventid="1102" points="271" swimtime="00:01:27.28" resultid="2143" heatid="3445" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1118" points="202" swimtime="00:01:32.00" resultid="2144" heatid="3462" lane="3" entrytime="00:01:33.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Magalhaes Dabul" birthdate="2014-01-05" gender="M" nation="BRA" license="391023" swrid="5602555" athleteid="2466" externalid="391023">
              <RESULTS>
                <RESULT eventid="1095" points="94" swimtime="00:01:38.51" resultid="2467" heatid="3441" lane="3" entrytime="00:02:01.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="63" reactiontime="+101" swimtime="00:00:55.28" resultid="2468" heatid="3422" lane="4" entrytime="00:01:04.17" entrycourse="SCM" />
                <RESULT eventid="1111" points="70" swimtime="00:00:52.71" resultid="2469" heatid="3458" lane="5" entrytime="00:01:03.07" entrycourse="SCM" />
                <RESULT eventid="1131" points="102" swimtime="00:00:43.07" resultid="2470" heatid="3473" lane="1" entrytime="00:00:50.20" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinícius" lastname="Oliveira Cruz" birthdate="2005-07-02" gender="M" nation="BRA" license="298495" swrid="5653299" athleteid="2626" externalid="298495" level="ADTRISC">
              <RESULTS>
                <RESULT eventid="1152" points="720" swimtime="00:03:56.71" resultid="2627" heatid="3501" lane="4" entrytime="00:04:03.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                    <SPLIT distance="100" swimtime="00:00:56.74" />
                    <SPLIT distance="150" swimtime="00:01:26.59" />
                    <SPLIT distance="200" swimtime="00:01:57.00" />
                    <SPLIT distance="250" swimtime="00:02:26.66" />
                    <SPLIT distance="300" swimtime="00:02:56.52" />
                    <SPLIT distance="350" swimtime="00:03:26.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="566" swimtime="00:00:57.74" resultid="2628" heatid="3602" lane="3" entrytime="00:00:58.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="698" swimtime="00:00:50.54" resultid="2629" heatid="3581" lane="4" entrytime="00:00:51.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="646" swimtime="00:00:23.31" resultid="3614" heatid="3540" lane="6" late="yes" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Fontana Moraes" birthdate="2006-08-17" gender="M" nation="BRA" license="296593" swrid="5600163" athleteid="1807" externalid="296593">
              <RESULTS>
                <RESULT eventid="1200" points="184" reactiontime="+79" swimtime="00:01:24.85" resultid="1808" heatid="3530" lane="5" entrytime="00:01:19.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="296" swimtime="00:05:18.32" resultid="1809" heatid="3500" lane="7" entrytime="00:04:56.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:11.54" />
                    <SPLIT distance="150" swimtime="00:01:51.69" />
                    <SPLIT distance="200" swimtime="00:02:32.93" />
                    <SPLIT distance="250" swimtime="00:03:14.39" />
                    <SPLIT distance="300" swimtime="00:03:56.44" />
                    <SPLIT distance="350" swimtime="00:04:38.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="243" swimtime="00:00:32.28" resultid="1810" heatid="3546" lane="2" entrytime="00:00:29.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="De Macedo Martynychen" birthdate="2015-06-12" gender="F" nation="BRA" license="399681" swrid="5652885" athleteid="2570" externalid="399681">
              <RESULTS>
                <RESULT eventid="1092" points="44" swimtime="00:02:21.98" resultid="2571" heatid="3436" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="49" swimtime="00:01:08.54" resultid="2572" heatid="3418" lane="8" />
                <RESULT eventid="1108" points="48" swimtime="00:01:06.67" resultid="2573" heatid="3454" lane="6" />
                <RESULT eventid="1128" points="61" swimtime="00:00:58.15" resultid="2574" heatid="3466" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13038" nation="BRA" region="PR" clubid="1428" swrid="93759" name="Associação De Pais E Atletas De Natação Ws/Crb" shortname="Apan/Ws">
          <ATHLETES>
            <ATHLETE firstname="Isadora" lastname="Rosa Silva" birthdate="2011-03-25" gender="F" nation="BRA" license="392120" swrid="5602579" athleteid="1478" externalid="392120">
              <RESULTS>
                <RESULT eventid="1208" points="215" swimtime="00:00:38.24" resultid="1479" heatid="3534" lane="5" entrytime="00:00:45.57" entrycourse="SCM" />
                <RESULT eventid="1160" points="191" swimtime="00:01:48.27" resultid="1480" heatid="3502" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="167" swimtime="00:00:51.51" resultid="1481" heatid="3605" lane="1" entrytime="00:00:58.34" entrycourse="SCM" />
                <RESULT eventid="1240" points="194" swimtime="00:01:26.70" resultid="1482" heatid="3564" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabelly" lastname="Mendonca Bello" birthdate="2008-04-15" gender="F" nation="BRA" license="376996" swrid="5600217" athleteid="1444" externalid="376996" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1208" points="420" swimtime="00:00:30.61" resultid="1445" heatid="3538" lane="1" entrytime="00:00:31.58" entrycourse="SCM" />
                <RESULT eventid="1160" points="367" swimtime="00:01:27.07" resultid="1446" heatid="3504" lane="4" entrytime="00:01:32.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" status="DSQ" swimtime="00:02:54.06" resultid="1447" heatid="3552" lane="8" />
                <RESULT eventid="1304" points="335" swimtime="00:00:40.84" resultid="1448" heatid="3606" lane="7" entrytime="00:00:39.38" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Bobko Ganacim" birthdate="2013-08-02" gender="F" nation="BRA" license="397332" swrid="5641754" athleteid="1483" externalid="397332">
              <RESULTS>
                <RESULT eventid="1086" points="124" swimtime="00:03:41.17" resultid="1484" heatid="3425" lane="6" entrytime="00:04:09.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.79" />
                    <SPLIT distance="100" swimtime="00:01:43.10" />
                    <SPLIT distance="150" swimtime="00:02:41.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" reactiontime="+78" status="DSQ" swimtime="00:00:52.63" resultid="1485" heatid="3408" lane="7" entrytime="00:00:53.73" entrycourse="SCM" />
                <RESULT eventid="1138" points="157" swimtime="00:00:42.49" resultid="1486" heatid="3478" lane="2" entrytime="00:00:46.84" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Bernardi Iurk" birthdate="2012-04-14" gender="M" nation="BRA" license="406940" athleteid="1514" externalid="406940">
              <RESULTS>
                <RESULT eventid="1089" points="99" swimtime="00:03:34.66" resultid="1515" heatid="3430" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.74" />
                    <SPLIT distance="100" swimtime="00:01:42.28" />
                    <SPLIT distance="150" swimtime="00:02:40.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="88" reactiontime="+104" swimtime="00:00:49.67" resultid="1516" heatid="3411" lane="4" />
                <RESULT eventid="1141" points="117" swimtime="00:00:41.18" resultid="1517" heatid="3483" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="De Reginalda" birthdate="2011-07-22" gender="M" nation="BRA" license="400323" athleteid="1491" externalid="400323">
              <RESULTS>
                <RESULT eventid="1200" points="290" swimtime="00:01:13.00" resultid="1492" heatid="3529" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="135" swimtime="00:00:39.22" resultid="1493" heatid="3541" lane="2" />
                <RESULT eventid="1280" points="288" reactiontime="+47" swimtime="00:00:33.48" resultid="1494" heatid="3590" lane="2" />
                <RESULT eventid="1248" points="307" swimtime="00:01:06.42" resultid="1495" heatid="3571" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Sieck" birthdate="2011-01-20" gender="F" nation="BRA" license="382234" swrid="5602584" athleteid="1469" externalid="382234">
              <RESULTS>
                <RESULT eventid="1208" points="217" swimtime="00:00:38.10" resultid="1470" heatid="3534" lane="4" entrytime="00:00:41.95" entrycourse="SCM" />
                <RESULT eventid="1176" status="DSQ" swimtime="00:00:43.14" resultid="1471" heatid="3516" lane="1" entrytime="00:00:46.85" entrycourse="SCM" />
                <RESULT eventid="1288" points="121" swimtime="00:01:49.04" resultid="1472" heatid="3595" lane="7" entrytime="00:01:48.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="205" swimtime="00:01:25.15" resultid="1473" heatid="3564" lane="4" entrytime="00:01:33.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Da Reginalda" birthdate="2012-11-09" gender="M" nation="BRA" license="400275" athleteid="1496" externalid="400275">
              <RESULTS>
                <RESULT eventid="1089" points="186" swimtime="00:02:54.03" resultid="1497" heatid="3430" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                    <SPLIT distance="100" swimtime="00:01:19.47" />
                    <SPLIT distance="150" swimtime="00:02:04.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="183" swimtime="00:00:38.89" resultid="1498" heatid="3413" lane="8" />
                <RESULT eventid="1141" points="204" swimtime="00:00:34.21" resultid="1499" heatid="3482" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Dos Santos" birthdate="2013-06-26" gender="F" nation="BRA" license="387512" swrid="5588662" athleteid="1487" externalid="387512">
              <RESULTS>
                <RESULT eventid="1086" points="147" swimtime="00:03:28.77" resultid="1488" heatid="3424" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                    <SPLIT distance="100" swimtime="00:01:33.38" />
                    <SPLIT distance="150" swimtime="00:02:31.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="147" reactiontime="+104" swimtime="00:00:47.82" resultid="1489" heatid="3408" lane="1" entrytime="00:00:56.13" entrycourse="SCM" />
                <RESULT eventid="1138" points="186" swimtime="00:00:40.14" resultid="1490" heatid="3478" lane="8" entrytime="00:00:51.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Gramms Dallarosa" birthdate="2015-01-14" gender="F" nation="BRA" license="406868" athleteid="1507" externalid="406868">
              <RESULTS>
                <RESULT eventid="1080" points="61" swimtime="00:01:03.95" resultid="1508" heatid="3417" lane="7" />
                <RESULT eventid="1128" points="66" swimtime="00:00:56.57" resultid="1509" heatid="3465" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Zanchetta Silva" birthdate="2010-08-05" gender="F" nation="BRA" license="406865" athleteid="1504" externalid="406865">
              <RESULTS>
                <RESULT eventid="1208" points="160" swimtime="00:00:42.17" resultid="1505" heatid="3533" lane="5" />
                <RESULT eventid="1272" points="101" reactiontime="+59" swimtime="00:00:54.13" resultid="1506" heatid="3587" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Ferreira" birthdate="2012-12-29" gender="F" nation="BRA" license="382235" swrid="5602538" athleteid="1474" externalid="382235">
              <RESULTS>
                <RESULT eventid="1074" points="217" reactiontime="+76" swimtime="00:00:42.00" resultid="1475" heatid="3409" lane="6" entrytime="00:00:47.01" entrycourse="SCM" />
                <RESULT eventid="1118" points="145" swimtime="00:01:42.67" resultid="1476" heatid="3462" lane="6" entrytime="00:02:06.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="246" swimtime="00:00:36.57" resultid="1477" heatid="3479" lane="3" entrytime="00:00:41.04" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marjori" lastname="Leticia Oliveira" birthdate="2011-05-23" gender="F" nation="BRA" license="406869" athleteid="1510" externalid="406869">
              <RESULTS>
                <RESULT eventid="1208" points="206" swimtime="00:00:38.80" resultid="1511" heatid="3534" lane="7" />
                <RESULT eventid="1272" points="187" reactiontime="+54" swimtime="00:00:44.10" resultid="1512" heatid="3586" lane="3" />
                <RESULT eventid="1240" status="DSQ" swimtime="00:00:00.00" resultid="1513" heatid="3562" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Arceli Silva" birthdate="2008-03-04" gender="M" nation="BRA" license="331565" swrid="5385686" athleteid="1449" externalid="331565" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1200" points="332" reactiontime="+72" swimtime="00:01:09.78" resultid="1450" heatid="3531" lane="6" entrytime="00:01:11.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="374" swimtime="00:00:30.18" resultid="1451" heatid="3519" lane="3" />
                <RESULT eventid="1232" points="295" swimtime="00:02:44.56" resultid="1452" heatid="3560" lane="8" entrytime="00:02:45.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                    <SPLIT distance="100" swimtime="00:01:11.36" />
                    <SPLIT distance="150" swimtime="00:02:04.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="340" swimtime="00:01:08.41" resultid="1453" heatid="3601" lane="1" entrytime="00:01:10.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Zeclhynski Silva" birthdate="2006-09-14" gender="F" nation="BRA" license="330727" swrid="5600283" athleteid="1429" externalid="330727" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1208" points="593" swimtime="00:00:27.29" resultid="1430" heatid="3539" lane="4" entrytime="00:00:27.37" entrycourse="SCM" />
                <RESULT eventid="1192" points="583" reactiontime="+66" swimtime="00:01:05.68" resultid="1431" heatid="3527" lane="4" entrytime="00:01:04.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="610" reactiontime="+67" swimtime="00:00:29.77" resultid="1432" heatid="3589" lane="4" entrytime="00:00:29.75" entrycourse="SCM" />
                <RESULT eventid="1240" points="592" swimtime="00:00:59.84" resultid="1433" heatid="3570" lane="4" entrytime="00:01:00.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Daniele Silva" birthdate="2010-07-06" gender="F" nation="BRA" license="359593" swrid="5588628" athleteid="1454" externalid="359593" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1208" points="442" swimtime="00:00:30.08" resultid="1455" heatid="3538" lane="8" entrytime="00:00:31.69" entrycourse="SCM" />
                <RESULT eventid="1192" points="383" swimtime="00:01:15.55" resultid="1456" heatid="3526" lane="8" entrytime="00:01:21.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="306" swimtime="00:00:42.08" resultid="1457" heatid="3604" lane="7" />
                <RESULT eventid="1240" points="442" swimtime="00:01:05.94" resultid="1458" heatid="3566" lane="2" entrytime="00:01:14.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Da Costa Riekes" birthdate="2008-06-19" gender="F" nation="BRA" license="331686" swrid="5600143" athleteid="1439" externalid="331686" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1208" points="467" swimtime="00:00:29.55" resultid="1440" heatid="3539" lane="2" entrytime="00:00:30.12" entrycourse="SCM" />
                <RESULT eventid="1176" points="443" swimtime="00:00:31.98" resultid="1441" heatid="3516" lane="3" entrytime="00:00:33.88" entrycourse="SCM" />
                <RESULT eventid="1288" points="354" swimtime="00:01:16.36" resultid="1442" heatid="3596" lane="2" entrytime="00:01:14.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="484" swimtime="00:01:03.97" resultid="1443" heatid="3570" lane="8" entrytime="00:01:04.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Alexandre Azevedo" birthdate="2008-05-20" gender="M" nation="BRA" license="398694" athleteid="1459" externalid="398694">
              <RESULTS>
                <RESULT eventid="1168" points="192" swimtime="00:01:35.79" resultid="1460" heatid="3507" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="275" swimtime="00:00:30.98" resultid="1461" heatid="3545" lane="6" entrytime="00:00:31.23" entrycourse="SCM" />
                <RESULT eventid="1312" points="188" swimtime="00:00:43.48" resultid="1462" heatid="3609" lane="8" />
                <RESULT eventid="1248" points="242" swimtime="00:01:11.91" resultid="1463" heatid="3572" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leon" lastname="Bernardo Bello" birthdate="2014-11-23" gender="M" nation="BRA" license="400324" athleteid="1500" externalid="400324">
              <RESULTS>
                <RESULT eventid="1095" points="100" swimtime="00:01:36.32" resultid="1501" heatid="3439" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="101" reactiontime="+86" swimtime="00:00:47.45" resultid="1502" heatid="3420" lane="5" />
                <RESULT eventid="1131" points="120" swimtime="00:00:40.80" resultid="1503" heatid="3471" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Reis" birthdate="2008-04-07" gender="F" nation="BRA" license="378820" swrid="5600243" athleteid="1464" externalid="378820" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1208" points="215" swimtime="00:00:38.25" resultid="1465" heatid="3535" lane="5" entrytime="00:00:38.42" entrycourse="SCM" />
                <RESULT eventid="1176" points="168" swimtime="00:00:44.10" resultid="1466" heatid="3515" lane="2" />
                <RESULT eventid="1272" points="193" swimtime="00:00:43.66" resultid="1467" heatid="3588" lane="8" entrytime="00:00:45.21" entrycourse="SCM" />
                <RESULT eventid="1240" points="222" swimtime="00:01:22.87" resultid="1468" heatid="3565" lane="2" entrytime="00:01:23.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonia" lastname="Adam  Fracaro" birthdate="2010-04-27" gender="F" nation="BRA" license="382212" swrid="5588512" athleteid="1434" externalid="382212">
              <RESULTS>
                <RESULT eventid="1144" points="321" swimtime="00:05:37.79" resultid="1435" heatid="3492" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.83" />
                    <SPLIT distance="100" swimtime="00:01:16.20" />
                    <SPLIT distance="150" swimtime="00:01:58.52" />
                    <SPLIT distance="200" swimtime="00:02:41.68" />
                    <SPLIT distance="250" swimtime="00:03:26.36" />
                    <SPLIT distance="300" swimtime="00:04:10.52" />
                    <SPLIT distance="350" swimtime="00:04:56.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="327" swimtime="00:00:33.28" resultid="1436" heatid="3536" lane="5" entrytime="00:00:34.12" entrycourse="SCM" />
                <RESULT eventid="1272" points="260" reactiontime="+70" swimtime="00:00:39.53" resultid="1437" heatid="3588" lane="7" entrytime="00:00:41.56" entrycourse="SCM" />
                <RESULT eventid="1240" points="339" swimtime="00:01:12.04" resultid="1438" heatid="3566" lane="5" entrytime="00:01:14.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16131" nation="BRA" region="PR" clubid="2737" swrid="93766" name="Associação Nadar Colombo" shortname="Equipe Nadar">
          <ATHLETES>
            <ATHLETE firstname="Tayna" lastname="Macedo Gabardo" birthdate="2012-12-01" gender="F" nation="BRA" license="406704" athleteid="2770" externalid="406704">
              <RESULTS>
                <RESULT eventid="1074" points="144" reactiontime="+77" swimtime="00:00:48.10" resultid="2771" heatid="3407" lane="4" />
                <RESULT eventid="1138" points="174" swimtime="00:00:41.01" resultid="2772" heatid="3476" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Pavin" birthdate="2008-07-17" gender="F" nation="BRA" license="406703" athleteid="2768" externalid="406703">
              <RESULTS>
                <RESULT eventid="1208" points="283" swimtime="00:00:34.92" resultid="2769" heatid="3533" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Luiz Sartori" birthdate="2008-04-07" gender="M" nation="BRA" license="384742" swrid="5622287" athleteid="2749" externalid="384742">
              <RESULTS>
                <RESULT eventid="1184" points="379" swimtime="00:00:30.03" resultid="2750" heatid="3517" lane="3" />
                <RESULT eventid="1216" points="409" swimtime="00:00:27.15" resultid="2751" heatid="3548" lane="8" entrytime="00:00:27.79" entrycourse="SCM" />
                <RESULT eventid="1280" points="311" swimtime="00:00:32.60" resultid="2752" heatid="3591" lane="8" />
                <RESULT eventid="1248" points="431" swimtime="00:00:59.33" resultid="2753" heatid="3571" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaylaine" lastname="Sofia Vargas Bueno" birthdate="2006-11-28" gender="F" nation="BRA" license="384739" swrid="5622307" athleteid="2741" externalid="384739">
              <RESULTS>
                <RESULT eventid="1208" points="297" swimtime="00:00:34.36" resultid="2742" heatid="3536" lane="4" entrytime="00:00:33.87" entrycourse="SCM" />
                <RESULT eventid="1160" points="216" swimtime="00:01:43.79" resultid="2743" heatid="3504" lane="7" entrytime="00:01:40.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="257" swimtime="00:00:44.62" resultid="2744" heatid="3604" lane="1" />
                <RESULT eventid="1240" points="304" swimtime="00:01:14.69" resultid="2745" heatid="3566" lane="7" entrytime="00:01:14.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Krik" birthdate="2010-11-24" gender="F" nation="BRA" license="406702" athleteid="2765" externalid="406702">
              <RESULTS>
                <RESULT eventid="1208" points="169" swimtime="00:00:41.41" resultid="2766" heatid="3534" lane="6" />
                <RESULT eventid="1304" points="150" swimtime="00:00:53.29" resultid="2767" heatid="3603" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Carvalho" birthdate="2011-10-20" gender="F" nation="BRA" license="399927" swrid="5652882" athleteid="2758" externalid="399927">
              <RESULTS>
                <RESULT eventid="1208" points="256" swimtime="00:00:36.07" resultid="2759" heatid="3535" lane="6" entrytime="00:00:39.40" entrycourse="SCM" />
                <RESULT eventid="1160" points="232" swimtime="00:01:41.37" resultid="2760" heatid="3503" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="210" swimtime="00:00:47.72" resultid="2761" heatid="3605" lane="2" entrytime="00:00:51.67" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Felipe Glir" birthdate="2006-10-11" gender="M" nation="BRA" license="384741" swrid="5622280" athleteid="2746" externalid="384741">
              <RESULTS>
                <RESULT eventid="1216" points="366" swimtime="00:00:28.16" resultid="2747" heatid="3548" lane="7" entrytime="00:00:27.68" entrycourse="SCM" />
                <RESULT eventid="1248" points="344" swimtime="00:01:03.97" resultid="2748" heatid="3578" lane="1" entrytime="00:01:04.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Rafael D Agostin Batistao" birthdate="2008-05-13" gender="M" nation="BRA" license="384738" swrid="5622300" athleteid="2738" externalid="384738">
              <RESULTS>
                <RESULT eventid="1168" points="326" swimtime="00:01:20.32" resultid="2739" heatid="3508" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="311" swimtime="00:00:36.82" resultid="2740" heatid="3609" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Glir" birthdate="2010-07-01" gender="M" nation="BRA" license="406701" athleteid="2762" externalid="406701">
              <RESULTS>
                <RESULT eventid="1312" points="150" swimtime="00:00:46.87" resultid="2763" heatid="3608" lane="8" />
                <RESULT eventid="1248" points="203" swimtime="00:01:16.22" resultid="2764" heatid="3573" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Rosa De Souza" birthdate="2009-01-01" gender="F" nation="BRA" license="399926" swrid="5653301" athleteid="2754" externalid="399926">
              <RESULTS>
                <RESULT eventid="1208" points="288" swimtime="00:00:34.71" resultid="2755" heatid="3534" lane="3" />
                <RESULT eventid="1304" points="235" swimtime="00:00:45.92" resultid="2756" heatid="3603" lane="3" />
                <RESULT eventid="1240" points="255" swimtime="00:01:19.14" resultid="2757" heatid="3564" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13068" nation="BRA" region="PR" clubid="2826" swrid="93787" name="Sociedade Morgenau" shortname="Morgenau">
          <ATHLETES>
            <ATHLETE firstname="Herick" lastname="Dos Santos" birthdate="2009-06-11" gender="M" nation="BRA" license="406724" athleteid="3030" externalid="406724">
              <RESULTS>
                <RESULT eventid="1152" points="116" swimtime="00:07:14.12" resultid="3031" heatid="3497" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.60" />
                    <SPLIT distance="100" swimtime="00:01:36.59" />
                    <SPLIT distance="150" swimtime="00:02:33.38" />
                    <SPLIT distance="200" swimtime="00:03:31.44" />
                    <SPLIT distance="250" swimtime="00:04:29.75" />
                    <SPLIT distance="300" swimtime="00:05:26.25" />
                    <SPLIT distance="350" swimtime="00:06:21.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="171" swimtime="00:00:36.26" resultid="3032" heatid="3540" lane="5" />
                <RESULT eventid="1280" points="116" reactiontime="+69" swimtime="00:00:45.22" resultid="3033" heatid="3590" lane="4" />
                <RESULT eventid="1248" points="136" swimtime="00:01:27.00" resultid="3034" heatid="3572" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Liz Skowronski" birthdate="2008-01-24" gender="F" nation="BRA" license="358245" swrid="5600202" athleteid="2835" externalid="358245">
              <RESULTS>
                <RESULT eventid="1144" points="386" swimtime="00:05:17.55" resultid="2836" heatid="3493" lane="7" entrytime="00:05:27.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:15.07" />
                    <SPLIT distance="150" swimtime="00:01:54.44" />
                    <SPLIT distance="200" swimtime="00:02:34.98" />
                    <SPLIT distance="250" swimtime="00:03:15.27" />
                    <SPLIT distance="300" swimtime="00:03:56.58" />
                    <SPLIT distance="350" swimtime="00:04:37.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="353" reactiontime="+68" swimtime="00:01:17.65" resultid="2837" heatid="3526" lane="4" entrytime="00:01:17.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="343" swimtime="00:02:53.95" resultid="2838" heatid="3555" lane="1" entrytime="00:02:57.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                    <SPLIT distance="100" swimtime="00:01:22.14" />
                    <SPLIT distance="150" swimtime="00:02:14.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="259" swimtime="00:01:24.69" resultid="2839" heatid="3594" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="310" swimtime="00:00:37.30" resultid="2840" heatid="3589" lane="8" entrytime="00:00:35.92" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduarda" lastname="Azevedo Birsneek" birthdate="2010-03-31" gender="F" nation="BRA" license="391145" swrid="5389427" athleteid="2944" externalid="391145">
              <RESULTS>
                <RESULT eventid="1144" points="164" swimtime="00:07:02.45" resultid="2945" heatid="3490" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.34" />
                    <SPLIT distance="100" swimtime="00:01:36.42" />
                    <SPLIT distance="150" swimtime="00:02:29.69" />
                    <SPLIT distance="200" swimtime="00:03:23.88" />
                    <SPLIT distance="250" swimtime="00:04:19.18" />
                    <SPLIT distance="300" swimtime="00:05:13.35" />
                    <SPLIT distance="350" swimtime="00:06:07.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="186" reactiontime="+74" swimtime="00:01:36.12" resultid="2946" heatid="3523" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="123" swimtime="00:00:49.01" resultid="2947" heatid="3515" lane="3" />
                <RESULT eventid="1272" points="199" reactiontime="+52" swimtime="00:00:43.18" resultid="2948" heatid="3587" lane="3" entrytime="00:00:52.43" entrycourse="SCM" />
                <RESULT eventid="1240" points="158" swimtime="00:01:32.84" resultid="2949" heatid="3564" lane="3" entrytime="00:01:46.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Vitoria De Lima" birthdate="2011-06-10" gender="F" nation="BRA" license="400090" swrid="5652904" athleteid="2991" externalid="400090">
              <RESULTS>
                <RESULT eventid="1208" points="165" swimtime="00:00:41.80" resultid="2992" heatid="3535" lane="8" entrytime="00:00:41.69" entrycourse="SCM" />
                <RESULT eventid="1272" status="DNS" swimtime="00:00:00.00" resultid="2993" heatid="3586" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Capoia Soares" birthdate="2011-11-07" gender="M" nation="BRA" license="393257" swrid="5616440" athleteid="2966" externalid="393257">
              <RESULTS>
                <RESULT eventid="1200" points="75" reactiontime="+107" swimtime="00:01:54.34" resultid="2967" heatid="3528" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="56" swimtime="00:00:56.74" resultid="2968" heatid="3519" lane="6" />
                <RESULT eventid="1280" reactiontime="+79" status="DSQ" swimtime="00:00:49.49" resultid="2969" heatid="3592" lane="2" entrytime="00:00:55.98" entrycourse="SCM" />
                <RESULT eventid="1248" points="96" swimtime="00:01:37.82" resultid="2970" heatid="3575" lane="1" entrytime="00:01:48.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Isabel Santos" birthdate="2005-12-20" gender="F" nation="BRA" license="391141" swrid="5600191" athleteid="2929" externalid="391141">
              <RESULTS>
                <RESULT eventid="1144" points="247" swimtime="00:06:08.31" resultid="2930" heatid="3489" lane="3" />
                <RESULT eventid="1176" points="237" swimtime="00:00:39.35" resultid="2931" heatid="3516" lane="8" entrytime="00:00:48.02" entrycourse="SCM" />
                <RESULT eventid="1224" status="DNS" swimtime="00:00:00.00" resultid="2932" heatid="3552" lane="4" />
                <RESULT eventid="1240" points="282" swimtime="00:01:16.58" resultid="2933" heatid="3565" lane="1" entrytime="00:01:27.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Andreis Ramos" birthdate="2007-03-26" gender="M" nation="BRA" license="406719" athleteid="3005" externalid="406719">
              <RESULTS>
                <RESULT eventid="1184" points="279" swimtime="00:00:33.28" resultid="3006" heatid="3519" lane="7" />
                <RESULT eventid="1216" points="337" swimtime="00:00:28.96" resultid="3007" heatid="3542" lane="4" />
                <RESULT eventid="1312" status="DSQ" swimtime="00:00:42.18" resultid="3008" heatid="3609" lane="6" />
                <RESULT eventid="1280" points="214" reactiontime="+40" swimtime="00:00:36.91" resultid="3009" heatid="3591" lane="4" />
                <RESULT eventid="1248" points="309" swimtime="00:01:06.29" resultid="3010" heatid="3571" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jhenyffer" lastname="Stefany De Santana Szaida" birthdate="2006-09-16" gender="F" nation="BRA" license="369326" swrid="5600264" athleteid="2882" externalid="369326">
              <RESULTS>
                <RESULT eventid="1176" points="320" swimtime="00:00:35.64" resultid="2883" heatid="3516" lane="6" entrytime="00:00:36.70" entrycourse="SCM" />
                <RESULT eventid="1224" points="264" swimtime="00:03:09.78" resultid="2884" heatid="3553" lane="5" entrytime="00:03:10.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                    <SPLIT distance="100" swimtime="00:01:26.88" />
                    <SPLIT distance="150" swimtime="00:02:23.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="240" reactiontime="+65" swimtime="00:00:40.59" resultid="2885" heatid="3588" lane="3" entrytime="00:00:39.63" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mayara" lastname="Fieber" birthdate="2008-08-20" gender="F" nation="BRA" license="391147" swrid="5600161" athleteid="2956" externalid="391147">
              <RESULTS>
                <RESULT eventid="1208" points="337" swimtime="00:00:32.93" resultid="2957" heatid="3536" lane="1" entrytime="00:00:36.50" entrycourse="SCM" />
                <RESULT eventid="1192" points="258" reactiontime="+67" swimtime="00:01:26.14" resultid="2958" heatid="3525" lane="1" entrytime="00:01:36.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="272" swimtime="00:00:43.76" resultid="2959" heatid="3603" lane="6" />
                <RESULT eventid="1240" points="318" swimtime="00:01:13.61" resultid="2960" heatid="3565" lane="7" entrytime="00:01:23.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Paes Pereira" birthdate="2013-03-11" gender="M" nation="BRA" license="391137" swrid="5602567" athleteid="2921" externalid="391137">
              <RESULTS>
                <RESULT eventid="1141" points="92" swimtime="00:00:44.51" resultid="2922" heatid="3483" lane="5" entrytime="00:00:46.38" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stella" lastname="Magalhaes Birnbaum" birthdate="2009-05-14" gender="F" nation="BRA" license="399684" swrid="5653298" athleteid="2987" externalid="399684">
              <RESULTS>
                <RESULT eventid="1208" points="359" swimtime="00:00:32.24" resultid="2988" heatid="3536" lane="7" entrytime="00:00:35.20" entrycourse="SCM" />
                <RESULT eventid="1192" points="285" reactiontime="+88" swimtime="00:01:23.37" resultid="2989" heatid="3523" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="338" swimtime="00:01:12.10" resultid="2990" heatid="3566" lane="8" entrytime="00:01:17.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Portella Da Silva" birthdate="2010-07-19" gender="M" nation="BRA" license="399534" athleteid="2857" externalid="399534">
              <RESULTS>
                <RESULT eventid="1312" status="DSQ" swimtime="00:00:45.40" resultid="2858" heatid="3610" lane="8" />
                <RESULT eventid="1280" points="132" reactiontime="+48" swimtime="00:00:43.40" resultid="2859" heatid="3591" lane="6" />
                <RESULT eventid="1248" points="144" swimtime="00:01:25.51" resultid="2860" heatid="3572" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabryel" lastname="Denk" birthdate="2011-05-09" gender="M" nation="BRA" license="391138" swrid="5602531" athleteid="2923" externalid="391138">
              <RESULTS>
                <RESULT eventid="1152" points="266" swimtime="00:05:29.92" resultid="2924" heatid="3498" lane="2" entrytime="00:05:52.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.06" />
                    <SPLIT distance="100" swimtime="00:01:19.46" />
                    <SPLIT distance="150" swimtime="00:02:01.12" />
                    <SPLIT distance="200" swimtime="00:02:43.74" />
                    <SPLIT distance="250" swimtime="00:03:25.24" />
                    <SPLIT distance="300" swimtime="00:04:07.27" />
                    <SPLIT distance="350" swimtime="00:04:49.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="216" swimtime="00:00:33.55" resultid="2925" heatid="3544" lane="2" entrytime="00:00:36.83" entrycourse="SCM" />
                <RESULT eventid="1312" points="137" swimtime="00:00:48.31" resultid="2926" heatid="3610" lane="1" entrytime="00:00:51.95" entrycourse="SCM" />
                <RESULT eventid="1280" points="180" reactiontime="+50" swimtime="00:00:39.10" resultid="2927" heatid="3590" lane="5" />
                <RESULT eventid="1264" points="289" swimtime="00:21:20.90" resultid="2928" heatid="3585" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                    <SPLIT distance="100" swimtime="00:01:18.94" />
                    <SPLIT distance="150" swimtime="00:02:02.06" />
                    <SPLIT distance="250" swimtime="00:03:28.83" />
                    <SPLIT distance="300" swimtime="00:04:12.54" />
                    <SPLIT distance="350" swimtime="00:04:55.23" />
                    <SPLIT distance="400" swimtime="00:05:39.06" />
                    <SPLIT distance="450" swimtime="00:06:21.12" />
                    <SPLIT distance="500" swimtime="00:07:03.39" />
                    <SPLIT distance="550" swimtime="00:07:46.49" />
                    <SPLIT distance="600" swimtime="00:08:29.51" />
                    <SPLIT distance="650" swimtime="00:09:13.00" />
                    <SPLIT distance="700" swimtime="00:09:55.51" />
                    <SPLIT distance="750" swimtime="00:10:38.91" />
                    <SPLIT distance="800" swimtime="00:11:22.04" />
                    <SPLIT distance="850" swimtime="00:12:04.98" />
                    <SPLIT distance="900" swimtime="00:12:47.92" />
                    <SPLIT distance="950" swimtime="00:13:30.84" />
                    <SPLIT distance="1000" swimtime="00:14:13.81" />
                    <SPLIT distance="1050" swimtime="00:14:56.42" />
                    <SPLIT distance="1100" swimtime="00:15:39.54" />
                    <SPLIT distance="1150" swimtime="00:16:22.64" />
                    <SPLIT distance="1200" swimtime="00:17:05.42" />
                    <SPLIT distance="1250" swimtime="00:17:48.43" />
                    <SPLIT distance="1300" swimtime="00:18:31.70" />
                    <SPLIT distance="1350" swimtime="00:19:14.14" />
                    <SPLIT distance="1400" swimtime="00:19:57.31" />
                    <SPLIT distance="1450" swimtime="00:20:40.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Alves" birthdate="2012-10-12" gender="M" nation="BRA" license="369324" swrid="5588674" athleteid="2877" externalid="369324">
              <RESULTS>
                <RESULT eventid="1089" points="209" swimtime="00:02:47.32" resultid="2878" heatid="3433" lane="4" entrytime="00:02:50.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.17" />
                    <SPLIT distance="100" swimtime="00:01:20.43" />
                    <SPLIT distance="150" swimtime="00:02:06.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="228" reactiontime="+69" swimtime="00:00:36.15" resultid="2879" heatid="3415" lane="4" entrytime="00:00:36.40" entrycourse="SCM" />
                <RESULT eventid="1105" points="175" swimtime="00:01:27.94" resultid="2880" heatid="3448" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="234" swimtime="00:00:32.68" resultid="2881" heatid="3487" lane="3" entrytime="00:00:33.60" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Kozera Chiarato" birthdate="2010-05-28" gender="M" nation="BRA" license="406722" athleteid="3021" externalid="406722">
              <RESULTS>
                <RESULT eventid="1184" points="243" swimtime="00:00:34.84" resultid="3022" heatid="3517" lane="5" />
                <RESULT eventid="1168" points="200" swimtime="00:01:34.38" resultid="3023" heatid="3508" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="240" swimtime="00:00:32.43" resultid="3024" heatid="3543" lane="8" />
                <RESULT eventid="1312" points="195" swimtime="00:00:42.98" resultid="3025" heatid="3608" lane="3" />
                <RESULT eventid="1248" points="214" swimtime="00:01:14.88" resultid="3026" heatid="3574" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Matos Oliveira" birthdate="2007-10-26" gender="M" nation="BRA" license="391136" swrid="5600215" athleteid="2915" externalid="391136">
              <RESULTS>
                <RESULT eventid="1184" points="261" swimtime="00:00:34.03" resultid="2916" heatid="3521" lane="8" entrytime="00:00:40.49" entrycourse="SCM" />
                <RESULT eventid="1152" points="351" swimtime="00:05:00.74" resultid="2917" heatid="3499" lane="8" entrytime="00:05:31.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                    <SPLIT distance="100" swimtime="00:01:09.20" />
                    <SPLIT distance="150" swimtime="00:01:48.01" />
                    <SPLIT distance="200" swimtime="00:02:27.11" />
                    <SPLIT distance="250" swimtime="00:03:05.97" />
                    <SPLIT distance="300" swimtime="00:03:44.42" />
                    <SPLIT distance="350" swimtime="00:04:23.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="258" swimtime="00:02:52.17" resultid="2918" heatid="3557" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:19.87" />
                    <SPLIT distance="150" swimtime="00:02:13.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="209" swimtime="00:00:42.00" resultid="2919" heatid="3608" lane="2" />
                <RESULT eventid="1264" points="339" swimtime="00:20:13.88" resultid="2920" heatid="3583" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                    <SPLIT distance="100" swimtime="00:01:13.45" />
                    <SPLIT distance="150" swimtime="00:01:53.83" />
                    <SPLIT distance="200" swimtime="00:02:34.31" />
                    <SPLIT distance="250" swimtime="00:03:15.34" />
                    <SPLIT distance="300" swimtime="00:03:56.18" />
                    <SPLIT distance="350" swimtime="00:04:36.87" />
                    <SPLIT distance="400" swimtime="00:05:17.69" />
                    <SPLIT distance="450" swimtime="00:05:58.51" />
                    <SPLIT distance="500" swimtime="00:06:39.24" />
                    <SPLIT distance="550" swimtime="00:07:20.32" />
                    <SPLIT distance="600" swimtime="00:08:01.32" />
                    <SPLIT distance="650" swimtime="00:08:42.74" />
                    <SPLIT distance="700" swimtime="00:09:23.41" />
                    <SPLIT distance="750" swimtime="00:10:04.40" />
                    <SPLIT distance="800" swimtime="00:10:45.53" />
                    <SPLIT distance="850" swimtime="00:11:25.94" />
                    <SPLIT distance="900" swimtime="00:12:07.36" />
                    <SPLIT distance="950" swimtime="00:12:48.52" />
                    <SPLIT distance="1000" swimtime="00:13:29.46" />
                    <SPLIT distance="1050" swimtime="00:14:10.48" />
                    <SPLIT distance="1100" swimtime="00:14:51.31" />
                    <SPLIT distance="1150" swimtime="00:15:32.45" />
                    <SPLIT distance="1200" swimtime="00:16:13.18" />
                    <SPLIT distance="1250" swimtime="00:16:54.52" />
                    <SPLIT distance="1300" swimtime="00:17:35.49" />
                    <SPLIT distance="1350" swimtime="00:18:16.62" />
                    <SPLIT distance="1400" swimtime="00:18:56.91" />
                    <SPLIT distance="1450" swimtime="00:19:36.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Bora" birthdate="2005-01-06" gender="F" nation="BRA" license="358252" swrid="5600153" athleteid="2872" externalid="358252">
              <RESULTS>
                <RESULT eventid="1144" points="365" swimtime="00:05:23.49" resultid="2873" heatid="3489" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="100" swimtime="00:01:16.64" />
                    <SPLIT distance="150" swimtime="00:01:57.83" />
                    <SPLIT distance="200" swimtime="00:02:39.07" />
                    <SPLIT distance="250" swimtime="00:03:20.33" />
                    <SPLIT distance="300" swimtime="00:04:02.10" />
                    <SPLIT distance="350" swimtime="00:04:43.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="301" reactiontime="+66" swimtime="00:01:21.84" resultid="2874" heatid="3526" lane="1" entrytime="00:01:20.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="307" swimtime="00:03:00.47" resultid="2875" heatid="3555" lane="7" entrytime="00:02:56.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.81" />
                    <SPLIT distance="100" swimtime="00:01:24.68" />
                    <SPLIT distance="150" swimtime="00:02:20.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="265" swimtime="00:01:24.10" resultid="2876" heatid="3595" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cecilia Carstens" birthdate="2014-02-22" gender="F" nation="BRA" license="406721" athleteid="3016" externalid="406721">
              <RESULTS>
                <RESULT eventid="1080" points="70" reactiontime="+80" swimtime="00:01:01.24" resultid="3017" heatid="3416" lane="3" />
                <RESULT eventid="1068" points="97" swimtime="00:01:01.55" resultid="3018" heatid="3399" lane="5" />
                <RESULT eventid="1108" points="48" swimtime="00:01:07.06" resultid="3019" heatid="3454" lane="7" />
                <RESULT eventid="1128" points="60" swimtime="00:00:58.38" resultid="3020" heatid="3466" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maryana" lastname="Lemos Carvalho" birthdate="2014-02-10" gender="F" nation="BRA" license="406718" athleteid="3001" externalid="406718">
              <RESULTS>
                <RESULT eventid="1092" points="88" swimtime="00:01:52.96" resultid="3002" heatid="3435" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="67" reactiontime="+82" swimtime="00:01:02.13" resultid="3003" heatid="3417" lane="3" />
                <RESULT eventid="1128" points="102" swimtime="00:00:48.98" resultid="3004" heatid="3465" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Nitz Costa" birthdate="2015-02-09" gender="F" nation="BRA" license="397328" swrid="5641773" athleteid="2982" externalid="397328">
              <RESULTS>
                <RESULT eventid="1092" points="162" swimtime="00:01:32.02" resultid="2983" heatid="3436" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="160" reactiontime="+75" swimtime="00:00:46.43" resultid="2984" heatid="3419" lane="5" entrytime="00:00:49.83" entrycourse="SCM" />
                <RESULT eventid="1108" points="128" swimtime="00:00:48.30" resultid="2985" heatid="3455" lane="8" entrytime="00:01:02.67" entrycourse="SCM" />
                <RESULT eventid="1128" points="146" swimtime="00:00:43.46" resultid="2986" heatid="3468" lane="6" entrytime="00:00:46.87" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Lima" birthdate="2006-12-03" gender="M" nation="BRA" license="366749" swrid="5600201" athleteid="2896" externalid="366749">
              <RESULTS>
                <RESULT eventid="1152" points="519" swimtime="00:04:24.10" resultid="2897" heatid="3496" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                    <SPLIT distance="100" swimtime="00:01:02.88" />
                    <SPLIT distance="150" swimtime="00:01:36.82" />
                    <SPLIT distance="200" swimtime="00:02:10.71" />
                    <SPLIT distance="250" swimtime="00:02:44.40" />
                    <SPLIT distance="300" swimtime="00:03:18.45" />
                    <SPLIT distance="350" swimtime="00:03:51.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="530" swimtime="00:00:24.91" resultid="2898" heatid="3550" lane="7" entrytime="00:00:25.30" entrycourse="SCM" />
                <RESULT eventid="1296" points="462" swimtime="00:01:01.79" resultid="2899" heatid="3602" lane="1" entrytime="00:01:02.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="549" swimtime="00:00:54.75" resultid="2900" heatid="3580" lane="4" entrytime="00:00:55.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Madalena De Lima" birthdate="2006-05-04" gender="M" nation="BRA" license="307786" swrid="5600206" athleteid="2832" externalid="307786">
              <RESULTS>
                <RESULT eventid="1152" points="461" swimtime="00:04:34.57" resultid="2833" heatid="3501" lane="7" entrytime="00:04:37.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.31" />
                    <SPLIT distance="100" swimtime="00:01:02.61" />
                    <SPLIT distance="150" swimtime="00:01:36.40" />
                    <SPLIT distance="200" swimtime="00:02:10.64" />
                    <SPLIT distance="250" swimtime="00:02:45.83" />
                    <SPLIT distance="300" swimtime="00:03:22.03" />
                    <SPLIT distance="350" swimtime="00:03:59.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="429" swimtime="00:18:42.69" resultid="2834" heatid="3585" lane="4" entrytime="00:18:40.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.36" />
                    <SPLIT distance="100" swimtime="00:01:03.78" />
                    <SPLIT distance="150" swimtime="00:01:38.64" />
                    <SPLIT distance="200" swimtime="00:02:13.96" />
                    <SPLIT distance="250" swimtime="00:02:49.56" />
                    <SPLIT distance="300" swimtime="00:03:25.36" />
                    <SPLIT distance="350" swimtime="00:04:01.68" />
                    <SPLIT distance="400" swimtime="00:04:38.09" />
                    <SPLIT distance="450" swimtime="00:05:14.76" />
                    <SPLIT distance="500" swimtime="00:05:52.18" />
                    <SPLIT distance="550" swimtime="00:06:29.37" />
                    <SPLIT distance="600" swimtime="00:07:06.58" />
                    <SPLIT distance="650" swimtime="00:07:43.37" />
                    <SPLIT distance="700" swimtime="00:08:20.14" />
                    <SPLIT distance="750" swimtime="00:08:57.11" />
                    <SPLIT distance="800" swimtime="00:09:34.68" />
                    <SPLIT distance="850" swimtime="00:10:12.69" />
                    <SPLIT distance="900" swimtime="00:10:50.59" />
                    <SPLIT distance="950" swimtime="00:11:28.84" />
                    <SPLIT distance="1000" swimtime="00:12:07.18" />
                    <SPLIT distance="1050" swimtime="00:12:45.93" />
                    <SPLIT distance="1100" swimtime="00:13:25.22" />
                    <SPLIT distance="1150" swimtime="00:14:04.76" />
                    <SPLIT distance="1200" swimtime="00:14:45.63" />
                    <SPLIT distance="1250" swimtime="00:15:26.49" />
                    <SPLIT distance="1300" swimtime="00:16:06.98" />
                    <SPLIT distance="1350" swimtime="00:16:46.63" />
                    <SPLIT distance="1400" swimtime="00:17:26.57" />
                    <SPLIT distance="1450" swimtime="00:18:05.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Fernanda Pinto" birthdate="2004-09-17" gender="F" nation="BRA" license="391144" swrid="5600157" athleteid="2939" externalid="391144">
              <RESULTS>
                <RESULT eventid="1208" points="312" swimtime="00:00:33.80" resultid="2940" heatid="3536" lane="8" entrytime="00:00:36.68" entrycourse="SCM" />
                <RESULT eventid="1176" points="225" swimtime="00:00:40.07" resultid="2941" heatid="3515" lane="4" />
                <RESULT eventid="1272" points="215" reactiontime="+74" swimtime="00:00:42.10" resultid="2942" heatid="3587" lane="6" entrytime="00:00:52.73" entrycourse="SCM" />
                <RESULT eventid="1240" points="286" swimtime="00:01:16.25" resultid="2943" heatid="3565" lane="3" entrytime="00:01:21.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Felipe Kuhn" birthdate="2014-03-22" gender="M" nation="BRA" license="392121" swrid="5602536" athleteid="2961" externalid="392121">
              <RESULTS>
                <RESULT eventid="1095" points="99" swimtime="00:01:36.80" resultid="2962" heatid="3442" lane="7" entrytime="00:01:41.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="89" swimtime="00:00:55.85" resultid="2963" heatid="3404" lane="6" entrytime="00:00:59.07" entrycourse="SCM" />
                <RESULT eventid="1111" status="SICK" swimtime="00:00:00.00" resultid="2964" heatid="3456" lane="4" />
                <RESULT eventid="1131" status="SICK" swimtime="00:00:00.00" resultid="2965" heatid="3473" lane="6" entrytime="00:00:44.35" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benito" lastname="Alves Sant&apos;Ana" birthdate="2009-06-01" gender="M" nation="BRA" license="376585" swrid="5351951" athleteid="2846" externalid="376585">
              <RESULTS>
                <RESULT eventid="1200" reactiontime="+71" status="DSQ" swimtime="00:01:11.74" resultid="2847" heatid="3531" lane="3" entrytime="00:01:10.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="473" swimtime="00:04:32.23" resultid="2848" heatid="3501" lane="8" entrytime="00:04:46.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                    <SPLIT distance="100" swimtime="00:01:03.02" />
                    <SPLIT distance="150" swimtime="00:01:36.68" />
                    <SPLIT distance="200" swimtime="00:02:12.00" />
                    <SPLIT distance="250" swimtime="00:02:46.32" />
                    <SPLIT distance="300" swimtime="00:03:18.86" />
                    <SPLIT distance="350" swimtime="00:03:57.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="406" swimtime="00:02:28.04" resultid="2849" heatid="3561" lane="8" entrytime="00:02:29.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:01:10.22" />
                    <SPLIT distance="150" swimtime="00:01:55.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="310" swimtime="00:01:10.55" resultid="2850" heatid="3601" lane="7" entrytime="00:01:10.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="520" swimtime="00:17:32.83" resultid="2851" heatid="3583" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                    <SPLIT distance="100" swimtime="00:01:04.80" />
                    <SPLIT distance="150" swimtime="00:01:39.59" />
                    <SPLIT distance="200" swimtime="00:02:14.29" />
                    <SPLIT distance="250" swimtime="00:02:48.74" />
                    <SPLIT distance="300" swimtime="00:03:23.68" />
                    <SPLIT distance="350" swimtime="00:03:58.81" />
                    <SPLIT distance="400" swimtime="00:04:35.43" />
                    <SPLIT distance="450" swimtime="00:05:10.12" />
                    <SPLIT distance="500" swimtime="00:05:45.05" />
                    <SPLIT distance="550" swimtime="00:06:21.23" />
                    <SPLIT distance="600" swimtime="00:06:55.50" />
                    <SPLIT distance="650" swimtime="00:07:32.50" />
                    <SPLIT distance="700" swimtime="00:08:07.00" />
                    <SPLIT distance="750" swimtime="00:08:40.80" />
                    <SPLIT distance="800" swimtime="00:09:17.03" />
                    <SPLIT distance="850" swimtime="00:09:51.88" />
                    <SPLIT distance="900" swimtime="00:10:28.35" />
                    <SPLIT distance="950" swimtime="00:11:04.04" />
                    <SPLIT distance="1000" swimtime="00:11:39.62" />
                    <SPLIT distance="1050" swimtime="00:12:15.60" />
                    <SPLIT distance="1100" swimtime="00:12:50.80" />
                    <SPLIT distance="1150" swimtime="00:13:27.12" />
                    <SPLIT distance="1200" swimtime="00:14:03.45" />
                    <SPLIT distance="1250" swimtime="00:14:38.35" />
                    <SPLIT distance="1300" swimtime="00:15:13.62" />
                    <SPLIT distance="1350" swimtime="00:15:50.24" />
                    <SPLIT distance="1400" swimtime="00:16:25.67" />
                    <SPLIT distance="1450" swimtime="00:17:00.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Bilecki" birthdate="2007-05-28" gender="M" nation="BRA" license="406726" athleteid="3040" externalid="406726">
              <RESULTS>
                <RESULT eventid="1184" points="282" swimtime="00:00:33.15" resultid="3041" heatid="3518" lane="8" />
                <RESULT eventid="1216" points="311" swimtime="00:00:29.75" resultid="3042" heatid="3541" lane="1" />
                <RESULT eventid="1296" points="222" swimtime="00:01:18.82" resultid="3043" heatid="3598" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="306" swimtime="00:01:06.54" resultid="3044" heatid="3573" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Geovana" lastname="Dos Santos" birthdate="2011-01-20" gender="F" nation="BRA" license="367254" swrid="5602533" athleteid="2867" externalid="367254">
              <RESULTS>
                <RESULT eventid="1144" points="283" swimtime="00:05:52.17" resultid="2868" heatid="3491" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                    <SPLIT distance="100" swimtime="00:01:19.68" />
                    <SPLIT distance="150" swimtime="00:02:04.68" />
                    <SPLIT distance="200" swimtime="00:02:49.63" />
                    <SPLIT distance="250" swimtime="00:03:36.08" />
                    <SPLIT distance="300" swimtime="00:04:21.75" />
                    <SPLIT distance="350" swimtime="00:05:07.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="302" swimtime="00:00:34.14" resultid="2869" heatid="3536" lane="2" entrytime="00:00:35.09" entrycourse="SCM" />
                <RESULT eventid="1272" points="264" reactiontime="+52" swimtime="00:00:39.33" resultid="2870" heatid="3588" lane="6" entrytime="00:00:39.76" entrycourse="SCM" />
                <RESULT eventid="1240" points="281" swimtime="00:01:16.67" resultid="2871" heatid="3565" lane="4" entrytime="00:01:20.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Henrique Opuchkevich" birthdate="2011-02-22" gender="M" nation="BRA" license="406720" athleteid="3011" externalid="406720">
              <RESULTS>
                <RESULT eventid="1168" points="181" swimtime="00:01:37.60" resultid="3012" heatid="3509" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="185" swimtime="00:00:35.36" resultid="3013" heatid="3544" lane="8" />
                <RESULT eventid="1312" points="172" swimtime="00:00:44.83" resultid="3014" heatid="3609" lane="7" />
                <RESULT eventid="1248" points="199" swimtime="00:01:16.75" resultid="3015" heatid="3572" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Luiza Rimbano De Jesus" birthdate="2008-09-02" gender="F" nation="BRA" license="366819" swrid="5653297" athleteid="2976" externalid="366819">
              <RESULTS>
                <RESULT eventid="1144" points="370" swimtime="00:05:22.16" resultid="2977" heatid="3490" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.73" />
                    <SPLIT distance="100" swimtime="00:01:11.60" />
                    <SPLIT distance="150" swimtime="00:01:51.06" />
                    <SPLIT distance="200" swimtime="00:02:31.40" />
                    <SPLIT distance="250" swimtime="00:03:12.70" />
                    <SPLIT distance="300" swimtime="00:03:56.16" />
                    <SPLIT distance="350" swimtime="00:04:40.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="486" swimtime="00:00:29.16" resultid="2978" heatid="3539" lane="6" entrytime="00:00:29.71" entrycourse="SCM" />
                <RESULT eventid="1160" points="379" swimtime="00:01:26.10" resultid="2979" heatid="3504" lane="5" entrytime="00:01:32.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="328" swimtime="00:01:18.36" resultid="2980" heatid="3595" lane="5" entrytime="00:01:23.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="470" swimtime="00:01:04.61" resultid="2981" heatid="3570" lane="1" entrytime="00:01:04.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Seiffert Mafra" birthdate="2013-01-11" gender="F" nation="BRA" license="406729" athleteid="3054" externalid="406729">
              <RESULTS>
                <RESULT eventid="1086" points="102" swimtime="00:03:55.41" resultid="3055" heatid="3425" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.67" />
                    <SPLIT distance="100" swimtime="00:01:49.50" />
                    <SPLIT distance="150" swimtime="00:02:53.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="67" reactiontime="+132" swimtime="00:01:02.16" resultid="3056" heatid="3405" lane="4" />
                <RESULT eventid="1102" points="105" swimtime="00:01:59.45" resultid="3057" heatid="3444" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="129" swimtime="00:00:45.35" resultid="3058" heatid="3477" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Fernanda De Lima" birthdate="2013-09-26" gender="F" nation="BRA" license="378290" swrid="5588693" athleteid="2901" externalid="378290">
              <RESULTS>
                <RESULT eventid="1086" points="143" swimtime="00:03:30.53" resultid="2902" heatid="3424" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.02" />
                    <SPLIT distance="100" swimtime="00:01:41.73" />
                    <SPLIT distance="150" swimtime="00:02:36.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="141" reactiontime="+68" swimtime="00:00:48.51" resultid="2903" heatid="3409" lane="7" entrytime="00:00:47.67" entrycourse="SCM" />
                <RESULT eventid="1138" points="182" swimtime="00:00:40.42" resultid="2904" heatid="3479" lane="2" entrytime="00:00:43.15" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauren" lastname="Dziura" birthdate="2010-01-11" gender="F" nation="BRA" license="369416" swrid="5588668" athleteid="2891" externalid="369416">
              <RESULTS>
                <RESULT eventid="1144" points="371" swimtime="00:05:21.79" resultid="2892" heatid="3490" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.59" />
                    <SPLIT distance="100" swimtime="00:01:15.11" />
                    <SPLIT distance="150" swimtime="00:01:56.10" />
                    <SPLIT distance="200" swimtime="00:02:37.72" />
                    <SPLIT distance="250" swimtime="00:03:17.89" />
                    <SPLIT distance="300" swimtime="00:04:00.05" />
                    <SPLIT distance="350" swimtime="00:04:41.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="271" reactiontime="+67" swimtime="00:01:24.77" resultid="2893" heatid="3525" lane="2" entrytime="00:01:25.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="323" swimtime="00:02:57.50" resultid="2894" heatid="3554" lane="1" entrytime="00:03:06.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                    <SPLIT distance="100" swimtime="00:01:26.14" />
                    <SPLIT distance="150" swimtime="00:02:19.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="258" swimtime="00:01:24.82" resultid="2895" heatid="3595" lane="2" entrytime="00:01:34.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Marcos Pinto" birthdate="2006-01-26" gender="M" nation="BRA" license="391143" swrid="5600209" athleteid="2934" externalid="391143">
              <RESULTS>
                <RESULT eventid="1168" points="178" swimtime="00:01:38.13" resultid="2935" heatid="3508" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="235" swimtime="00:05:43.49" resultid="2936" heatid="3498" lane="1" entrytime="00:06:04.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                    <SPLIT distance="100" swimtime="00:01:19.71" />
                    <SPLIT distance="150" swimtime="00:02:02.90" />
                    <SPLIT distance="200" swimtime="00:02:45.44" />
                    <SPLIT distance="250" swimtime="00:03:28.63" />
                    <SPLIT distance="300" swimtime="00:04:12.81" />
                    <SPLIT distance="350" swimtime="00:04:57.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="191" swimtime="00:03:10.20" resultid="2937" heatid="3558" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.73" />
                    <SPLIT distance="100" swimtime="00:01:33.62" />
                    <SPLIT distance="150" swimtime="00:02:27.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="260" swimtime="00:01:10.18" resultid="2938" heatid="3576" lane="8" entrytime="00:01:14.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Barros Zagonel" birthdate="2006-06-01" gender="M" nation="BRA" license="347856" swrid="5622261" athleteid="2827" externalid="347856" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1168" points="318" swimtime="00:01:20.98" resultid="2828" heatid="3511" lane="8" entrytime="00:01:26.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="373" swimtime="00:00:27.99" resultid="2829" heatid="3542" lane="1" />
                <RESULT eventid="1312" points="358" swimtime="00:00:35.13" resultid="2830" heatid="3611" lane="6" entrytime="00:00:36.01" entrycourse="SCM" />
                <RESULT eventid="1248" points="344" swimtime="00:01:03.98" resultid="2831" heatid="3573" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="De Mello Araujo" birthdate="2012-08-14" gender="M" nation="BRA" license="406727" athleteid="3045" externalid="406727">
              <RESULTS>
                <RESULT eventid="1105" status="DSQ" swimtime="00:01:38.37" resultid="3046" heatid="3449" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" status="DSQ" swimtime="00:00:36.95" resultid="3047" heatid="3483" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Tomaz Zmievski" birthdate="2012-09-20" gender="F" nation="BRA" license="406725" athleteid="3035" externalid="406725">
              <RESULTS>
                <RESULT eventid="1086" points="163" swimtime="00:03:21.88" resultid="3036" heatid="3424" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.29" />
                    <SPLIT distance="100" swimtime="00:01:34.04" />
                    <SPLIT distance="150" swimtime="00:02:29.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="110" reactiontime="+95" swimtime="00:00:52.62" resultid="3037" heatid="3406" lane="4" />
                <RESULT eventid="1102" points="123" swimtime="00:01:53.54" resultid="3038" heatid="3443" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="195" swimtime="00:00:39.51" resultid="3039" heatid="3476" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Gabriel Sarmento Buski" birthdate="2010-04-05" gender="M" nation="BRA" license="399533" athleteid="2852" externalid="399533">
              <RESULTS>
                <RESULT eventid="1168" points="227" swimtime="00:01:30.62" resultid="2853" heatid="3507" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" status="DSQ" swimtime="00:05:20.30" resultid="2854" heatid="3496" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.47" />
                    <SPLIT distance="100" swimtime="00:01:13.24" />
                    <SPLIT distance="150" swimtime="00:01:54.27" />
                    <SPLIT distance="200" swimtime="00:02:35.92" />
                    <SPLIT distance="250" swimtime="00:03:18.89" />
                    <SPLIT distance="300" swimtime="00:04:00.09" />
                    <SPLIT distance="350" swimtime="00:04:42.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" status="DSQ" swimtime="00:00:41.33" resultid="2855" heatid="3608" lane="4" />
                <RESULT eventid="1264" points="304" swimtime="00:20:59.22" resultid="2856" heatid="3585" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:15.44" />
                    <SPLIT distance="150" swimtime="00:01:57.06" />
                    <SPLIT distance="200" swimtime="00:02:39.36" />
                    <SPLIT distance="250" swimtime="00:03:21.58" />
                    <SPLIT distance="300" swimtime="00:04:03.10" />
                    <SPLIT distance="350" swimtime="00:04:44.91" />
                    <SPLIT distance="400" swimtime="00:05:26.89" />
                    <SPLIT distance="450" swimtime="00:06:08.83" />
                    <SPLIT distance="500" swimtime="00:06:51.00" />
                    <SPLIT distance="550" swimtime="00:07:34.24" />
                    <SPLIT distance="600" swimtime="00:08:16.67" />
                    <SPLIT distance="650" swimtime="00:08:58.57" />
                    <SPLIT distance="700" swimtime="00:09:41.53" />
                    <SPLIT distance="750" swimtime="00:10:24.37" />
                    <SPLIT distance="800" swimtime="00:11:07.35" />
                    <SPLIT distance="850" swimtime="00:11:50.56" />
                    <SPLIT distance="900" swimtime="00:12:33.08" />
                    <SPLIT distance="950" swimtime="00:13:16.66" />
                    <SPLIT distance="1000" swimtime="00:13:59.49" />
                    <SPLIT distance="1050" swimtime="00:14:41.77" />
                    <SPLIT distance="1100" swimtime="00:15:24.18" />
                    <SPLIT distance="1150" swimtime="00:16:06.58" />
                    <SPLIT distance="1200" swimtime="00:16:48.96" />
                    <SPLIT distance="1250" swimtime="00:17:31.97" />
                    <SPLIT distance="1300" swimtime="00:18:13.73" />
                    <SPLIT distance="1350" swimtime="00:18:56.38" />
                    <SPLIT distance="1400" swimtime="00:19:39.06" />
                    <SPLIT distance="1450" swimtime="00:20:21.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaylane" lastname="Marques Ferreira" birthdate="2010-03-06" gender="F" nation="BRA" license="391146" swrid="5600211" athleteid="2950" externalid="391146">
              <RESULTS>
                <RESULT eventid="1144" points="148" swimtime="00:07:16.53" resultid="2951" heatid="3491" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.11" />
                    <SPLIT distance="100" swimtime="00:01:38.45" />
                    <SPLIT distance="150" swimtime="00:02:33.63" />
                    <SPLIT distance="200" swimtime="00:03:29.82" />
                    <SPLIT distance="250" swimtime="00:04:27.61" />
                    <SPLIT distance="300" swimtime="00:05:25.43" />
                    <SPLIT distance="350" swimtime="00:06:22.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="240" swimtime="00:00:36.87" resultid="2952" heatid="3535" lane="2" entrytime="00:00:39.69" entrycourse="SCM" />
                <RESULT eventid="1176" points="242" swimtime="00:00:39.07" resultid="2953" heatid="3516" lane="7" entrytime="00:00:46.49" entrycourse="SCM" />
                <RESULT eventid="1288" points="165" swimtime="00:01:38.41" resultid="2954" heatid="3594" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="222" swimtime="00:01:22.89" resultid="2955" heatid="3564" lane="5" entrytime="00:01:36.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thiago" lastname="Kozera Chiarato" birthdate="2008-01-22" gender="M" nation="BRA" license="406728" athleteid="3048" externalid="406728">
              <RESULTS>
                <RESULT eventid="1184" points="307" swimtime="00:00:32.24" resultid="3049" heatid="3518" lane="4" />
                <RESULT eventid="1216" points="326" swimtime="00:00:29.27" resultid="3050" heatid="3541" lane="3" />
                <RESULT eventid="1312" points="265" swimtime="00:00:38.80" resultid="3051" heatid="3609" lane="5" />
                <RESULT eventid="1296" points="244" swimtime="00:01:16.38" resultid="3052" heatid="3600" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="301" swimtime="00:01:06.88" resultid="3053" heatid="3571" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="De Mello Araujo" birthdate="2010-11-03" gender="F" nation="BRA" license="406723" athleteid="3027" externalid="406723">
              <RESULTS>
                <RESULT eventid="1192" points="152" reactiontime="+74" swimtime="00:01:42.63" resultid="3028" heatid="3524" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1160" points="195" swimtime="00:01:47.52" resultid="3029" heatid="3503" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Lara" birthdate="2014-09-02" gender="F" nation="BRA" license="406686" athleteid="2994" externalid="406686">
              <RESULTS>
                <RESULT eventid="1128" points="49" swimtime="00:01:02.32" resultid="2995" heatid="3466" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kedny" lastname="Correa" birthdate="2004-11-05" gender="M" nation="BRA" license="383858" swrid="5600142" athleteid="2905" externalid="383858">
              <RESULTS>
                <RESULT eventid="1184" points="396" swimtime="00:00:29.60" resultid="2906" heatid="3521" lane="5" entrytime="00:00:30.38" entrycourse="SCM" />
                <RESULT eventid="1152" points="466" swimtime="00:04:33.69" resultid="2907" heatid="3501" lane="1" entrytime="00:04:43.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.76" />
                    <SPLIT distance="100" swimtime="00:01:04.47" />
                    <SPLIT distance="150" swimtime="00:01:37.98" />
                    <SPLIT distance="200" swimtime="00:02:12.48" />
                    <SPLIT distance="250" swimtime="00:02:47.56" />
                    <SPLIT distance="300" swimtime="00:03:23.32" />
                    <SPLIT distance="350" swimtime="00:03:59.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="429" swimtime="00:00:26.73" resultid="2908" heatid="3542" lane="6" />
                <RESULT eventid="1296" points="295" swimtime="00:01:11.73" resultid="2909" heatid="3601" lane="2" entrytime="00:01:10.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="453" swimtime="00:18:21.89" resultid="2910" heatid="3585" lane="5" entrytime="00:19:07.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.18" />
                    <SPLIT distance="100" swimtime="00:01:04.43" />
                    <SPLIT distance="150" swimtime="00:01:39.08" />
                    <SPLIT distance="200" swimtime="00:02:14.10" />
                    <SPLIT distance="250" swimtime="00:02:49.46" />
                    <SPLIT distance="300" swimtime="00:03:25.21" />
                    <SPLIT distance="350" swimtime="00:04:01.35" />
                    <SPLIT distance="400" swimtime="00:04:38.01" />
                    <SPLIT distance="450" swimtime="00:05:14.59" />
                    <SPLIT distance="500" swimtime="00:05:51.92" />
                    <SPLIT distance="550" swimtime="00:06:29.23" />
                    <SPLIT distance="600" swimtime="00:07:06.72" />
                    <SPLIT distance="650" swimtime="00:07:44.02" />
                    <SPLIT distance="700" swimtime="00:08:21.46" />
                    <SPLIT distance="750" swimtime="00:08:59.28" />
                    <SPLIT distance="800" swimtime="00:09:37.25" />
                    <SPLIT distance="850" swimtime="00:10:15.26" />
                    <SPLIT distance="900" swimtime="00:10:53.08" />
                    <SPLIT distance="950" swimtime="00:11:31.28" />
                    <SPLIT distance="1000" swimtime="00:12:08.67" />
                    <SPLIT distance="1050" swimtime="00:12:46.37" />
                    <SPLIT distance="1100" swimtime="00:13:24.29" />
                    <SPLIT distance="1150" swimtime="00:14:02.45" />
                    <SPLIT distance="1200" swimtime="00:14:39.88" />
                    <SPLIT distance="1250" swimtime="00:15:17.26" />
                    <SPLIT distance="1300" swimtime="00:15:54.76" />
                    <SPLIT distance="1350" swimtime="00:16:32.45" />
                    <SPLIT distance="1400" swimtime="00:17:10.32" />
                    <SPLIT distance="1450" swimtime="00:17:47.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monike" lastname="Lemos Carvalho" birthdate="2008-03-28" gender="F" nation="BRA" license="307796" swrid="5600199" athleteid="2911" externalid="307796">
              <RESULTS>
                <RESULT eventid="1192" points="352" reactiontime="+72" swimtime="00:01:17.73" resultid="2912" heatid="3526" lane="6" entrytime="00:01:19.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="327" swimtime="00:00:41.14" resultid="2913" heatid="3603" lane="4" />
                <RESULT eventid="1240" points="406" swimtime="00:01:07.84" resultid="2914" heatid="3567" lane="4" entrytime="00:01:10.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Mingorance Martins" birthdate="2007-10-13" gender="M" nation="BRA" license="393920" swrid="5622295" athleteid="2971" externalid="393920">
              <RESULTS>
                <RESULT eventid="1152" points="442" swimtime="00:04:38.57" resultid="2972" heatid="3495" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:05.86" />
                    <SPLIT distance="150" swimtime="00:01:41.66" />
                    <SPLIT distance="200" swimtime="00:02:17.86" />
                    <SPLIT distance="250" swimtime="00:02:53.12" />
                    <SPLIT distance="300" swimtime="00:03:28.68" />
                    <SPLIT distance="350" swimtime="00:04:04.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="482" swimtime="00:00:25.71" resultid="2973" heatid="3549" lane="3" entrytime="00:00:26.03" entrycourse="SCM" />
                <RESULT eventid="1264" points="385" swimtime="00:19:24.04" resultid="2974" heatid="3583" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                    <SPLIT distance="100" swimtime="00:01:14.20" />
                    <SPLIT distance="150" swimtime="00:01:53.89" />
                    <SPLIT distance="200" swimtime="00:02:34.00" />
                    <SPLIT distance="250" swimtime="00:03:14.46" />
                    <SPLIT distance="300" swimtime="00:03:54.00" />
                    <SPLIT distance="350" swimtime="00:04:33.91" />
                    <SPLIT distance="400" swimtime="00:05:13.96" />
                    <SPLIT distance="450" swimtime="00:05:54.12" />
                    <SPLIT distance="500" swimtime="00:06:34.67" />
                    <SPLIT distance="550" swimtime="00:07:15.72" />
                    <SPLIT distance="600" swimtime="00:07:56.00" />
                    <SPLIT distance="650" swimtime="00:08:35.68" />
                    <SPLIT distance="700" swimtime="00:09:14.97" />
                    <SPLIT distance="750" swimtime="00:09:54.28" />
                    <SPLIT distance="800" swimtime="00:10:32.90" />
                    <SPLIT distance="850" swimtime="00:11:11.81" />
                    <SPLIT distance="900" swimtime="00:11:49.76" />
                    <SPLIT distance="950" swimtime="00:12:28.75" />
                    <SPLIT distance="1000" swimtime="00:13:08.18" />
                    <SPLIT distance="1050" swimtime="00:13:46.82" />
                    <SPLIT distance="1100" swimtime="00:14:25.24" />
                    <SPLIT distance="1150" swimtime="00:15:03.01" />
                    <SPLIT distance="1200" swimtime="00:15:40.34" />
                    <SPLIT distance="1250" swimtime="00:16:17.93" />
                    <SPLIT distance="1300" swimtime="00:16:55.65" />
                    <SPLIT distance="1350" swimtime="00:17:33.74" />
                    <SPLIT distance="1400" swimtime="00:18:12.27" />
                    <SPLIT distance="1450" swimtime="00:18:48.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="492" swimtime="00:00:56.77" resultid="2975" heatid="3580" lane="1" entrytime="00:00:57.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Vitor Navarro Zanini" birthdate="2008-06-30" gender="M" nation="BRA" license="369415" swrid="5600273" athleteid="2886" externalid="369415">
              <RESULTS>
                <RESULT eventid="1168" points="333" swimtime="00:01:19.68" resultid="2887" heatid="3510" lane="6" entrytime="00:01:30.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="326" swimtime="00:05:08.22" resultid="2888" heatid="3498" lane="6" entrytime="00:05:46.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.25" />
                    <SPLIT distance="100" swimtime="00:01:13.98" />
                    <SPLIT distance="150" swimtime="00:01:54.40" />
                    <SPLIT distance="200" swimtime="00:02:34.12" />
                    <SPLIT distance="250" swimtime="00:03:13.28" />
                    <SPLIT distance="300" swimtime="00:03:51.92" />
                    <SPLIT distance="350" swimtime="00:04:30.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="304" swimtime="00:02:43.02" resultid="2889" heatid="3558" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:20.58" />
                    <SPLIT distance="150" swimtime="00:02:07.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="350" swimtime="00:00:35.40" resultid="2890" heatid="3610" lane="3" entrytime="00:00:41.98" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Rodrigues Galvao" birthdate="2007-04-19" gender="M" nation="BRA" license="376586" swrid="5600247" athleteid="2841" externalid="376586">
              <RESULTS>
                <RESULT eventid="1184" points="519" swimtime="00:00:27.06" resultid="2842" heatid="3521" lane="4" entrytime="00:00:29.79" entrycourse="SCM" />
                <RESULT eventid="1216" points="495" swimtime="00:00:25.48" resultid="2843" heatid="3549" lane="2" entrytime="00:00:26.35" entrycourse="SCM" />
                <RESULT eventid="1296" points="450" swimtime="00:01:02.31" resultid="2844" heatid="3602" lane="8" entrytime="00:01:03.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="493" swimtime="00:00:56.76" resultid="2845" heatid="3580" lane="8" entrytime="00:00:58.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcus" lastname="Vinicius De Almeida" birthdate="2009-06-16" gender="M" nation="BRA" license="348099" swrid="5600272" athleteid="2861" externalid="348099">
              <RESULTS>
                <RESULT eventid="1200" points="395" reactiontime="+72" swimtime="00:01:05.84" resultid="2862" heatid="3531" lane="4" entrytime="00:01:08.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="453" swimtime="00:01:11.94" resultid="2863" heatid="3512" lane="7" entrytime="00:01:18.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="457" swimtime="00:00:32.37" resultid="2864" heatid="3608" lane="6" />
                <RESULT eventid="1280" points="398" reactiontime="+55" swimtime="00:00:30.05" resultid="2865" heatid="3593" lane="1" entrytime="00:00:32.23" entrycourse="SCM" />
                <RESULT eventid="1264" points="474" swimtime="00:18:05.90" resultid="2866" heatid="3583" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                    <SPLIT distance="100" swimtime="00:01:05.63" />
                    <SPLIT distance="150" swimtime="00:01:40.16" />
                    <SPLIT distance="200" swimtime="00:02:15.50" />
                    <SPLIT distance="250" swimtime="00:02:50.40" />
                    <SPLIT distance="300" swimtime="00:03:25.53" />
                    <SPLIT distance="350" swimtime="00:04:00.74" />
                    <SPLIT distance="400" swimtime="00:04:36.72" />
                    <SPLIT distance="450" swimtime="00:05:12.63" />
                    <SPLIT distance="500" swimtime="00:05:49.01" />
                    <SPLIT distance="550" swimtime="00:06:25.78" />
                    <SPLIT distance="600" swimtime="00:07:02.03" />
                    <SPLIT distance="650" swimtime="00:07:38.95" />
                    <SPLIT distance="700" swimtime="00:08:15.68" />
                    <SPLIT distance="750" swimtime="00:08:52.81" />
                    <SPLIT distance="800" swimtime="00:09:30.26" />
                    <SPLIT distance="850" swimtime="00:10:07.34" />
                    <SPLIT distance="900" swimtime="00:10:44.31" />
                    <SPLIT distance="950" swimtime="00:11:21.17" />
                    <SPLIT distance="1000" swimtime="00:11:58.09" />
                    <SPLIT distance="1050" swimtime="00:12:34.20" />
                    <SPLIT distance="1100" swimtime="00:13:11.40" />
                    <SPLIT distance="1150" swimtime="00:13:48.49" />
                    <SPLIT distance="1200" swimtime="00:14:25.69" />
                    <SPLIT distance="1250" swimtime="00:15:02.80" />
                    <SPLIT distance="1300" swimtime="00:15:39.67" />
                    <SPLIT distance="1350" swimtime="00:16:16.34" />
                    <SPLIT distance="1400" swimtime="00:16:53.28" />
                    <SPLIT distance="1450" swimtime="00:17:30.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Melo" birthdate="2015-02-07" gender="F" nation="BRA" license="406717" athleteid="2996" externalid="406717">
              <RESULTS>
                <RESULT eventid="1092" points="112" swimtime="00:01:44.05" resultid="2997" heatid="3437" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="125" swimtime="00:00:50.49" resultid="2998" heatid="3418" lane="6" />
                <RESULT eventid="1108" points="62" swimtime="00:01:01.54" resultid="2999" heatid="3452" lane="2" />
                <RESULT eventid="1128" points="132" swimtime="00:00:44.97" resultid="3000" heatid="3466" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1007" nation="BRA" region="PR" clubid="3059" swrid="93785" name="Santa Mônica Clube De Campo" shortname="Santa Mônica">
          <ATHLETES>
            <ATHLETE firstname="Mathias" lastname="Lopes Batista" birthdate="2012-08-22" gender="M" nation="BRA" license="399740" swrid="5652889" athleteid="3312" externalid="399740">
              <RESULTS>
                <RESULT eventid="1077" points="121" reactiontime="+82" swimtime="00:00:44.59" resultid="3313" heatid="3414" lane="1" entrytime="00:00:47.50" entrycourse="SCM" />
                <RESULT eventid="1141" points="129" swimtime="00:00:39.80" resultid="3314" heatid="3485" lane="8" entrytime="00:00:38.92" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Luiz Cruz" birthdate="2012-10-13" gender="M" nation="BRA" license="393209" swrid="5616447" athleteid="3289" externalid="393209">
              <RESULTS>
                <RESULT eventid="1089" points="159" swimtime="00:03:03.37" resultid="3290" heatid="3431" lane="5" entrytime="00:03:14.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.49" />
                    <SPLIT distance="100" swimtime="00:01:28.56" />
                    <SPLIT distance="150" swimtime="00:02:16.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="88" swimtime="00:02:04.23" resultid="3291" heatid="3396" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" status="DSQ" swimtime="00:01:52.43" resultid="3292" heatid="3464" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="150" swimtime="00:00:37.89" resultid="3293" heatid="3484" lane="6" entrytime="00:00:41.31" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Cavassin Ieger" birthdate="2011-08-31" gender="M" nation="BRA" license="367149" swrid="5588743" athleteid="3138" externalid="367149">
              <RESULTS>
                <RESULT eventid="1168" points="236" swimtime="00:01:29.42" resultid="3139" heatid="3510" lane="7" entrytime="00:01:34.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="290" swimtime="00:05:20.64" resultid="3140" heatid="3496" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                    <SPLIT distance="100" swimtime="00:01:14.36" />
                    <SPLIT distance="150" swimtime="00:01:56.08" />
                    <SPLIT distance="200" swimtime="00:02:37.22" />
                    <SPLIT distance="250" swimtime="00:03:19.36" />
                    <SPLIT distance="300" swimtime="00:04:00.63" />
                    <SPLIT distance="350" swimtime="00:04:42.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="232" swimtime="00:00:40.56" resultid="3141" heatid="3610" lane="6" entrytime="00:00:43.58" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Leticia Durat" birthdate="2008-02-09" gender="F" nation="BRA" license="331636" swrid="5600200" athleteid="3082" externalid="331636">
              <RESULTS>
                <RESULT eventid="1208" points="409" swimtime="00:00:30.89" resultid="3083" heatid="3538" lane="5" entrytime="00:00:30.38" entrycourse="SCM" />
                <RESULT eventid="1160" status="DSQ" swimtime="00:01:29.66" resultid="3084" heatid="3505" lane="6" entrytime="00:01:26.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="402" swimtime="00:01:08.07" resultid="3085" heatid="3563" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Giuseppe Bulla Lanaro" birthdate="2007-05-22" gender="M" nation="BRA" license="331630" swrid="5600174" athleteid="3069" externalid="331630">
              <RESULTS>
                <RESULT eventid="1152" points="601" swimtime="00:04:11.46" resultid="3070" heatid="3501" lane="5" entrytime="00:04:12.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.50" />
                    <SPLIT distance="100" swimtime="00:00:58.97" />
                    <SPLIT distance="150" swimtime="00:01:30.62" />
                    <SPLIT distance="200" swimtime="00:02:02.42" />
                    <SPLIT distance="250" swimtime="00:02:34.60" />
                    <SPLIT distance="300" swimtime="00:03:07.30" />
                    <SPLIT distance="350" swimtime="00:03:40.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="530" swimtime="00:00:24.91" resultid="3071" heatid="3550" lane="8" entrytime="00:00:25.49" entrycourse="SCM" />
                <RESULT eventid="1296" points="496" swimtime="00:01:00.33" resultid="3072" heatid="3602" lane="7" entrytime="00:01:02.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="584" swimtime="00:00:53.63" resultid="3073" heatid="3581" lane="7" entrytime="00:00:54.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Zanotto De Souza" birthdate="2013-08-24" gender="M" nation="BRA" license="388361" swrid="5588974" athleteid="3271" externalid="388361">
              <RESULTS>
                <RESULT eventid="1089" points="202" swimtime="00:02:49.34" resultid="3272" heatid="3432" lane="3" entrytime="00:02:58.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                    <SPLIT distance="100" swimtime="00:01:23.07" />
                    <SPLIT distance="150" swimtime="00:02:08.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="172" reactiontime="+68" swimtime="00:00:39.69" resultid="3273" heatid="3415" lane="1" entrytime="00:00:40.83" entrycourse="SCM" />
                <RESULT eventid="1105" points="150" swimtime="00:01:32.67" resultid="3274" heatid="3448" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="205" swimtime="00:00:34.18" resultid="3275" heatid="3487" lane="7" entrytime="00:00:34.41" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Borges Piekarzievicz" birthdate="2013-09-10" gender="M" nation="BRA" license="403142" swrid="5676294" athleteid="3335" externalid="403142">
              <RESULTS>
                <RESULT eventid="1077" points="51" swimtime="00:00:59.45" resultid="3336" heatid="3412" lane="3" />
                <RESULT eventid="1141" points="91" swimtime="00:00:44.74" resultid="3337" heatid="3482" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Analyce" lastname="Nunes Porto Luz" birthdate="2006-10-29" gender="F" nation="BRA" license="369322" swrid="5600226" athleteid="3074" externalid="369322">
              <RESULTS>
                <RESULT eventid="1144" points="521" swimtime="00:04:47.40" resultid="3075" heatid="3494" lane="2" entrytime="00:04:46.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:07.87" />
                    <SPLIT distance="150" swimtime="00:01:43.55" />
                    <SPLIT distance="200" swimtime="00:02:19.70" />
                    <SPLIT distance="250" swimtime="00:02:55.95" />
                    <SPLIT distance="300" swimtime="00:03:33.06" />
                    <SPLIT distance="350" swimtime="00:04:10.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="460" swimtime="00:00:31.58" resultid="3076" heatid="3516" lane="5" entrytime="00:00:32.89" entrycourse="SCM" />
                <RESULT eventid="1288" points="426" swimtime="00:01:11.78" resultid="3077" heatid="3596" lane="6" entrytime="00:01:10.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Breno" lastname="Borges Piekarzievicz" birthdate="2011-11-11" gender="M" nation="BRA" license="403144" swrid="5676295" athleteid="3341" externalid="403144">
              <RESULTS>
                <RESULT eventid="1168" status="DSQ" swimtime="00:01:49.67" resultid="3342" heatid="3507" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="122" swimtime="00:00:40.55" resultid="3343" heatid="3541" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Prestes" birthdate="2014-01-16" gender="M" nation="BRA" license="382249" swrid="5602574" athleteid="3240" externalid="382249">
              <RESULTS>
                <RESULT eventid="1095" points="117" swimtime="00:01:31.66" resultid="3241" heatid="3442" lane="2" entrytime="00:01:36.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="136" swimtime="00:00:48.48" resultid="3242" heatid="3404" lane="5" entrytime="00:00:56.12" entrycourse="SCM" />
                <RESULT eventid="1111" points="65" swimtime="00:00:54.09" resultid="3243" heatid="3458" lane="1" />
                <RESULT eventid="1131" points="136" swimtime="00:00:39.15" resultid="3244" heatid="3474" lane="2" entrytime="00:00:41.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathalia" lastname="Lourenco Osorio" birthdate="2007-04-14" gender="F" nation="BRA" license="307465" swrid="5600203" athleteid="3064" externalid="307465">
              <RESULTS>
                <RESULT eventid="1208" points="543" swimtime="00:00:28.10" resultid="3065" heatid="3534" lane="2" />
                <RESULT eventid="1192" points="524" reactiontime="+70" swimtime="00:01:08.06" resultid="3066" heatid="3527" lane="5" entrytime="00:01:09.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="463" swimtime="00:00:36.65" resultid="3067" heatid="3606" lane="6" entrytime="00:00:38.20" entrycourse="SCM" />
                <RESULT eventid="1272" points="502" reactiontime="+76" swimtime="00:00:31.77" resultid="3068" heatid="3589" lane="6" entrytime="00:00:32.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Ruschel" birthdate="2009-12-28" gender="F" nation="BRA" license="371384" swrid="5600251" athleteid="3176" externalid="371384">
              <RESULTS>
                <RESULT eventid="1256" points="398" swimtime="00:20:34.10" resultid="3177" heatid="3582" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.55" />
                    <SPLIT distance="100" swimtime="00:01:15.79" />
                    <SPLIT distance="150" swimtime="00:01:57.50" />
                    <SPLIT distance="200" swimtime="00:02:38.87" />
                    <SPLIT distance="250" swimtime="00:03:20.41" />
                    <SPLIT distance="300" swimtime="00:04:01.77" />
                    <SPLIT distance="350" swimtime="00:04:44.35" />
                    <SPLIT distance="400" swimtime="00:05:26.18" />
                    <SPLIT distance="450" swimtime="00:06:06.44" />
                    <SPLIT distance="500" swimtime="00:06:47.96" />
                    <SPLIT distance="550" swimtime="00:07:29.56" />
                    <SPLIT distance="600" swimtime="00:08:11.71" />
                    <SPLIT distance="650" swimtime="00:08:53.16" />
                    <SPLIT distance="700" swimtime="00:09:35.06" />
                    <SPLIT distance="750" swimtime="00:10:16.98" />
                    <SPLIT distance="800" swimtime="00:10:58.53" />
                    <SPLIT distance="850" swimtime="00:11:39.80" />
                    <SPLIT distance="900" swimtime="00:12:21.48" />
                    <SPLIT distance="950" swimtime="00:13:02.32" />
                    <SPLIT distance="1000" swimtime="00:13:44.20" />
                    <SPLIT distance="1050" swimtime="00:14:25.61" />
                    <SPLIT distance="1100" swimtime="00:15:07.24" />
                    <SPLIT distance="1150" swimtime="00:15:48.29" />
                    <SPLIT distance="1200" swimtime="00:16:30.11" />
                    <SPLIT distance="1250" swimtime="00:17:10.95" />
                    <SPLIT distance="1300" swimtime="00:17:52.82" />
                    <SPLIT distance="1350" swimtime="00:18:33.77" />
                    <SPLIT distance="1400" swimtime="00:19:14.49" />
                    <SPLIT distance="1450" swimtime="00:19:55.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="484" swimtime="00:01:03.96" resultid="3178" heatid="3569" lane="2" entrytime="00:01:06.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabrizio" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="M" nation="BRA" license="344303" swrid="5559846" athleteid="3091" externalid="344303">
              <RESULTS>
                <RESULT eventid="1184" points="446" swimtime="00:00:28.45" resultid="3092" heatid="3522" lane="8" entrytime="00:00:29.46" entrycourse="SCM" />
                <RESULT eventid="1216" points="404" swimtime="00:00:27.26" resultid="3093" heatid="3548" lane="2" entrytime="00:00:27.53" entrycourse="SCM" />
                <RESULT eventid="1296" points="428" swimtime="00:01:03.40" resultid="3094" heatid="3599" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="437" swimtime="00:00:59.07" resultid="3095" heatid="3579" lane="1" entrytime="00:01:00.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Celli Schneider" birthdate="2013-02-04" gender="M" nation="BRA" license="377317" swrid="5588588" athleteid="3205" externalid="377317">
              <RESULTS>
                <RESULT eventid="1077" points="150" reactiontime="+68" swimtime="00:00:41.54" resultid="3206" heatid="3414" lane="5" entrytime="00:00:41.45" entrycourse="SCM" />
                <RESULT eventid="1105" points="125" swimtime="00:01:38.32" resultid="3207" heatid="3450" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="182" swimtime="00:00:35.51" resultid="3208" heatid="3486" lane="5" entrytime="00:00:35.57" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lais" lastname="Manika Broto" birthdate="2013-03-27" gender="F" nation="BRA" license="378054" swrid="5588795" athleteid="3226" externalid="378054">
              <RESULTS>
                <RESULT eventid="1086" points="264" swimtime="00:02:51.81" resultid="3227" heatid="3426" lane="3" entrytime="00:03:06.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:01:24.19" />
                    <SPLIT distance="150" swimtime="00:02:10.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" status="DSQ" swimtime="00:00:42.73" resultid="3228" heatid="3409" lane="5" entrytime="00:00:45.24" entrycourse="SCM" />
                <RESULT eventid="1102" points="241" swimtime="00:01:30.72" resultid="3229" heatid="3447" lane="8" entrytime="00:01:49.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="278" swimtime="00:00:35.10" resultid="3230" heatid="3480" lane="7" entrytime="00:00:38.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Hugo Dos Santos" birthdate="2014-07-25" gender="M" nation="BRA" license="397420" swrid="5641766" athleteid="3307" externalid="397420">
              <RESULTS>
                <RESULT eventid="1095" points="85" swimtime="00:01:41.86" resultid="3308" heatid="3442" lane="1" entrytime="00:01:51.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="74" swimtime="00:00:52.62" resultid="3309" heatid="3423" lane="8" entrytime="00:00:58.01" entrycourse="SCM" />
                <RESULT eventid="1111" points="42" swimtime="00:01:02.13" resultid="3310" heatid="3457" lane="6" />
                <RESULT eventid="1131" points="91" swimtime="00:00:44.80" resultid="3311" heatid="3473" lane="7" entrytime="00:00:50.00" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Ieger" birthdate="2009-02-20" gender="M" nation="BRA" license="356888" swrid="5600180" athleteid="3112" externalid="356888">
              <RESULTS>
                <RESULT eventid="1168" points="391" swimtime="00:01:15.54" resultid="3113" heatid="3512" lane="2" entrytime="00:01:16.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="402" swimtime="00:00:27.30" resultid="3114" heatid="3549" lane="1" entrytime="00:00:26.62" entrycourse="SCM" />
                <RESULT eventid="1248" points="403" swimtime="00:01:00.67" resultid="3115" heatid="3579" lane="7" entrytime="00:01:00.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Fontoura Barros" birthdate="2011-08-04" gender="F" nation="BRA" license="403143" swrid="5676298" athleteid="3338" externalid="403143">
              <RESULTS>
                <RESULT eventid="1208" points="150" swimtime="00:00:43.14" resultid="3339" heatid="3533" lane="4" />
                <RESULT eventid="1160" points="144" swimtime="00:01:58.87" resultid="3340" heatid="3502" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Garcia Reschetti Rubbo" birthdate="2011-08-06" gender="F" nation="BRA" license="367053" swrid="5588720" athleteid="3126" externalid="367053" level="DCOMP IT">
              <RESULTS>
                <RESULT eventid="1144" points="257" swimtime="00:06:03.35" resultid="3127" heatid="3492" lane="3" entrytime="00:06:25.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                    <SPLIT distance="100" swimtime="00:01:23.46" />
                    <SPLIT distance="150" swimtime="00:02:10.11" />
                    <SPLIT distance="200" swimtime="00:02:56.46" />
                    <SPLIT distance="250" swimtime="00:03:43.82" />
                    <SPLIT distance="300" swimtime="00:04:31.60" />
                    <SPLIT distance="350" swimtime="00:05:19.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="266" swimtime="00:00:35.61" resultid="3128" heatid="3536" lane="6" entrytime="00:00:34.95" entrycourse="SCM" />
                <RESULT eventid="1160" points="255" swimtime="00:01:38.25" resultid="3129" heatid="3504" lane="1" entrytime="00:01:40.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cardim Martins" birthdate="2010-09-01" gender="F" nation="BRA" license="390920" swrid="5600130" athleteid="3377" externalid="390920">
              <RESULTS>
                <RESULT eventid="1144" points="281" swimtime="00:05:53.02" resultid="3378" heatid="3491" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                    <SPLIT distance="100" swimtime="00:01:22.26" />
                    <SPLIT distance="150" swimtime="00:02:06.00" />
                    <SPLIT distance="200" swimtime="00:02:50.66" />
                    <SPLIT distance="250" swimtime="00:03:35.88" />
                    <SPLIT distance="300" swimtime="00:04:21.68" />
                    <SPLIT distance="350" swimtime="00:05:08.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="218" swimtime="00:00:40.47" resultid="3379" heatid="3514" lane="6" />
                <RESULT eventid="1272" points="238" reactiontime="+61" swimtime="00:00:40.70" resultid="3380" heatid="3587" lane="5" entrytime="00:00:47.80" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Gabriel Broto" birthdate="2014-09-14" gender="M" nation="BRA" license="402171" swrid="5661345" athleteid="3332" externalid="402171">
              <RESULTS>
                <RESULT eventid="1095" points="31" swimtime="00:02:22.17" resultid="3333" heatid="3440" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:07.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="29" reactiontime="+78" swimtime="00:01:11.92" resultid="3334" heatid="3421" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Gelenski Pelaio" birthdate="2005-10-10" gender="M" nation="BRA" license="281473" swrid="5600173" athleteid="3162" externalid="281473" level="UNIDOMBOSC">
              <RESULTS>
                <RESULT eventid="1184" points="558" swimtime="00:00:26.41" resultid="3163" heatid="3522" lane="5" entrytime="00:00:26.11" entrycourse="SCM" />
                <RESULT eventid="1216" points="507" swimtime="00:00:25.27" resultid="3164" heatid="3550" lane="2" entrytime="00:00:24.52" entrycourse="SCM" />
                <RESULT eventid="1296" points="514" swimtime="00:00:59.62" resultid="3165" heatid="3602" lane="5" entrytime="00:00:58.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="544" swimtime="00:00:54.90" resultid="3166" heatid="3581" lane="1" entrytime="00:00:54.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="Cirilo Da Cunha" birthdate="2013-05-26" gender="F" nation="BRA" license="377316" swrid="5588595" athleteid="3200" externalid="377316">
              <RESULTS>
                <RESULT eventid="1062" status="DSQ" swimtime="00:02:04.23" resultid="3201" heatid="3393" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1086" points="257" swimtime="00:02:53.32" resultid="3202" heatid="3426" lane="4" entrytime="00:03:04.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.76" />
                    <SPLIT distance="100" swimtime="00:01:23.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1118" points="127" swimtime="00:01:47.52" resultid="3203" heatid="3461" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="228" swimtime="00:00:37.53" resultid="3204" heatid="3479" lane="4" entrytime="00:00:39.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Pinterich Almeida" birthdate="2005-03-13" gender="M" nation="BRA" license="330749" swrid="5600235" athleteid="3118" externalid="330749">
              <RESULTS>
                <RESULT eventid="1152" points="596" swimtime="00:04:12.15" resultid="3119" heatid="3495" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.17" />
                    <SPLIT distance="100" swimtime="00:00:59.96" />
                    <SPLIT distance="150" swimtime="00:01:31.84" />
                    <SPLIT distance="200" swimtime="00:02:04.29" />
                    <SPLIT distance="250" swimtime="00:02:36.31" />
                    <SPLIT distance="300" swimtime="00:03:08.83" />
                    <SPLIT distance="350" swimtime="00:03:41.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="520" reactiontime="+47" swimtime="00:00:27.48" resultid="3120" heatid="3593" lane="5" entrytime="00:00:27.29" entrycourse="SCM" />
                <RESULT eventid="1248" points="617" swimtime="00:00:52.67" resultid="3121" heatid="3581" lane="5" entrytime="00:00:52.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Aparecida Lourenço Alves" birthdate="2013-11-06" gender="F" nation="BRA" license="387374" swrid="5588530" athleteid="3249" externalid="387374">
              <RESULTS>
                <RESULT eventid="1074" points="124" swimtime="00:00:50.58" resultid="3250" heatid="3409" lane="8" entrytime="00:00:50.76" entrycourse="SCM" />
                <RESULT eventid="1138" points="159" swimtime="00:00:42.30" resultid="3251" heatid="3479" lane="8" entrytime="00:00:43.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emily" lastname="Sayuri Tangueria De Lima" birthdate="2010-06-11" gender="F" nation="BRA" license="367215" swrid="5588901" athleteid="3154" externalid="367215">
              <RESULTS>
                <RESULT eventid="1144" points="409" swimtime="00:05:11.40" resultid="3155" heatid="3491" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.34" />
                    <SPLIT distance="100" swimtime="00:01:14.06" />
                    <SPLIT distance="150" swimtime="00:01:53.49" />
                    <SPLIT distance="200" swimtime="00:02:33.33" />
                    <SPLIT distance="250" swimtime="00:03:14.35" />
                    <SPLIT distance="300" swimtime="00:03:54.04" />
                    <SPLIT distance="350" swimtime="00:04:32.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1176" points="368" swimtime="00:00:34.01" resultid="3156" heatid="3514" lane="4" />
                <RESULT eventid="1288" points="348" swimtime="00:01:16.82" resultid="3157" heatid="3596" lane="8" entrytime="00:01:21.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Novakoski" birthdate="2009-03-05" gender="F" nation="BRA" license="339136" swrid="5600225" athleteid="3100" externalid="339136">
              <RESULTS>
                <RESULT eventid="1208" points="419" swimtime="00:00:30.62" resultid="3101" heatid="3538" lane="7" entrytime="00:00:31.40" entrycourse="SCM" />
                <RESULT eventid="1256" points="365" swimtime="00:21:10.54" resultid="3102" heatid="3582" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                    <SPLIT distance="100" swimtime="00:01:16.72" />
                    <SPLIT distance="150" swimtime="00:01:57.66" />
                    <SPLIT distance="200" swimtime="00:02:38.97" />
                    <SPLIT distance="250" swimtime="00:03:20.57" />
                    <SPLIT distance="300" swimtime="00:04:01.81" />
                    <SPLIT distance="350" swimtime="00:04:43.77" />
                    <SPLIT distance="400" swimtime="00:05:25.44" />
                    <SPLIT distance="450" swimtime="00:06:06.99" />
                    <SPLIT distance="500" swimtime="00:06:48.49" />
                    <SPLIT distance="550" swimtime="00:07:30.19" />
                    <SPLIT distance="600" swimtime="00:08:11.80" />
                    <SPLIT distance="650" swimtime="00:08:53.38" />
                    <SPLIT distance="700" swimtime="00:09:35.90" />
                    <SPLIT distance="750" swimtime="00:10:18.69" />
                    <SPLIT distance="800" swimtime="00:11:01.51" />
                    <SPLIT distance="850" swimtime="00:11:44.94" />
                    <SPLIT distance="900" swimtime="00:12:28.62" />
                    <SPLIT distance="950" swimtime="00:13:11.63" />
                    <SPLIT distance="1000" swimtime="00:13:55.09" />
                    <SPLIT distance="1050" swimtime="00:14:39.12" />
                    <SPLIT distance="1100" swimtime="00:15:23.17" />
                    <SPLIT distance="1150" swimtime="00:16:07.89" />
                    <SPLIT distance="1200" swimtime="00:16:51.60" />
                    <SPLIT distance="1250" swimtime="00:17:34.87" />
                    <SPLIT distance="1300" swimtime="00:18:18.96" />
                    <SPLIT distance="1350" swimtime="00:19:03.05" />
                    <SPLIT distance="1400" swimtime="00:19:47.56" />
                    <SPLIT distance="1450" swimtime="00:20:31.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="434" swimtime="00:01:06.37" resultid="3103" heatid="3568" lane="5" entrytime="00:01:08.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose" lastname="Vinicius Batistella" birthdate="2012-05-15" gender="M" nation="BRA" license="403785" swrid="5684613" athleteid="3359" externalid="403785">
              <RESULTS>
                <RESULT eventid="1089" points="127" swimtime="00:03:17.23" resultid="3360" heatid="3430" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.53" />
                    <SPLIT distance="100" swimtime="00:01:32.45" />
                    <SPLIT distance="150" swimtime="00:02:25.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="151" swimtime="00:00:37.80" resultid="3361" heatid="3483" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Helena Vieira Jussen" birthdate="2011-12-29" gender="F" nation="BRA" license="372282" swrid="5588740" athleteid="3179" externalid="372282">
              <RESULTS>
                <RESULT eventid="1144" points="238" swimtime="00:06:12.99" resultid="3180" heatid="3492" lane="6" entrytime="00:06:37.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.42" />
                    <SPLIT distance="100" swimtime="00:01:24.42" />
                    <SPLIT distance="150" swimtime="00:02:13.11" />
                    <SPLIT distance="200" swimtime="00:03:01.47" />
                    <SPLIT distance="250" swimtime="00:03:50.39" />
                    <SPLIT distance="300" swimtime="00:04:39.12" />
                    <SPLIT distance="350" swimtime="00:05:27.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="264" swimtime="00:00:35.70" resultid="3181" heatid="3535" lane="4" entrytime="00:00:37.43" entrycourse="SCM" />
                <RESULT eventid="1304" points="287" swimtime="00:00:42.97" resultid="3182" heatid="3605" lane="5" entrytime="00:00:44.25" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Victoria De Medeiros Da Rocha" birthdate="2014-08-14" gender="F" nation="BRA" license="403782" swrid="5684611" athleteid="3351" externalid="403782">
              <RESULTS>
                <RESULT eventid="1080" points="55" reactiontime="+82" swimtime="00:01:06.21" resultid="3352" heatid="3417" lane="6" />
                <RESULT eventid="1068" points="52" swimtime="00:01:15.69" resultid="3353" heatid="3399" lane="6" />
                <RESULT eventid="1108" points="28" swimtime="00:01:20.19" resultid="3354" heatid="3453" lane="4" />
                <RESULT eventid="1128" points="71" swimtime="00:00:55.33" resultid="3355" heatid="3467" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Marini" birthdate="2014-04-09" gender="M" nation="BRA" license="382247" swrid="5684582" athleteid="3231" externalid="382247">
              <RESULTS>
                <RESULT eventid="1095" points="110" swimtime="00:01:33.42" resultid="3232" heatid="3439" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="82" reactiontime="+78" swimtime="00:00:50.75" resultid="3233" heatid="3421" lane="1" />
                <RESULT eventid="1111" points="56" swimtime="00:00:56.58" resultid="3234" heatid="3457" lane="8" />
                <RESULT eventid="1131" points="109" swimtime="00:00:42.17" resultid="3235" heatid="3471" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Nogueira Silva" birthdate="2011-08-13" gender="M" nation="BRA" license="367150" swrid="5588832" athleteid="3142" externalid="367150">
              <RESULTS>
                <RESULT eventid="1168" points="252" swimtime="00:01:27.46" resultid="3143" heatid="3508" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="322" swimtime="00:05:09.48" resultid="3144" heatid="3496" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.96" />
                    <SPLIT distance="100" swimtime="00:01:14.03" />
                    <SPLIT distance="150" swimtime="00:01:52.58" />
                    <SPLIT distance="200" swimtime="00:02:32.44" />
                    <SPLIT distance="250" swimtime="00:03:12.31" />
                    <SPLIT distance="300" swimtime="00:03:51.52" />
                    <SPLIT distance="350" swimtime="00:04:31.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="295" swimtime="00:00:30.27" resultid="3145" heatid="3545" lane="1" entrytime="00:00:31.71" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabio" lastname="C Burak" birthdate="2009-08-29" gender="M" nation="BRA" license="343297" swrid="5600126" athleteid="3285" externalid="343297">
              <RESULTS>
                <RESULT eventid="1200" points="421" reactiontime="+78" swimtime="00:01:04.48" resultid="3286" heatid="3531" lane="7" entrytime="00:01:13.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="440" swimtime="00:01:12.67" resultid="3287" heatid="3512" lane="6" entrytime="00:01:14.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="376" swimtime="00:00:27.91" resultid="3288" heatid="3547" lane="3" entrytime="00:00:28.20" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Strapasson" birthdate="2012-03-01" gender="M" nation="BRA" license="371377" swrid="5602585" athleteid="3167" externalid="371377">
              <RESULTS>
                <RESULT eventid="1089" points="255" swimtime="00:02:36.56" resultid="3168" heatid="3432" lane="2" entrytime="00:03:06.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.71" />
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                    <SPLIT distance="150" swimtime="00:01:56.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="244" swimtime="00:01:28.43" resultid="3169" heatid="3398" lane="5" entrytime="00:01:35.30" entrycourse="SCM" />
                <RESULT eventid="1105" points="203" swimtime="00:01:23.84" resultid="3170" heatid="3450" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="256" swimtime="00:00:31.75" resultid="3171" heatid="3488" lane="2" entrytime="00:00:32.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Julia Rocha" birthdate="2014-02-10" gender="F" nation="BRA" license="397158" swrid="5641767" athleteid="3298" externalid="397158">
              <RESULTS>
                <RESULT eventid="1080" points="158" reactiontime="+60" swimtime="00:00:46.65" resultid="3299" heatid="3419" lane="4" entrytime="00:00:48.80" entrycourse="SCM" />
                <RESULT eventid="1068" points="99" swimtime="00:01:01.29" resultid="3300" heatid="3400" lane="2" />
                <RESULT eventid="1108" points="95" swimtime="00:00:53.29" resultid="3301" heatid="3454" lane="3" entrytime="00:01:12.35" entrycourse="SCM" />
                <RESULT eventid="1128" points="192" swimtime="00:00:39.68" resultid="3302" heatid="3469" lane="3" entrytime="00:00:40.22" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="De Castro Paiva Maciel" birthdate="2008-04-10" gender="M" nation="BRA" license="378333" swrid="5622275" athleteid="3078" externalid="378333">
              <RESULTS>
                <RESULT eventid="1184" points="424" swimtime="00:00:28.95" resultid="3079" heatid="3521" lane="6" entrytime="00:00:31.48" entrycourse="SCM" />
                <RESULT eventid="1216" points="404" swimtime="00:00:27.26" resultid="3080" heatid="3547" lane="1" entrytime="00:00:28.75" entrycourse="SCM" />
                <RESULT eventid="1248" points="417" swimtime="00:00:59.98" resultid="3081" heatid="3574" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Prestes Alves Pinto" birthdate="2012-01-19" gender="F" nation="BRA" license="377324" swrid="5588867" athleteid="3221" externalid="377324">
              <RESULTS>
                <RESULT eventid="1086" points="327" swimtime="00:02:40.05" resultid="3222" heatid="3428" lane="1" entrytime="00:02:45.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.34" />
                    <SPLIT distance="100" swimtime="00:01:18.12" />
                    <SPLIT distance="150" swimtime="00:02:00.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="256" swimtime="00:00:39.75" resultid="3223" heatid="3410" lane="7" entrytime="00:00:38.84" entrycourse="SCM" />
                <RESULT eventid="1102" points="238" swimtime="00:01:31.07" resultid="3224" heatid="3446" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="310" swimtime="00:00:33.87" resultid="3225" heatid="3481" lane="1" entrytime="00:00:33.99" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Marques" birthdate="2007-06-29" gender="M" nation="BRA" license="367257" swrid="5600213" athleteid="3374" externalid="367257">
              <RESULTS>
                <RESULT eventid="1152" points="342" swimtime="00:05:03.38" resultid="3375" heatid="3500" lane="5" entrytime="00:04:48.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.58" />
                    <SPLIT distance="100" swimtime="00:01:08.87" />
                    <SPLIT distance="150" swimtime="00:01:46.76" />
                    <SPLIT distance="200" swimtime="00:02:25.50" />
                    <SPLIT distance="250" swimtime="00:03:05.39" />
                    <SPLIT distance="300" swimtime="00:03:45.31" />
                    <SPLIT distance="350" swimtime="00:04:25.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="353" swimtime="00:01:03.39" resultid="3376" heatid="3578" lane="4" entrytime="00:01:01.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Zattar" birthdate="2012-04-19" gender="F" nation="BRA" license="401736" swrid="5661351" athleteid="3323" externalid="401736">
              <RESULTS>
                <RESULT eventid="1062" points="186" swimtime="00:01:49.09" resultid="3324" heatid="3392" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="245" reactiontime="+77" swimtime="00:00:40.35" resultid="3325" heatid="3406" lane="7" />
                <RESULT eventid="1102" points="196" swimtime="00:01:37.19" resultid="3326" heatid="3443" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="249" swimtime="00:00:36.44" resultid="3327" heatid="3477" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="Moreira Furtado" birthdate="2011-01-27" gender="F" nation="BRA" license="403783" swrid="5684587" athleteid="3356" externalid="403783">
              <RESULTS>
                <RESULT eventid="1208" points="176" swimtime="00:00:40.90" resultid="3357" heatid="3533" lane="2" />
                <RESULT eventid="1240" points="174" swimtime="00:01:29.84" resultid="3358" heatid="3563" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Lucachinski Villatore" birthdate="2013-10-04" gender="M" nation="BRA" license="382248" swrid="5588778" athleteid="3236" externalid="382248">
              <RESULTS>
                <RESULT eventid="1089" points="86" swimtime="00:03:44.37" resultid="3237" heatid="3430" lane="4" entrytime="00:04:40.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.85" />
                    <SPLIT distance="100" swimtime="00:01:45.21" />
                    <SPLIT distance="150" swimtime="00:02:45.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="69" reactiontime="+77" swimtime="00:00:53.74" resultid="3238" heatid="3411" lane="3" />
                <RESULT eventid="1141" points="81" swimtime="00:00:46.57" resultid="3239" heatid="3483" lane="3" entrytime="00:00:46.86" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Andrade Guarido" birthdate="2014-05-17" gender="M" nation="BRA" license="400031" swrid="5652873" athleteid="3315" externalid="400031">
              <RESULTS>
                <RESULT eventid="1083" points="67" reactiontime="+29" swimtime="00:00:54.39" resultid="3316" heatid="3421" lane="7" />
                <RESULT eventid="1071" points="91" swimtime="00:00:55.36" resultid="3317" heatid="3403" lane="1" />
                <RESULT eventid="1131" points="99" swimtime="00:00:43.55" resultid="3318" heatid="3472" lane="4" entrytime="00:00:52.23" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Fachini Kovalski" birthdate="2012-05-15" gender="M" nation="BRA" license="403404" swrid="5676297" athleteid="3348" externalid="403404">
              <RESULTS>
                <RESULT eventid="1077" points="74" reactiontime="+80" swimtime="00:00:52.47" resultid="3349" heatid="3412" lane="2" />
                <RESULT eventid="1141" points="103" swimtime="00:00:43.00" resultid="3350" heatid="3482" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Guizun Jannuzzi" birthdate="2011-12-27" gender="M" nation="BRA" license="367148" swrid="5588732" athleteid="3134" externalid="367148">
              <RESULTS>
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="3135" heatid="3509" lane="4" entrytime="00:01:53.48" entrycourse="SCM" />
                <RESULT eventid="1152" status="DNS" swimtime="00:00:00.00" resultid="3136" heatid="3498" lane="7" entrytime="00:05:57.53" entrycourse="SCM" />
                <RESULT eventid="1216" status="DNS" swimtime="00:00:00.00" resultid="3137" heatid="3544" lane="3" entrytime="00:00:34.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Vianna" birthdate="2011-01-31" gender="M" nation="BRA" license="371380" swrid="5588947" athleteid="3172" externalid="371380">
              <RESULTS>
                <RESULT eventid="1152" points="329" swimtime="00:05:07.38" resultid="3173" heatid="3497" lane="4" entrytime="00:06:22.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:14.78" />
                    <SPLIT distance="150" swimtime="00:01:54.16" />
                    <SPLIT distance="200" swimtime="00:02:33.57" />
                    <SPLIT distance="250" swimtime="00:03:12.18" />
                    <SPLIT distance="300" swimtime="00:03:51.00" />
                    <SPLIT distance="350" swimtime="00:04:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="329" swimtime="00:00:29.18" resultid="3174" heatid="3546" lane="8" entrytime="00:00:30.56" entrycourse="SCM" />
                <RESULT eventid="1248" points="330" swimtime="00:01:04.83" resultid="3175" heatid="3577" lane="3" entrytime="00:01:06.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Gouvea" birthdate="2013-04-19" gender="M" nation="BRA" license="387378" swrid="5588729" athleteid="3259" externalid="387378">
              <RESULTS>
                <RESULT eventid="1089" points="112" swimtime="00:03:26.09" resultid="3260" heatid="3431" lane="2" entrytime="00:03:30.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.64" />
                    <SPLIT distance="100" swimtime="00:01:35.30" />
                    <SPLIT distance="150" swimtime="00:02:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="114" swimtime="00:01:53.97" resultid="3261" heatid="3396" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="144" swimtime="00:00:38.39" resultid="3262" heatid="3484" lane="5" entrytime="00:00:39.48" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Coelho Oliveira" birthdate="2015-03-03" gender="F" nation="BRA" license="406839" athleteid="3385" externalid="406839">
              <RESULTS>
                <RESULT eventid="1080" points="65" reactiontime="+47" swimtime="00:01:02.72" resultid="3386" heatid="3418" lane="2" />
                <RESULT eventid="1068" points="61" swimtime="00:01:11.91" resultid="3387" heatid="3400" lane="1" />
                <RESULT eventid="1128" points="72" swimtime="00:00:55.10" resultid="3388" heatid="3465" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Augusto Vaz" birthdate="2011-06-25" gender="M" nation="BRA" license="401737" swrid="5661339" athleteid="3328" externalid="401737">
              <RESULTS>
                <RESULT eventid="1184" points="194" swimtime="00:00:37.52" resultid="3329" heatid="3519" lane="1" />
                <RESULT eventid="1152" status="DSQ" swimtime="00:00:00.00" resultid="3330" heatid="3496" lane="2" />
                <RESULT eventid="1216" points="241" swimtime="00:00:32.38" resultid="3331" heatid="3542" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Schlickmann Assis" birthdate="2003-07-24" gender="F" nation="BRA" license="303874" swrid="5600257" athleteid="3116" externalid="303874">
              <RESULTS>
                <RESULT eventid="1176" points="479" swimtime="00:00:31.15" resultid="3117" heatid="3515" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Camily Moraes" birthdate="2014-07-13" gender="F" nation="BRA" license="397159" swrid="5641755" athleteid="3303" externalid="397159">
              <RESULTS>
                <RESULT eventid="1092" points="95" swimtime="00:01:49.76" resultid="3304" heatid="3437" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="111" swimtime="00:00:52.39" resultid="3305" heatid="3419" lane="1" entrytime="00:00:55.12" entrycourse="SCM" />
                <RESULT eventid="1128" points="129" swimtime="00:00:45.29" resultid="3306" heatid="3467" lane="4" entrytime="00:00:52.85" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietra" lastname="Vitoria Paczrowski" birthdate="2009-08-12" gender="F" nation="BRA" license="351253" swrid="5600275" athleteid="3108" externalid="351253" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1208" points="460" swimtime="00:00:29.69" resultid="3109" heatid="3539" lane="8" entrytime="00:00:30.22" entrycourse="SCM" />
                <RESULT eventid="1272" points="367" reactiontime="+53" swimtime="00:00:35.26" resultid="3110" heatid="3588" lane="4" entrytime="00:00:36.62" entrycourse="SCM" />
                <RESULT eventid="1240" points="435" swimtime="00:01:06.31" resultid="3111" heatid="3569" lane="1" entrytime="00:01:07.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Zanatta Flizikowski" birthdate="2010-01-08" gender="F" nation="BRA" license="367051" swrid="5588969" athleteid="3367" externalid="367051">
              <RESULTS>
                <RESULT eventid="1176" points="391" swimtime="00:00:33.33" resultid="3368" heatid="3515" lane="6" />
                <RESULT eventid="1240" points="427" swimtime="00:01:06.73" resultid="3369" heatid="3563" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wilson" lastname="Candido Souza" birthdate="2005-04-06" gender="M" nation="BRA" license="256803" swrid="5600129" athleteid="3158" externalid="256803">
              <RESULTS>
                <RESULT eventid="1168" points="501" swimtime="00:01:09.59" resultid="3159" heatid="3512" lane="4" entrytime="00:01:12.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="486" swimtime="00:00:31.73" resultid="3160" heatid="3612" lane="1" entrytime="00:00:32.61" entrycourse="SCM" />
                <RESULT eventid="1248" points="508" swimtime="00:00:56.19" resultid="3161" heatid="3580" lane="7" entrytime="00:00:56.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Coelho De Oliveira" birthdate="2012-11-11" gender="M" nation="BRA" license="385198" swrid="5588600" athleteid="3245" externalid="385198">
              <RESULTS>
                <RESULT eventid="1089" points="105" swimtime="00:03:30.01" resultid="3246" heatid="3429" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.42" />
                    <SPLIT distance="100" swimtime="00:01:40.12" />
                    <SPLIT distance="150" swimtime="00:02:38.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="102" swimtime="00:01:58.21" resultid="3247" heatid="3398" lane="8" entrytime="00:02:07.80" entrycourse="SCM" />
                <RESULT eventid="1141" points="131" swimtime="00:00:39.64" resultid="3248" heatid="3484" lane="7" entrytime="00:00:44.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Franchesca Costa" birthdate="2008-05-19" gender="F" nation="BRA" license="350213" swrid="5600168" athleteid="3150" externalid="350213">
              <RESULTS>
                <RESULT eventid="1208" points="365" swimtime="00:00:32.08" resultid="3151" heatid="3534" lane="8" />
                <RESULT eventid="1192" points="378" reactiontime="+62" swimtime="00:01:15.85" resultid="3152" heatid="3527" lane="1" entrytime="00:01:14.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="385" reactiontime="+63" swimtime="00:00:34.70" resultid="3153" heatid="3589" lane="1" entrytime="00:00:34.20" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otto" lastname="Hedeke" birthdate="2011-03-24" gender="M" nation="BRA" license="372643" swrid="5588738" athleteid="3183" externalid="372643">
              <RESULTS>
                <RESULT eventid="1152" points="253" swimtime="00:05:35.27" resultid="3184" heatid="3498" lane="8" entrytime="00:06:12.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.58" />
                    <SPLIT distance="100" swimtime="00:01:20.12" />
                    <SPLIT distance="150" swimtime="00:02:03.55" />
                    <SPLIT distance="200" swimtime="00:02:46.78" />
                    <SPLIT distance="250" swimtime="00:03:31.46" />
                    <SPLIT distance="300" swimtime="00:04:14.82" />
                    <SPLIT distance="350" swimtime="00:04:55.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="263" swimtime="00:22:00.59" resultid="3185" heatid="3584" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                    <SPLIT distance="100" swimtime="00:01:22.61" />
                    <SPLIT distance="150" swimtime="00:02:07.18" />
                    <SPLIT distance="200" swimtime="00:02:51.55" />
                    <SPLIT distance="250" swimtime="00:03:36.20" />
                    <SPLIT distance="300" swimtime="00:04:20.93" />
                    <SPLIT distance="350" swimtime="00:05:05.61" />
                    <SPLIT distance="400" swimtime="00:05:49.38" />
                    <SPLIT distance="450" swimtime="00:06:33.63" />
                    <SPLIT distance="500" swimtime="00:07:18.47" />
                    <SPLIT distance="550" swimtime="00:08:02.70" />
                    <SPLIT distance="600" swimtime="00:08:46.98" />
                    <SPLIT distance="650" swimtime="00:09:32.06" />
                    <SPLIT distance="700" swimtime="00:10:17.11" />
                    <SPLIT distance="750" swimtime="00:11:01.37" />
                    <SPLIT distance="800" swimtime="00:11:47.35" />
                    <SPLIT distance="850" swimtime="00:12:31.48" />
                    <SPLIT distance="900" swimtime="00:13:16.51" />
                    <SPLIT distance="950" swimtime="00:14:01.77" />
                    <SPLIT distance="1000" swimtime="00:14:46.85" />
                    <SPLIT distance="1050" swimtime="00:15:30.46" />
                    <SPLIT distance="1100" swimtime="00:16:15.25" />
                    <SPLIT distance="1150" swimtime="00:17:00.54" />
                    <SPLIT distance="1200" swimtime="00:17:43.71" />
                    <SPLIT distance="1250" swimtime="00:18:28.56" />
                    <SPLIT distance="1300" swimtime="00:19:13.02" />
                    <SPLIT distance="1350" swimtime="00:19:57.06" />
                    <SPLIT distance="1400" swimtime="00:20:40.47" />
                    <SPLIT distance="1450" swimtime="00:21:22.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Marques Machado" birthdate="2010-02-17" gender="M" nation="BRA" license="390918" swrid="5600212" athleteid="3281" externalid="390918">
              <RESULTS>
                <RESULT eventid="1184" status="DNS" swimtime="00:00:00.00" resultid="3282" heatid="3518" lane="7" />
                <RESULT eventid="1152" status="DNS" swimtime="00:00:00.00" resultid="3283" heatid="3495" lane="2" />
                <RESULT eventid="1248" status="DNS" swimtime="00:00:00.00" resultid="3284" heatid="3575" lane="2" entrytime="00:01:23.29" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cleverson" lastname="Cardoso" birthdate="2013-07-20" gender="M" nation="BRA" license="387382" swrid="5588577" athleteid="3267" externalid="387382">
              <RESULTS>
                <RESULT eventid="1077" points="85" reactiontime="+81" swimtime="00:00:50.19" resultid="3268" heatid="3413" lane="3" entrytime="00:00:51.67" entrycourse="SCM" />
                <RESULT eventid="1065" points="93" swimtime="00:02:01.81" resultid="3269" heatid="3397" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="93" swimtime="00:00:44.48" resultid="3270" heatid="3484" lane="8" entrytime="00:00:44.26" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Luis Santin Ronchi" birthdate="2007-11-14" gender="M" nation="BRA" license="336738" swrid="5600204" athleteid="3086" externalid="336738">
              <RESULTS>
                <RESULT eventid="1184" points="439" swimtime="00:00:28.61" resultid="3087" heatid="3519" lane="5" />
                <RESULT eventid="1168" points="425" swimtime="00:01:13.48" resultid="3088" heatid="3512" lane="5" entrytime="00:01:13.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="433" swimtime="00:02:24.85" resultid="3089" heatid="3561" lane="7" entrytime="00:02:20.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.59" />
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                    <SPLIT distance="150" swimtime="00:01:50.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="427" swimtime="00:00:33.12" resultid="3090" heatid="3611" lane="5" entrytime="00:00:33.48" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Rodrigues Bortoluzzi" birthdate="2013-10-07" gender="M" nation="BRA" license="387375" swrid="5652897" athleteid="3252" externalid="387375">
              <RESULTS>
                <RESULT eventid="1077" points="73" reactiontime="+142" swimtime="00:00:52.88" resultid="3253" heatid="3413" lane="6" entrytime="00:00:54.77" entrycourse="SCM" />
                <RESULT eventid="1141" points="125" swimtime="00:00:40.24" resultid="3254" heatid="3484" lane="4" entrytime="00:00:39.46" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Nalle Bejes" birthdate="2010-04-20" gender="F" nation="BRA" license="377323" swrid="5588826" athleteid="3217" externalid="377323">
              <RESULTS>
                <RESULT eventid="1144" points="386" swimtime="00:05:17.56" resultid="3218" heatid="3491" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                    <SPLIT distance="100" swimtime="00:01:15.13" />
                    <SPLIT distance="150" swimtime="00:01:55.10" />
                    <SPLIT distance="200" swimtime="00:02:35.58" />
                    <SPLIT distance="250" swimtime="00:03:16.12" />
                    <SPLIT distance="300" swimtime="00:03:57.26" />
                    <SPLIT distance="350" swimtime="00:04:37.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" status="DSQ" swimtime="00:03:00.10" resultid="3219" heatid="3553" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                    <SPLIT distance="100" swimtime="00:01:27.93" />
                    <SPLIT distance="150" swimtime="00:02:21.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="346" swimtime="00:00:40.39" resultid="3220" heatid="3604" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diego" lastname="Brasil Caropreso" birthdate="2009-10-29" gender="M" nation="BRA" license="399502" swrid="5653287" athleteid="3370" externalid="399502">
              <RESULTS>
                <RESULT eventid="1184" points="305" swimtime="00:00:32.28" resultid="3371" heatid="3520" lane="4" entrytime="00:00:42.57" entrycourse="SCM" />
                <RESULT eventid="1216" points="356" swimtime="00:00:28.43" resultid="3372" heatid="3547" lane="6" entrytime="00:00:28.33" entrycourse="SCM" />
                <RESULT eventid="1248" points="356" swimtime="00:01:03.21" resultid="3373" heatid="3578" lane="8" entrytime="00:01:05.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carol" lastname="Nalle Bejes" birthdate="2010-04-20" gender="F" nation="BRA" license="377315" swrid="5588824" athleteid="3196" externalid="377315">
              <RESULTS>
                <RESULT eventid="1144" points="372" swimtime="00:05:21.52" resultid="3197" heatid="3489" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="100" swimtime="00:01:15.59" />
                    <SPLIT distance="150" swimtime="00:01:56.39" />
                    <SPLIT distance="200" swimtime="00:02:36.98" />
                    <SPLIT distance="250" swimtime="00:03:17.54" />
                    <SPLIT distance="300" swimtime="00:03:59.62" />
                    <SPLIT distance="350" swimtime="00:04:41.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="348" swimtime="00:00:32.59" resultid="3198" heatid="3536" lane="3" entrytime="00:00:34.72" entrycourse="SCM" />
                <RESULT eventid="1304" points="408" swimtime="00:00:38.25" resultid="3199" heatid="3603" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Wenceslau Bitencourt" birthdate="2012-02-11" gender="M" nation="BRA" license="377318" swrid="5602591" athleteid="3209" externalid="377318">
              <RESULTS>
                <RESULT eventid="1089" points="198" swimtime="00:02:50.24" resultid="3210" heatid="3429" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                    <SPLIT distance="100" swimtime="00:01:23.65" />
                    <SPLIT distance="150" swimtime="00:02:07.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="162" reactiontime="+72" swimtime="00:00:40.55" resultid="3211" heatid="3414" lane="6" entrytime="00:00:43.76" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lis" lastname="Cristini Harmatiuk" birthdate="2014-07-19" gender="F" nation="BRA" license="396830" swrid="5641759" athleteid="3362" externalid="396830">
              <RESULTS>
                <RESULT eventid="1080" points="135" reactiontime="+67" swimtime="00:00:49.22" resultid="3363" heatid="3419" lane="3" entrytime="00:00:50.61" entrycourse="SCM" />
                <RESULT eventid="1068" points="162" swimtime="00:00:52.00" resultid="3364" heatid="3401" lane="6" entrytime="00:00:57.42" entrycourse="SCM" />
                <RESULT eventid="1108" points="95" swimtime="00:00:53.30" resultid="3365" heatid="3452" lane="4" />
                <RESULT eventid="1128" points="165" swimtime="00:00:41.73" resultid="3366" heatid="3469" lane="2" entrytime="00:00:43.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helenna" lastname="Banzatto Silva" birthdate="2013-07-11" gender="F" nation="BRA" license="393210" swrid="5616439" athleteid="3294" externalid="393210">
              <RESULTS>
                <RESULT eventid="1062" points="109" swimtime="00:02:10.24" resultid="3295" heatid="3392" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="40" swimtime="00:01:13.25" resultid="3296" heatid="3408" lane="8" entrytime="00:01:18.29" entrycourse="SCM" />
                <RESULT eventid="1138" points="47" swimtime="00:01:03.21" resultid="3297" heatid="3476" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="De Siqueira Machado" birthdate="2012-05-25" gender="F" nation="BRA" license="377312" swrid="5588649" athleteid="3186" externalid="377312">
              <RESULTS>
                <RESULT eventid="1086" points="262" swimtime="00:02:52.37" resultid="3187" heatid="3427" lane="6" entrytime="00:02:52.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="100" swimtime="00:01:22.22" />
                    <SPLIT distance="150" swimtime="00:02:08.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="237" swimtime="00:00:40.76" resultid="3188" heatid="3410" lane="1" entrytime="00:00:40.57" entrycourse="SCM" />
                <RESULT eventid="1102" points="250" swimtime="00:01:29.66" resultid="3189" heatid="3445" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="330" swimtime="00:00:33.15" resultid="3190" heatid="3481" lane="7" entrytime="00:00:33.78" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helloisa" lastname="De Bassani" birthdate="2012-09-23" gender="F" nation="BRA" license="403403" swrid="5676296" athleteid="3344" externalid="403403">
              <RESULTS>
                <RESULT eventid="1062" points="59" swimtime="00:02:39.30" resultid="3345" heatid="3394" lane="8" />
                <RESULT eventid="1074" points="72" reactiontime="+83" swimtime="00:01:00.61" resultid="3346" heatid="3406" lane="2" />
                <RESULT eventid="1138" points="116" swimtime="00:00:46.92" resultid="3347" heatid="3477" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Celli Schneider" birthdate="2011-02-21" gender="M" nation="BRA" license="367055" swrid="5588587" athleteid="3130" externalid="367055">
              <RESULTS>
                <RESULT eventid="1200" points="265" reactiontime="+46" swimtime="00:01:15.19" resultid="3131" heatid="3530" lane="3" entrytime="00:01:19.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="315" swimtime="00:05:11.63" resultid="3132" heatid="3495" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.27" />
                    <SPLIT distance="100" swimtime="00:01:15.89" />
                    <SPLIT distance="150" swimtime="00:01:56.15" />
                    <SPLIT distance="200" swimtime="00:02:35.85" />
                    <SPLIT distance="250" swimtime="00:03:14.90" />
                    <SPLIT distance="300" swimtime="00:03:54.48" />
                    <SPLIT distance="350" swimtime="00:04:32.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="276" reactiontime="+57" swimtime="00:00:33.93" resultid="3133" heatid="3592" lane="4" entrytime="00:00:35.17" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Hoffmann Zoschke" birthdate="2015-03-22" gender="M" nation="BRA" license="390917" swrid="5602547" athleteid="3276" externalid="390917">
              <RESULTS>
                <RESULT eventid="1095" points="124" swimtime="00:01:29.92" resultid="3277" heatid="3440" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="85" swimtime="00:00:56.60" resultid="3278" heatid="3404" lane="2" entrytime="00:01:01.35" entrycourse="SCM" />
                <RESULT eventid="1111" points="99" swimtime="00:00:46.92" resultid="3279" heatid="3458" lane="4" entrytime="00:00:58.15" entrycourse="SCM" />
                <RESULT eventid="1131" points="129" swimtime="00:00:39.88" resultid="3280" heatid="3473" lane="5" entrytime="00:00:43.26" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Ryan Rosa" birthdate="2014-01-14" gender="M" nation="BRA" license="400032" swrid="5652898" athleteid="3319" externalid="400032">
              <RESULTS>
                <RESULT eventid="1095" points="58" swimtime="00:01:55.43" resultid="3320" heatid="3440" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="74" swimtime="00:00:59.34" resultid="3321" heatid="3402" lane="2" />
                <RESULT eventid="1131" points="62" swimtime="00:00:50.67" resultid="3322" heatid="3472" lane="5" entrytime="00:00:52.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kethelyn" lastname="Ribeiro Da Silva Rodrigues" birthdate="2009-04-24" gender="F" nation="BRA" license="367052" swrid="5600244" athleteid="3122" externalid="367052">
              <RESULTS>
                <RESULT eventid="1208" points="417" swimtime="00:00:30.69" resultid="3123" heatid="3537" lane="3" entrytime="00:00:32.16" entrycourse="SCM" />
                <RESULT eventid="1272" points="281" reactiontime="+57" swimtime="00:00:38.51" resultid="3124" heatid="3587" lane="2" />
                <RESULT eventid="1240" points="411" swimtime="00:01:07.56" resultid="3125" heatid="3568" lane="1" entrytime="00:01:10.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Luiza Rocha Batista" birthdate="2013-11-24" gender="F" nation="BRA" license="387379" swrid="5588784" athleteid="3263" externalid="387379">
              <RESULTS>
                <RESULT eventid="1074" points="114" reactiontime="+71" swimtime="00:00:52.02" resultid="3264" heatid="3408" lane="6" entrytime="00:00:53.63" entrycourse="SCM" />
                <RESULT eventid="1118" points="79" swimtime="00:02:05.67" resultid="3265" heatid="3461" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="145" swimtime="00:00:43.57" resultid="3266" heatid="3479" lane="5" entrytime="00:00:40.87" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tais" lastname="Feltrin Martins" birthdate="2013-01-17" gender="F" nation="BRA" license="406840" athleteid="3389" externalid="406840">
              <RESULTS>
                <RESULT eventid="1074" points="85" reactiontime="+70" swimtime="00:00:57.24" resultid="3390" heatid="3407" lane="6" />
                <RESULT eventid="1138" points="80" swimtime="00:00:53.03" resultid="3391" heatid="3476" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Bello Costa Lange" birthdate="2013-07-17" gender="M" nation="BRA" license="377319" swrid="5588548" athleteid="3212" externalid="377319">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="3213" heatid="3432" lane="5" entrytime="00:02:57.70" entrycourse="SCM" />
                <RESULT eventid="1065" status="DNS" swimtime="00:00:00.00" resultid="3214" heatid="3396" lane="7" />
                <RESULT eventid="1105" points="145" swimtime="00:01:33.60" resultid="3215" heatid="3451" lane="7" entrytime="00:01:38.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1121" points="74" swimtime="00:01:53.78" resultid="3216" heatid="3463" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Blansky Hagebock" birthdate="2008-08-15" gender="M" nation="BRA" license="339123" swrid="5455418" athleteid="3104" externalid="339123">
              <RESULTS>
                <RESULT eventid="1184" points="421" swimtime="00:00:29.00" resultid="3105" heatid="3521" lane="3" entrytime="00:00:30.65" entrycourse="SCM" />
                <RESULT eventid="1216" points="462" swimtime="00:00:26.07" resultid="3106" heatid="3549" lane="8" entrytime="00:00:26.63" entrycourse="SCM" />
                <RESULT eventid="1248" points="511" swimtime="00:00:56.08" resultid="3107" heatid="3579" lane="4" entrytime="00:00:59.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="F" nation="BRA" license="344301" swrid="5569976" athleteid="3060" externalid="344301">
              <RESULTS>
                <RESULT eventid="1144" points="547" swimtime="00:04:42.67" resultid="3061" heatid="3492" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                    <SPLIT distance="100" swimtime="00:01:03.66" />
                    <SPLIT distance="150" swimtime="00:01:39.52" />
                    <SPLIT distance="200" swimtime="00:02:16.10" />
                    <SPLIT distance="250" swimtime="00:02:53.09" />
                    <SPLIT distance="300" swimtime="00:03:30.24" />
                    <SPLIT distance="350" swimtime="00:04:07.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="538" swimtime="00:01:06.43" resultid="3062" heatid="3596" lane="3" entrytime="00:01:06.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="558" swimtime="00:01:01.03" resultid="3063" heatid="3570" lane="2" entrytime="00:01:04.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mathias" lastname="Bernardo" birthdate="2014-05-17" gender="M" nation="BRA" license="387376" swrid="5652880" athleteid="3255" externalid="387376">
              <RESULTS>
                <RESULT eventid="1095" points="48" swimtime="00:02:02.82" resultid="3256" heatid="3441" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="38" swimtime="00:01:05.66" resultid="3257" heatid="3422" lane="3" entrytime="00:01:08.82" entrycourse="SCM" />
                <RESULT eventid="1131" points="74" swimtime="00:00:47.97" resultid="3258" heatid="3472" lane="2" entrytime="00:00:57.27" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Araujo Felix" birthdate="2010-05-27" gender="F" nation="BRA" license="393157" swrid="5622260" athleteid="3381" externalid="393157">
              <RESULTS>
                <RESULT eventid="1144" status="DNS" swimtime="00:00:00.00" resultid="3382" heatid="3489" lane="6" />
                <RESULT eventid="1176" status="DNS" swimtime="00:00:00.00" resultid="3383" heatid="3514" lane="3" />
                <RESULT eventid="1240" status="DNS" swimtime="00:00:00.00" resultid="3384" heatid="3563" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Inoue Kuroda" birthdate="2009-04-18" gender="M" nation="BRA" license="324700" swrid="5600190" athleteid="3096" externalid="324700">
              <RESULTS>
                <RESULT eventid="1200" points="400" reactiontime="+68" swimtime="00:01:05.59" resultid="3097" heatid="3532" lane="1" entrytime="00:01:08.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="434" swimtime="00:00:26.61" resultid="3098" heatid="3543" lane="2" />
                <RESULT eventid="1248" points="460" swimtime="00:00:58.06" resultid="3099" heatid="3579" lane="8" entrytime="00:01:00.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Bello Costa Lange" birthdate="2010-09-13" gender="M" nation="BRA" license="367152" swrid="5588547" athleteid="3146" externalid="367152">
              <RESULTS>
                <RESULT eventid="1184" points="303" swimtime="00:00:32.36" resultid="3147" heatid="3520" lane="7" />
                <RESULT eventid="1152" points="340" swimtime="00:05:03.98" resultid="3148" heatid="3497" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:10.88" />
                    <SPLIT distance="150" swimtime="00:01:49.38" />
                    <SPLIT distance="200" swimtime="00:02:28.30" />
                    <SPLIT distance="250" swimtime="00:03:07.24" />
                    <SPLIT distance="300" swimtime="00:03:46.55" />
                    <SPLIT distance="350" swimtime="00:04:25.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="301" swimtime="00:01:11.24" resultid="3149" heatid="3601" lane="8" entrytime="00:01:13.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauren" lastname="Kurecki" birthdate="2014-03-06" gender="F" nation="BRA" license="377314" swrid="5602549" athleteid="3191" externalid="377314">
              <RESULTS>
                <RESULT eventid="1092" points="258" swimtime="00:01:18.93" resultid="3192" heatid="3438" lane="4" entrytime="00:01:23.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="227" swimtime="00:00:46.45" resultid="3193" heatid="3401" lane="4" entrytime="00:00:47.75" entrycourse="SCM" />
                <RESULT eventid="1108" points="206" swimtime="00:00:41.26" resultid="3194" heatid="3455" lane="4" entrytime="00:00:46.20" entrycourse="SCM" />
                <RESULT eventid="1128" points="300" swimtime="00:00:34.25" resultid="3195" heatid="3469" lane="4" entrytime="00:00:37.67" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2864" nation="BRA" region="PR" clubid="1320" swrid="93756" name="Associacao De Pais E Amigos Da Natacao De Ponta Gr" shortname="Apan Ponta Grossa">
          <ATHLETES>
            <ATHLETE firstname="Arthur" lastname="Dolinski Thomassewski" birthdate="2006-12-15" gender="M" nation="BRA" license="400409" swrid="5653289" athleteid="1417" externalid="400409">
              <RESULTS>
                <RESULT eventid="1216" points="309" swimtime="00:00:29.79" resultid="1418" heatid="3540" lane="4" />
                <RESULT eventid="1312" points="259" swimtime="00:00:39.11" resultid="1419" heatid="3608" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Allana" lastname="Lacerda" birthdate="2005-03-15" gender="F" nation="BRA" license="295186" swrid="5600197" athleteid="1336" externalid="295186" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1176" points="385" swimtime="00:00:33.50" resultid="1337" heatid="3515" lane="7" />
                <RESULT eventid="1160" points="443" swimtime="00:01:21.78" resultid="1338" heatid="3506" lane="7" entrytime="00:01:21.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="420" swimtime="00:02:42.66" resultid="1339" heatid="3556" lane="3" entrytime="00:02:37.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.98" />
                    <SPLIT distance="100" swimtime="00:01:19.42" />
                    <SPLIT distance="150" swimtime="00:02:04.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="416" swimtime="00:00:37.99" resultid="1340" heatid="3606" lane="2" entrytime="00:00:38.27" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Victoria Borges" birthdate="2014-01-16" gender="F" nation="BRA" license="376737" swrid="5602587" athleteid="1389" externalid="376737">
              <RESULTS>
                <RESULT eventid="1092" points="149" swimtime="00:01:34.62" resultid="1390" heatid="3438" lane="1" entrytime="00:01:46.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1080" points="152" reactiontime="+73" swimtime="00:00:47.28" resultid="1391" heatid="3419" lane="2" entrytime="00:00:51.22" entrycourse="SCM" />
                <RESULT eventid="1108" points="72" swimtime="00:00:58.51" resultid="1392" heatid="3453" lane="8" />
                <RESULT eventid="1128" points="186" swimtime="00:00:40.10" resultid="1393" heatid="3469" lane="8" entrytime="00:00:45.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Chi Kravchychyn" birthdate="2009-09-27" gender="M" nation="BRA" license="344268" swrid="5600134" athleteid="1327" externalid="344268">
              <RESULTS>
                <RESULT eventid="1184" points="452" swimtime="00:00:28.33" resultid="1328" heatid="3520" lane="2" />
                <RESULT eventid="1168" points="502" swimtime="00:01:09.51" resultid="1329" heatid="3513" lane="7" entrytime="00:01:08.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="495" swimtime="00:02:18.51" resultid="1330" heatid="3561" lane="1" entrytime="00:02:20.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                    <SPLIT distance="100" swimtime="00:01:06.61" />
                    <SPLIT distance="150" swimtime="00:01:46.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="465" swimtime="00:00:32.19" resultid="1331" heatid="3612" lane="8" entrytime="00:00:32.83" entrycourse="SCM" />
                <RESULT eventid="1280" points="342" reactiontime="+68" swimtime="00:00:31.60" resultid="1332" heatid="3592" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fegert" birthdate="2009-04-13" gender="M" nation="BRA" license="353813" swrid="5622279" athleteid="1355" externalid="353813">
              <RESULTS>
                <RESULT eventid="1184" points="364" swimtime="00:00:30.46" resultid="1356" heatid="3520" lane="6" />
                <RESULT eventid="1216" points="384" swimtime="00:00:27.72" resultid="1357" heatid="3544" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Carraro Borges" birthdate="2009-05-11" gender="M" nation="BRA" license="345590" swrid="5622267" athleteid="1358" externalid="345590" level="SAGRADA FA">
              <RESULTS>
                <RESULT eventid="1152" points="412" swimtime="00:04:45.21" resultid="1359" heatid="3500" lane="3" entrytime="00:04:49.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.16" />
                    <SPLIT distance="100" swimtime="00:01:06.04" />
                    <SPLIT distance="150" swimtime="00:01:41.52" />
                    <SPLIT distance="200" swimtime="00:02:17.81" />
                    <SPLIT distance="250" swimtime="00:02:54.64" />
                    <SPLIT distance="300" swimtime="00:03:31.57" />
                    <SPLIT distance="350" swimtime="00:04:08.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="372" swimtime="00:00:28.03" resultid="1360" heatid="3543" lane="6" />
                <RESULT eventid="1264" points="422" swimtime="00:18:48.99" resultid="1361" heatid="3585" lane="3" entrytime="00:19:23.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.66" />
                    <SPLIT distance="100" swimtime="00:01:08.91" />
                    <SPLIT distance="150" swimtime="00:01:45.84" />
                    <SPLIT distance="200" swimtime="00:02:23.24" />
                    <SPLIT distance="250" swimtime="00:03:00.47" />
                    <SPLIT distance="300" swimtime="00:03:38.24" />
                    <SPLIT distance="350" swimtime="00:04:16.17" />
                    <SPLIT distance="400" swimtime="00:04:55.41" />
                    <SPLIT distance="450" swimtime="00:05:33.80" />
                    <SPLIT distance="500" swimtime="00:06:12.18" />
                    <SPLIT distance="550" swimtime="00:06:50.70" />
                    <SPLIT distance="600" swimtime="00:07:29.50" />
                    <SPLIT distance="650" swimtime="00:08:07.95" />
                    <SPLIT distance="700" swimtime="00:08:46.32" />
                    <SPLIT distance="750" swimtime="00:09:24.53" />
                    <SPLIT distance="800" swimtime="00:10:01.81" />
                    <SPLIT distance="850" swimtime="00:10:39.46" />
                    <SPLIT distance="900" swimtime="00:11:17.67" />
                    <SPLIT distance="950" swimtime="00:11:55.46" />
                    <SPLIT distance="1000" swimtime="00:12:33.89" />
                    <SPLIT distance="1050" swimtime="00:13:11.80" />
                    <SPLIT distance="1100" swimtime="00:13:49.74" />
                    <SPLIT distance="1150" swimtime="00:14:27.39" />
                    <SPLIT distance="1200" swimtime="00:15:05.50" />
                    <SPLIT distance="1250" swimtime="00:15:43.08" />
                    <SPLIT distance="1300" swimtime="00:16:20.52" />
                    <SPLIT distance="1350" swimtime="00:16:58.30" />
                    <SPLIT distance="1400" swimtime="00:17:36.04" />
                    <SPLIT distance="1450" swimtime="00:18:13.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Sabedotti" birthdate="2011-04-20" gender="F" nation="BRA" license="390877" swrid="5602580" athleteid="1397" externalid="390877">
              <RESULTS>
                <RESULT eventid="1208" points="407" swimtime="00:00:30.93" resultid="1398" heatid="3537" lane="5" entrytime="00:00:31.82" entrycourse="SCM" />
                <RESULT eventid="1176" points="349" swimtime="00:00:34.61" resultid="1399" heatid="3515" lane="1" />
                <RESULT eventid="1272" points="335" reactiontime="+56" swimtime="00:00:36.35" resultid="1400" heatid="3588" lane="5" entrytime="00:00:37.43" entrycourse="SCM" />
                <RESULT eventid="1240" points="390" swimtime="00:01:08.77" resultid="1401" heatid="3567" lane="5" entrytime="00:01:10.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Seifert Klas" birthdate="2012-12-17" gender="F" nation="BRA" license="406934" athleteid="1424" externalid="406934">
              <RESULTS>
                <RESULT eventid="1086" points="128" swimtime="00:03:38.56" resultid="1425" heatid="3425" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.70" />
                    <SPLIT distance="100" swimtime="00:01:42.72" />
                    <SPLIT distance="150" swimtime="00:02:42.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="132" reactiontime="+41" swimtime="00:00:49.52" resultid="1426" heatid="3407" lane="1" />
                <RESULT eventid="1138" points="143" swimtime="00:00:43.79" resultid="1427" heatid="3477" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yohan" lastname="Rigoni Moraes" birthdate="2002-04-03" gender="M" nation="BRA" license="272187" swrid="5600245" athleteid="1333" externalid="272187" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1168" points="603" swimtime="00:01:05.42" resultid="1334" heatid="3513" lane="3" entrytime="00:01:04.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="638" swimtime="00:00:28.97" resultid="1335" heatid="3612" lane="5" entrytime="00:00:29.46" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Hilgenberg Lievore" birthdate="2014-04-23" gender="M" nation="BRA" license="391167" swrid="5602546" athleteid="1407" externalid="391167">
              <RESULTS>
                <RESULT eventid="1095" points="133" swimtime="00:01:27.75" resultid="1408" heatid="3442" lane="3" entrytime="00:01:30.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="123" swimtime="00:00:44.41" resultid="1409" heatid="3423" lane="6" entrytime="00:00:48.58" entrycourse="SCM" />
                <RESULT eventid="1111" points="63" swimtime="00:00:54.66" resultid="1410" heatid="3457" lane="5" />
                <RESULT eventid="1131" points="145" swimtime="00:00:38.36" resultid="1411" heatid="3474" lane="6" entrytime="00:00:40.42" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Clara Domingues" birthdate="2012-01-19" gender="F" nation="BRA" license="377291" swrid="5588599" athleteid="1394" externalid="377291">
              <RESULTS>
                <RESULT eventid="1086" points="186" swimtime="00:03:13.17" resultid="1395" heatid="3424" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.90" />
                    <SPLIT distance="100" swimtime="00:01:35.48" />
                    <SPLIT distance="150" swimtime="00:02:25.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="135" reactiontime="+77" swimtime="00:00:49.20" resultid="1396" heatid="3408" lane="5" entrytime="00:00:51.30" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Delinski" birthdate="2009-11-28" gender="F" nation="BRA" license="385190" swrid="5600150" athleteid="1351" externalid="385190">
              <RESULTS>
                <RESULT eventid="1160" points="319" swimtime="00:01:31.21" resultid="1352" heatid="3504" lane="3" entrytime="00:01:32.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" status="DSQ" swimtime="00:03:11.17" resultid="1353" heatid="3552" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:01:30.53" />
                    <SPLIT distance="150" swimtime="00:02:23.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="311" swimtime="00:00:41.86" resultid="1354" heatid="3606" lane="8" entrytime="00:00:42.63" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Campagnoli" birthdate="2009-04-13" gender="F" nation="BRA" license="366915" swrid="5600128" athleteid="1341" externalid="366915">
              <RESULTS>
                <RESULT eventid="1208" points="478" swimtime="00:00:29.31" resultid="1342" heatid="3538" lane="6" entrytime="00:00:31.19" entrycourse="SCM" />
                <RESULT eventid="1192" points="423" reactiontime="+73" swimtime="00:01:13.11" resultid="1343" heatid="3527" lane="7" entrytime="00:01:14.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="459" reactiontime="+68" swimtime="00:00:32.73" resultid="1344" heatid="3589" lane="7" entrytime="00:00:33.73" entrycourse="SCM" />
                <RESULT eventid="1240" points="462" swimtime="00:01:04.99" resultid="1345" heatid="3569" lane="3" entrytime="00:01:06.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Clara Rigailo" birthdate="2013-04-06" gender="F" nation="BRA" license="396828" swrid="5641758" athleteid="1412" externalid="396828">
              <RESULTS>
                <RESULT eventid="1062" points="197" swimtime="00:01:47.13" resultid="1413" heatid="3393" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="140" reactiontime="+81" swimtime="00:00:48.58" resultid="1414" heatid="3408" lane="4" entrytime="00:00:50.78" entrycourse="SCM" />
                <RESULT eventid="1102" points="176" swimtime="00:01:40.68" resultid="1415" heatid="3443" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="202" swimtime="00:00:39.03" resultid="1416" heatid="3478" lane="3" entrytime="00:00:44.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariana" lastname="Brunetti Silva" birthdate="2014-03-24" gender="F" nation="BRA" license="390878" swrid="5602517" athleteid="1402" externalid="390878">
              <RESULTS>
                <RESULT eventid="1092" points="128" swimtime="00:01:39.67" resultid="1403" heatid="3438" lane="7" entrytime="00:01:44.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="107" swimtime="00:00:59.75" resultid="1404" heatid="3400" lane="4" entrytime="00:01:09.92" entrycourse="SCM" />
                <RESULT eventid="1108" points="61" swimtime="00:01:01.91" resultid="1405" heatid="3454" lane="5" entrytime="00:01:05.18" entrycourse="SCM" />
                <RESULT eventid="1128" points="133" swimtime="00:00:44.92" resultid="1406" heatid="3469" lane="1" entrytime="00:00:44.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Franca Berger" birthdate="2010-05-07" gender="F" nation="BRA" license="399692" swrid="5653290" athleteid="1379" externalid="399692">
              <RESULTS>
                <RESULT eventid="1208" points="262" swimtime="00:00:35.83" resultid="1380" heatid="3535" lane="3" entrytime="00:00:39.02" entrycourse="SCM" />
                <RESULT eventid="1160" points="227" swimtime="00:01:42.18" resultid="1381" heatid="3503" lane="4" entrytime="00:01:51.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="251" swimtime="00:00:44.95" resultid="1382" heatid="3605" lane="7" entrytime="00:00:51.87" entrycourse="SCM" />
                <RESULT eventid="1240" points="256" swimtime="00:01:19.07" resultid="1383" heatid="3564" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Carolina Babiuki" birthdate="2007-02-06" gender="F" nation="BRA" license="316227" swrid="5600131" athleteid="1346" externalid="316227" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1208" points="478" swimtime="00:00:29.32" resultid="1347" heatid="3539" lane="3" entrytime="00:00:28.97" entrycourse="SCM" />
                <RESULT eventid="1192" points="423" reactiontime="+72" swimtime="00:01:13.08" resultid="1348" heatid="3527" lane="2" entrytime="00:01:10.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="475" reactiontime="+68" swimtime="00:00:32.35" resultid="1349" heatid="3589" lane="2" entrytime="00:00:32.09" entrycourse="SCM" />
                <RESULT eventid="1240" points="440" swimtime="00:01:06.05" resultid="1350" heatid="3570" lane="6" entrytime="00:01:03.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Bischof Rogoski" birthdate="2014-10-03" gender="M" nation="BRA" license="401860" swrid="5661341" athleteid="1420" externalid="401860">
              <RESULTS>
                <RESULT eventid="1095" points="112" swimtime="00:01:32.99" resultid="1421" heatid="3440" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="90" swimtime="00:00:55.51" resultid="1422" heatid="3403" lane="4" />
                <RESULT eventid="1131" points="133" swimtime="00:00:39.48" resultid="1423" heatid="3470" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Gueiber Montes" birthdate="2009-03-09" gender="M" nation="BRA" license="342154" swrid="5600179" athleteid="1321" externalid="342154">
              <RESULTS>
                <RESULT eventid="1200" points="510" reactiontime="+60" swimtime="00:01:00.46" resultid="1322" heatid="3532" lane="3" entrytime="00:01:01.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="507" swimtime="00:00:25.27" resultid="1323" heatid="3549" lane="7" entrytime="00:00:26.38" entrycourse="SCM" />
                <RESULT eventid="1296" points="348" swimtime="00:01:07.89" resultid="1324" heatid="3597" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1280" points="488" reactiontime="+41" swimtime="00:00:28.07" resultid="1325" heatid="3593" lane="2" entrytime="00:00:28.69" entrycourse="SCM" />
                <RESULT eventid="1248" points="561" swimtime="00:00:54.36" resultid="1326" heatid="3580" lane="3" entrytime="00:00:56.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Brenda" lastname="Gabriele Carvalho" birthdate="2010-04-11" gender="F" nation="BRA" license="399557" swrid="5658060" athleteid="1367" externalid="399557">
              <RESULTS>
                <RESULT eventid="1208" points="231" swimtime="00:00:37.37" resultid="1368" heatid="3535" lane="1" entrytime="00:00:40.13" entrycourse="SCM" />
                <RESULT eventid="1160" points="239" swimtime="00:01:40.38" resultid="1369" heatid="3502" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="208" swimtime="00:00:47.82" resultid="1370" heatid="3604" lane="6" />
                <RESULT eventid="1272" points="250" reactiontime="+72" swimtime="00:00:40.04" resultid="1371" heatid="3587" lane="4" entrytime="00:00:47.77" entrycourse="SCM" />
                <RESULT eventid="1240" points="227" swimtime="00:01:22.35" resultid="1372" heatid="3565" lane="8" entrytime="00:01:32.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Campagnoli" birthdate="2013-03-13" gender="M" nation="BRA" license="370651" swrid="5602519" athleteid="1384" externalid="370651">
              <RESULTS>
                <RESULT eventid="1089" points="239" swimtime="00:02:39.95" resultid="1385" heatid="3434" lane="8" entrytime="00:02:45.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.82" />
                    <SPLIT distance="100" swimtime="00:01:18.39" />
                    <SPLIT distance="150" swimtime="00:02:00.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1077" points="234" reactiontime="+79" swimtime="00:00:35.86" resultid="1386" heatid="3413" lane="7" />
                <RESULT eventid="1121" points="209" swimtime="00:01:20.50" resultid="1387" heatid="3463" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="270" swimtime="00:00:31.16" resultid="1388" heatid="3488" lane="6" entrytime="00:00:31.90" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Augusto" lastname="Tramontin" birthdate="2011-11-29" gender="M" nation="BRA" license="399691" swrid="5652901" athleteid="1373" externalid="399691">
              <RESULTS>
                <RESULT eventid="1200" points="247" reactiontime="+93" swimtime="00:01:16.99" resultid="1374" heatid="3529" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="307" swimtime="00:00:29.87" resultid="1375" heatid="3545" lane="7" entrytime="00:00:31.45" entrycourse="SCM" />
                <RESULT eventid="1312" points="214" swimtime="00:00:41.66" resultid="1376" heatid="3609" lane="2" />
                <RESULT eventid="1280" reactiontime="+68" status="DSQ" swimtime="00:00:36.28" resultid="1377" heatid="3592" lane="5" entrytime="00:00:37.69" entrycourse="SCM" />
                <RESULT eventid="1248" points="291" swimtime="00:01:07.64" resultid="1378" heatid="3576" lane="1" entrytime="00:01:14.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yoseph" lastname="Rigoni Moraes" birthdate="2006-04-17" gender="M" nation="BRA" license="295182" swrid="5622302" athleteid="1362" externalid="295182" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1184" points="492" swimtime="00:00:27.54" resultid="1363" heatid="3522" lane="6" entrytime="00:00:28.50" entrycourse="SCM" />
                <RESULT eventid="1216" points="458" swimtime="00:00:26.15" resultid="1364" heatid="3549" lane="5" entrytime="00:00:26.01" entrycourse="SCM" />
                <RESULT eventid="1312" points="450" swimtime="00:00:32.54" resultid="1365" heatid="3611" lane="4" entrytime="00:00:33.43" entrycourse="SCM" />
                <RESULT eventid="1264" points="393" swimtime="00:19:15.38" resultid="1366" heatid="3584" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.76" />
                    <SPLIT distance="100" swimtime="00:01:03.83" />
                    <SPLIT distance="150" swimtime="00:01:41.23" />
                    <SPLIT distance="200" swimtime="00:02:18.97" />
                    <SPLIT distance="250" swimtime="00:02:57.38" />
                    <SPLIT distance="300" swimtime="00:03:35.96" />
                    <SPLIT distance="350" swimtime="00:04:14.49" />
                    <SPLIT distance="400" swimtime="00:04:54.10" />
                    <SPLIT distance="450" swimtime="00:05:33.43" />
                    <SPLIT distance="500" swimtime="00:06:13.03" />
                    <SPLIT distance="550" swimtime="00:06:53.05" />
                    <SPLIT distance="600" swimtime="00:07:33.36" />
                    <SPLIT distance="650" swimtime="00:08:12.94" />
                    <SPLIT distance="700" swimtime="00:08:52.12" />
                    <SPLIT distance="750" swimtime="00:09:30.67" />
                    <SPLIT distance="800" swimtime="00:10:09.62" />
                    <SPLIT distance="850" swimtime="00:10:48.48" />
                    <SPLIT distance="900" swimtime="00:11:27.56" />
                    <SPLIT distance="950" swimtime="00:12:07.99" />
                    <SPLIT distance="1000" swimtime="00:12:47.45" />
                    <SPLIT distance="1050" swimtime="00:13:26.01" />
                    <SPLIT distance="1100" swimtime="00:14:04.99" />
                    <SPLIT distance="1150" swimtime="00:14:44.27" />
                    <SPLIT distance="1200" swimtime="00:15:23.95" />
                    <SPLIT distance="1250" swimtime="00:16:03.38" />
                    <SPLIT distance="1300" swimtime="00:16:42.10" />
                    <SPLIT distance="1350" swimtime="00:17:19.67" />
                    <SPLIT distance="1400" swimtime="00:17:59.28" />
                    <SPLIT distance="1450" swimtime="00:18:38.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11303" nation="BRA" region="PR" clubid="1518" swrid="93760" name="Associação De Talentos Da Natação" shortname="Atn/Curitiba">
          <ATHLETES>
            <ATHLETE firstname="Felipe" lastname="Bortoleto" birthdate="2008-09-05" gender="M" nation="BRA" license="406709" athleteid="1648" externalid="406709">
              <RESULTS>
                <RESULT eventid="1200" points="281" reactiontime="+81" swimtime="00:01:13.73" resultid="1649" heatid="3528" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1184" points="327" swimtime="00:00:31.54" resultid="1650" heatid="3518" lane="5" />
                <RESULT eventid="1296" points="339" swimtime="00:01:08.50" resultid="1651" heatid="3598" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="390" swimtime="00:01:01.35" resultid="1652" heatid="3573" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jhon" lastname="Caleb Dos Santos" birthdate="2010-03-02" gender="M" nation="BRA" license="359020" swrid="5588574" athleteid="1563" externalid="359020">
              <RESULTS>
                <RESULT eventid="1200" points="359" reactiontime="+73" swimtime="00:01:07.94" resultid="1564" heatid="3528" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1168" points="367" swimtime="00:01:17.16" resultid="1565" heatid="3511" lane="5" entrytime="00:01:21.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1152" points="446" swimtime="00:04:37.69" resultid="1566" heatid="3497" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.75" />
                    <SPLIT distance="100" swimtime="00:01:03.26" />
                    <SPLIT distance="150" swimtime="00:01:38.27" />
                    <SPLIT distance="200" swimtime="00:02:14.08" />
                    <SPLIT distance="250" swimtime="00:02:49.07" />
                    <SPLIT distance="300" swimtime="00:03:25.41" />
                    <SPLIT distance="350" swimtime="00:04:02.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1232" points="419" swimtime="00:02:26.44" resultid="1567" heatid="3560" lane="3" entrytime="00:02:32.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.87" />
                    <SPLIT distance="100" swimtime="00:01:05.35" />
                    <SPLIT distance="150" swimtime="00:01:50.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1296" points="401" swimtime="00:01:04.79" resultid="1568" heatid="3601" lane="6" entrytime="00:01:08.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yohanna" lastname="Vitoria Sousa" birthdate="2012-01-20" gender="F" nation="BRA" license="406710" athleteid="1653" externalid="406710">
              <RESULTS>
                <RESULT eventid="1074" points="86" reactiontime="+80" swimtime="00:00:57.15" resultid="1654" heatid="3405" lane="3" />
                <RESULT eventid="1138" points="133" swimtime="00:00:44.91" resultid="1655" heatid="3476" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Zaleski Dallazem" birthdate="2009-05-16" gender="M" nation="BRA" license="344286" swrid="5600280" athleteid="1553" externalid="344286" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1168" points="387" swimtime="00:01:15.81" resultid="1554" heatid="3512" lane="8" entrytime="00:01:20.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="377" swimtime="00:00:27.90" resultid="1555" heatid="3547" lane="7" entrytime="00:00:28.69" entrycourse="SCM" />
                <RESULT eventid="1312" points="385" swimtime="00:00:34.28" resultid="1556" heatid="3611" lane="1" entrytime="00:00:38.81" entrycourse="SCM" />
                <RESULT eventid="1248" points="399" swimtime="00:01:00.87" resultid="1557" heatid="3572" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Guedes Braga" birthdate="2013-04-09" gender="F" nation="BRA" license="385009" swrid="5602534" athleteid="1584" externalid="385009">
              <RESULTS>
                <RESULT eventid="1086" points="220" swimtime="00:03:02.50" resultid="1585" heatid="3427" lane="7" entrytime="00:02:57.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:01:27.15" />
                    <SPLIT distance="150" swimtime="00:02:16.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="211" reactiontime="+77" swimtime="00:00:42.39" resultid="1586" heatid="3405" lane="5" />
                <RESULT eventid="1102" points="186" swimtime="00:01:38.97" resultid="1587" heatid="3446" lane="4" entrytime="00:01:53.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="264" swimtime="00:00:35.70" resultid="1588" heatid="3480" lane="6" entrytime="00:00:35.85" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Kerppers Kreia" birthdate="2006-12-01" gender="M" nation="BRA" license="366815" swrid="5600195" athleteid="1538" externalid="366815">
              <RESULTS>
                <RESULT eventid="1184" points="368" swimtime="00:00:30.33" resultid="1539" heatid="3519" lane="2" />
                <RESULT eventid="1216" points="425" swimtime="00:00:26.81" resultid="1540" heatid="3548" lane="3" entrytime="00:00:27.33" entrycourse="SCM" />
                <RESULT eventid="1248" points="464" swimtime="00:00:57.90" resultid="1541" heatid="3579" lane="6" entrytime="00:00:59.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Leal Kuss" birthdate="2012-10-20" gender="M" nation="BRA" license="385085" swrid="5588768" athleteid="1589" externalid="385085">
              <RESULTS>
                <RESULT eventid="1077" points="119" reactiontime="+76" swimtime="00:00:44.85" resultid="1590" heatid="3413" lane="5" entrytime="00:00:50.94" entrycourse="SCM" />
                <RESULT eventid="1105" points="130" swimtime="00:01:37.18" resultid="1591" heatid="3448" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="169" swimtime="00:00:36.40" resultid="1592" heatid="3486" lane="6" entrytime="00:00:35.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Castellano Purkot" birthdate="2010-01-25" gender="M" nation="BRA" license="392484" swrid="5622268" athleteid="1628" externalid="392484">
              <RESULTS>
                <RESULT eventid="1216" points="308" swimtime="00:00:29.84" resultid="1629" heatid="3545" lane="5" entrytime="00:00:30.84" entrycourse="SCM" />
                <RESULT eventid="1280" points="217" reactiontime="+71" swimtime="00:00:36.79" resultid="1630" heatid="3590" lane="6" />
                <RESULT eventid="1248" points="282" swimtime="00:01:08.33" resultid="1631" heatid="3576" lane="3" entrytime="00:01:11.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Navarro Silva" birthdate="2011-01-10" gender="F" nation="BRA" license="406711" athleteid="1656" externalid="406711">
              <RESULTS>
                <RESULT eventid="1208" points="253" swimtime="00:00:36.24" resultid="1657" heatid="3533" lane="1" />
                <RESULT eventid="1192" points="240" reactiontime="+86" swimtime="00:01:28.30" resultid="1658" heatid="3523" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="251" reactiontime="+66" swimtime="00:00:40.01" resultid="1659" heatid="3586" lane="5" />
                <RESULT eventid="1240" points="252" swimtime="00:01:19.48" resultid="1660" heatid="3564" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Goncalves Ghion" birthdate="2014-10-15" gender="F" nation="BRA" license="406912" athleteid="1664" externalid="406912">
              <RESULTS>
                <RESULT eventid="1068" points="91" swimtime="00:01:02.99" resultid="1665" heatid="3400" lane="8" />
                <RESULT eventid="1128" points="92" swimtime="00:00:50.77" resultid="1666" heatid="3465" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Muller" birthdate="2009-10-10" gender="F" nation="BRA" license="376952" swrid="5600221" athleteid="1574" externalid="376952">
              <RESULTS>
                <RESULT eventid="1208" points="381" swimtime="00:00:31.61" resultid="1575" heatid="3538" lane="2" entrytime="00:00:31.23" entrycourse="SCM" />
                <RESULT eventid="1160" points="442" swimtime="00:01:21.82" resultid="1576" heatid="3506" lane="8" entrytime="00:01:21.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="352" swimtime="00:02:52.48" resultid="1577" heatid="3552" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                    <SPLIT distance="100" swimtime="00:01:27.49" />
                    <SPLIT distance="150" swimtime="00:02:13.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="435" swimtime="00:00:37.42" resultid="1578" heatid="3606" lane="3" entrytime="00:00:37.75" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelo" lastname="Correia Bonfim" birthdate="2009-06-21" gender="M" nation="BRA" license="391663" swrid="5622271" athleteid="1623" externalid="391663">
              <RESULTS>
                <RESULT eventid="1168" points="311" swimtime="00:01:21.52" resultid="1624" heatid="3511" lane="1" entrytime="00:01:26.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="361" swimtime="00:00:28.31" resultid="1625" heatid="3546" lane="6" entrytime="00:00:29.43" entrycourse="SCM" />
                <RESULT eventid="1280" points="274" reactiontime="+50" swimtime="00:00:34.02" resultid="1626" heatid="3591" lane="2" />
                <RESULT eventid="1248" points="381" swimtime="00:01:01.81" resultid="1627" heatid="3573" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Manuela Souza" birthdate="2016-07-07" gender="F" nation="BRA" license="406759" athleteid="1661" externalid="406759">
              <RESULTS>
                <RESULT eventid="1114" points="66" swimtime="00:00:29.32" resultid="1662" heatid="3460" lane="4" />
                <RESULT eventid="1134" points="62" swimtime="00:00:26.31" resultid="1663" heatid="3475" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="James" lastname="Roberto Zoschke" birthdate="1976-02-08" gender="M" nation="BRA" license="312251" swrid="5688617" athleteid="1546" externalid="312251">
              <RESULTS>
                <RESULT eventid="1168" points="459" swimtime="00:01:11.62" resultid="1547" heatid="3513" lane="8" entrytime="00:01:11.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="469" swimtime="00:00:32.10" resultid="1548" heatid="3611" lane="3" entrytime="00:00:33.77" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Camila" lastname="Duarte De Almeida" birthdate="2009-11-26" gender="F" nation="BRA" license="378819" swrid="5600152" athleteid="1579" externalid="378819">
              <RESULTS>
                <RESULT eventid="1208" points="427" swimtime="00:00:30.44" resultid="1580" heatid="3538" lane="3" entrytime="00:00:30.75" entrycourse="SCM" />
                <RESULT eventid="1176" points="359" swimtime="00:00:34.28" resultid="1581" heatid="3516" lane="2" entrytime="00:00:37.40" entrycourse="SCM" />
                <RESULT eventid="1304" points="295" swimtime="00:00:42.60" resultid="1582" heatid="3604" lane="4" />
                <RESULT eventid="1240" points="409" swimtime="00:01:07.69" resultid="1583" heatid="3569" lane="8" entrytime="00:01:07.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Faria Del Valle" birthdate="2009-08-28" gender="M" nation="BRA" license="376328" swrid="5600155" athleteid="1569" externalid="376328">
              <RESULTS>
                <RESULT eventid="1216" points="513" swimtime="00:00:25.18" resultid="1570" heatid="3548" lane="1" entrytime="00:00:27.69" entrycourse="SCM" />
                <RESULT eventid="1312" points="430" swimtime="00:00:33.04" resultid="1571" heatid="3611" lane="7" entrytime="00:00:37.88" entrycourse="SCM" />
                <RESULT eventid="1280" points="351" reactiontime="+49" swimtime="00:00:31.32" resultid="1572" heatid="3591" lane="3" />
                <RESULT eventid="1248" points="475" swimtime="00:00:57.44" resultid="1573" heatid="3579" lane="5" entrytime="00:00:59.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Sofia Silva" birthdate="2007-05-28" gender="F" nation="BRA" license="390921" swrid="5600260" athleteid="1608" externalid="390921">
              <RESULTS>
                <RESULT eventid="1208" points="215" swimtime="00:00:38.27" resultid="1609" heatid="3535" lane="7" entrytime="00:00:39.92" entrycourse="SCM" />
                <RESULT eventid="1176" points="167" swimtime="00:00:44.22" resultid="1610" heatid="3514" lane="5" />
                <RESULT eventid="1160" points="225" swimtime="00:01:42.52" resultid="1611" heatid="3503" lane="3" entrytime="00:01:54.26" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="217" swimtime="00:03:22.76" resultid="1612" heatid="3553" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.19" />
                    <SPLIT distance="100" swimtime="00:01:38.64" />
                    <SPLIT distance="150" swimtime="00:02:36.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="200" swimtime="00:00:48.46" resultid="1613" heatid="3605" lane="6" entrytime="00:00:50.15" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Vinicius Zonta" birthdate="2012-11-14" gender="M" nation="BRA" license="399517" swrid="5652903" athleteid="1644" externalid="399517">
              <RESULTS>
                <RESULT eventid="1089" status="DSQ" swimtime="00:02:41.08" resultid="1645" heatid="3433" lane="2" entrytime="00:02:53.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.88" />
                    <SPLIT distance="100" swimtime="00:01:15.13" />
                    <SPLIT distance="150" swimtime="00:01:58.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="173" swimtime="00:01:28.28" resultid="1646" heatid="3450" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="234" swimtime="00:00:32.70" resultid="1647" heatid="3486" lane="7" entrytime="00:00:36.14" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mauricio" lastname="Furtado Niwa" birthdate="1978-05-30" gender="M" nation="BRA" license="398757" swrid="5653291" athleteid="1549" externalid="398757">
              <RESULTS>
                <RESULT eventid="1184" points="493" swimtime="00:00:27.52" resultid="1550" heatid="3522" lane="3" entrytime="00:00:28.09" entrycourse="SCM" />
                <RESULT eventid="1216" points="461" swimtime="00:00:26.08" resultid="1551" heatid="3542" lane="8" />
                <RESULT eventid="1296" points="483" swimtime="00:01:00.87" resultid="1552" heatid="3602" lane="2" entrytime="00:01:01.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Kerniski Demantova" birthdate="1982-05-25" gender="M" nation="BRA" license="398222" swrid="5653293" athleteid="1542" externalid="398222">
              <RESULTS>
                <RESULT eventid="1184" points="361" swimtime="00:00:30.54" resultid="1543" heatid="3519" lane="4" />
                <RESULT eventid="1152" points="403" swimtime="00:04:47.34" resultid="1544" heatid="3500" lane="6" entrytime="00:04:52.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:09.07" />
                    <SPLIT distance="150" swimtime="00:01:45.70" />
                    <SPLIT distance="200" swimtime="00:02:22.65" />
                    <SPLIT distance="250" swimtime="00:02:59.39" />
                    <SPLIT distance="300" swimtime="00:03:35.84" />
                    <SPLIT distance="350" swimtime="00:04:12.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1264" points="319" swimtime="00:20:38.41" resultid="1545" heatid="3585" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:14.87" />
                    <SPLIT distance="150" swimtime="00:01:54.69" />
                    <SPLIT distance="200" swimtime="00:02:34.73" />
                    <SPLIT distance="250" swimtime="00:03:15.23" />
                    <SPLIT distance="300" swimtime="00:03:55.60" />
                    <SPLIT distance="350" swimtime="00:04:35.99" />
                    <SPLIT distance="400" swimtime="00:05:16.36" />
                    <SPLIT distance="450" swimtime="00:05:56.85" />
                    <SPLIT distance="500" swimtime="00:06:37.72" />
                    <SPLIT distance="550" swimtime="00:07:18.85" />
                    <SPLIT distance="600" swimtime="00:07:59.74" />
                    <SPLIT distance="650" swimtime="00:08:40.57" />
                    <SPLIT distance="700" swimtime="00:09:21.83" />
                    <SPLIT distance="750" swimtime="00:10:03.25" />
                    <SPLIT distance="800" swimtime="00:10:45.37" />
                    <SPLIT distance="850" swimtime="00:11:27.10" />
                    <SPLIT distance="900" swimtime="00:12:09.65" />
                    <SPLIT distance="950" swimtime="00:12:51.65" />
                    <SPLIT distance="1000" swimtime="00:13:34.26" />
                    <SPLIT distance="1050" swimtime="00:14:16.26" />
                    <SPLIT distance="1100" swimtime="00:14:58.90" />
                    <SPLIT distance="1150" swimtime="00:15:41.60" />
                    <SPLIT distance="1200" swimtime="00:16:24.77" />
                    <SPLIT distance="1250" swimtime="00:17:08.26" />
                    <SPLIT distance="1300" swimtime="00:17:50.90" />
                    <SPLIT distance="1350" swimtime="00:18:33.14" />
                    <SPLIT distance="1400" swimtime="00:19:15.71" />
                    <SPLIT distance="1450" swimtime="00:19:57.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Neves Vianna" birthdate="2007-12-30" gender="F" nation="BRA" license="391106" swrid="5600223" athleteid="1614" externalid="391106">
              <RESULTS>
                <RESULT eventid="1144" points="228" swimtime="00:06:18.35" resultid="1615" heatid="3491" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.28" />
                    <SPLIT distance="100" swimtime="00:01:25.10" />
                    <SPLIT distance="150" swimtime="00:02:12.81" />
                    <SPLIT distance="200" swimtime="00:03:01.42" />
                    <SPLIT distance="250" swimtime="00:03:50.51" />
                    <SPLIT distance="300" swimtime="00:04:40.54" />
                    <SPLIT distance="350" swimtime="00:05:30.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1192" points="213" reactiontime="+70" swimtime="00:01:31.83" resultid="1616" heatid="3525" lane="7" entrytime="00:01:33.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="197" reactiontime="+50" swimtime="00:00:43.38" resultid="1617" heatid="3588" lane="1" entrytime="00:00:43.62" entrycourse="SCM" />
                <RESULT eventid="1240" points="223" swimtime="00:01:22.85" resultid="1618" heatid="3565" lane="6" entrytime="00:01:22.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Garcia De Fraga" birthdate="2009-03-24" gender="M" nation="BRA" license="342147" swrid="5600172" athleteid="1523" externalid="342147" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1200" points="546" reactiontime="+61" swimtime="00:00:59.12" resultid="1524" heatid="3532" lane="5" entrytime="00:01:01.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="508" swimtime="00:00:25.26" resultid="1525" heatid="3543" lane="4" />
                <RESULT eventid="1232" points="574" swimtime="00:02:11.91" resultid="1526" heatid="3561" lane="6" entrytime="00:02:15.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.99" />
                    <SPLIT distance="100" swimtime="00:01:00.56" />
                    <SPLIT distance="150" swimtime="00:01:38.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="542" swimtime="00:00:54.97" resultid="1527" heatid="3574" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Riccieri" lastname="Rodrigues Muzolon" birthdate="2010-11-08" gender="M" nation="BRA" license="385439" swrid="5588887" athleteid="1593" externalid="385439">
              <RESULTS>
                <RESULT eventid="1184" status="DNS" swimtime="00:00:00.00" resultid="1594" heatid="3521" lane="1" entrytime="00:00:37.68" entrycourse="SCM" />
                <RESULT eventid="1168" status="DNS" swimtime="00:00:00.00" resultid="1595" heatid="3510" lane="5" entrytime="00:01:27.32" entrycourse="SCM" />
                <RESULT eventid="1152" status="DNS" swimtime="00:00:00.00" resultid="1596" heatid="3496" lane="4" />
                <RESULT eventid="1312" status="DNS" swimtime="00:00:00.00" resultid="1597" heatid="3610" lane="5" entrytime="00:00:41.60" entrycourse="SCM" />
                <RESULT eventid="1248" status="DNS" swimtime="00:00:00.00" resultid="1598" heatid="3574" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcos" lastname="Demchuk" birthdate="2011-06-15" gender="M" nation="BRA" license="388540" swrid="5602530" athleteid="1604" externalid="388540">
              <RESULTS>
                <RESULT eventid="1168" points="183" swimtime="00:01:37.32" resultid="1605" heatid="3509" lane="5" entrytime="00:01:59.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="221" swimtime="00:00:33.33" resultid="1606" heatid="3544" lane="5" entrytime="00:00:34.51" entrycourse="SCM" />
                <RESULT eventid="1312" points="172" swimtime="00:00:44.85" resultid="1607" heatid="3610" lane="2" entrytime="00:00:48.81" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Yuji Yamazato" birthdate="2008-10-01" gender="M" nation="BRA" license="392664" swrid="5622313" athleteid="1632" externalid="392664">
              <RESULTS>
                <RESULT eventid="1184" points="304" swimtime="00:00:32.34" resultid="1633" heatid="3517" lane="2" />
                <RESULT eventid="1216" points="344" swimtime="00:00:28.77" resultid="1634" heatid="3547" lane="8" entrytime="00:00:28.82" entrycourse="SCM" />
                <RESULT eventid="1296" status="DNS" swimtime="00:00:00.00" resultid="1635" heatid="3599" lane="7" />
                <RESULT eventid="1248" status="DNS" swimtime="00:00:00.00" resultid="1636" heatid="3577" lane="6" entrytime="00:01:07.19" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Fonseca Vendramin" birthdate="2008-09-28" gender="F" nation="BRA" license="393918" swrid="5622282" athleteid="1637" externalid="393918">
              <RESULTS>
                <RESULT eventid="1288" points="269" swimtime="00:01:23.63" resultid="1638" heatid="3595" lane="6" entrytime="00:01:25.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="348" swimtime="00:01:11.44" resultid="1639" heatid="3566" lane="6" entrytime="00:01:14.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Bordignon Becker" birthdate="2011-12-31" gender="M" nation="BRA" license="391107" swrid="5602516" athleteid="1619" externalid="391107">
              <RESULTS>
                <RESULT eventid="1216" points="167" swimtime="00:00:36.59" resultid="1620" heatid="3544" lane="7" entrytime="00:00:39.78" entrycourse="SCM" />
                <RESULT eventid="1280" points="94" reactiontime="+69" swimtime="00:00:48.50" resultid="1621" heatid="3592" lane="6" entrytime="00:00:49.72" entrycourse="SCM" />
                <RESULT eventid="1248" points="155" swimtime="00:01:23.35" resultid="1622" heatid="3575" lane="7" entrytime="00:01:29.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Garcia Fraga" birthdate="2003-10-07" gender="M" nation="BRA" license="283467" athleteid="1531" externalid="283467" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1216" points="490" swimtime="00:00:25.57" resultid="1532" heatid="3543" lane="1" />
                <RESULT eventid="1232" points="522" swimtime="00:02:16.15" resultid="1533" heatid="3558" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="100" swimtime="00:01:03.95" />
                    <SPLIT distance="150" swimtime="00:01:43.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Ocanha" birthdate="2005-06-21" gender="M" nation="BRA" license="313769" swrid="5600231" athleteid="1528" externalid="313769" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1216" points="556" swimtime="00:00:24.51" resultid="1529" heatid="3550" lane="3" entrytime="00:00:24.41" entrycourse="SCM" />
                <RESULT eventid="1312" points="555" swimtime="00:00:30.35" resultid="1530" heatid="3612" lane="3" entrytime="00:00:30.42" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isis" lastname="De Miranda" birthdate="2012-01-10" gender="F" nation="BRA" license="397278" swrid="5652886" athleteid="1640" externalid="397278">
              <RESULTS>
                <RESULT eventid="1086" points="280" swimtime="00:02:48.61" resultid="1641" heatid="3427" lane="8" entrytime="00:03:02.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:20.57" />
                    <SPLIT distance="150" swimtime="00:02:04.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1118" points="194" swimtime="00:01:33.21" resultid="1642" heatid="3462" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="249" swimtime="00:00:36.44" resultid="1643" heatid="3480" lane="8" entrytime="00:00:39.13" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Freitas Szucs" birthdate="2011-10-02" gender="M" nation="BRA" license="377272" swrid="5588708" athleteid="1558" externalid="377272">
              <RESULTS>
                <RESULT eventid="1184" points="155" swimtime="00:00:40.48" resultid="1559" heatid="3520" lane="5" entrytime="00:00:42.65" entrycourse="SCM" />
                <RESULT eventid="1216" points="185" swimtime="00:00:35.33" resultid="1560" heatid="3544" lane="6" entrytime="00:00:36.81" entrycourse="SCM" />
                <RESULT eventid="1312" status="DSQ" swimtime="00:00:48.07" resultid="1561" heatid="3610" lane="7" entrytime="00:00:51.59" entrycourse="SCM" />
                <RESULT eventid="1248" points="185" swimtime="00:01:18.60" resultid="1562" heatid="3575" lane="6" entrytime="00:01:21.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Angelo" lastname="De Queiroz Neto" birthdate="2003-10-31" gender="M" nation="BRA" license="342814" swrid="5600149" athleteid="1534" externalid="342814" level="AERC">
              <RESULTS>
                <RESULT eventid="1184" points="385" swimtime="00:00:29.88" resultid="1535" heatid="3522" lane="1" entrytime="00:00:29.44" entrycourse="SCM" />
                <RESULT eventid="1296" points="380" swimtime="00:01:05.91" resultid="1536" heatid="3601" lane="3" entrytime="00:01:05.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1248" points="412" swimtime="00:01:00.26" resultid="1537" heatid="3579" lane="3" entrytime="00:00:59.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Duarte De Almeida" birthdate="2013-12-09" gender="M" nation="BRA" license="385711" swrid="5588666" athleteid="1599" externalid="385711">
              <RESULTS>
                <RESULT eventid="1089" points="202" swimtime="00:02:49.26" resultid="1600" heatid="3432" lane="4" entrytime="00:02:56.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                    <SPLIT distance="100" swimtime="00:01:22.66" />
                    <SPLIT distance="150" swimtime="00:02:08.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="168" swimtime="00:01:39.99" resultid="1601" heatid="3397" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="190" swimtime="00:01:25.69" resultid="1602" heatid="3451" lane="2" entrytime="00:01:35.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="222" swimtime="00:00:33.26" resultid="1603" heatid="3486" lane="4" entrytime="00:00:34.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabiana" lastname="Zaleski Dallazem" birthdate="2009-05-16" gender="F" nation="BRA" license="344287" swrid="5600279" athleteid="1519" externalid="344287" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1208" points="450" swimtime="00:00:29.92" resultid="1520" heatid="3538" lane="4" entrytime="00:00:30.34" entrycourse="SCM" />
                <RESULT eventid="1192" points="466" reactiontime="+68" swimtime="00:01:10.76" resultid="1521" heatid="3527" lane="3" entrytime="00:01:09.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1272" points="471" reactiontime="+65" swimtime="00:00:32.44" resultid="1522" heatid="3589" lane="3" entrytime="00:00:32.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2539" nation="BRA" region="PR" clubid="1667" swrid="93771" name="Círculo Militar Do Paraná" shortname="Círculo Militar">
          <ATHLETES>
            <ATHLETE firstname="Bruno" lastname="Yamamoto" birthdate="2006-04-22" gender="M" nation="BRA" license="336569" athleteid="1699" externalid="336569">
              <RESULTS>
                <RESULT eventid="1184" points="346" swimtime="00:00:30.96" resultid="1700" heatid="3519" lane="8" />
                <RESULT eventid="1216" points="396" swimtime="00:00:27.44" resultid="1701" heatid="3541" lane="8" />
                <RESULT eventid="1248" points="377" swimtime="00:01:02.07" resultid="1702" heatid="3571" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Oliveira Martini" birthdate="2008-10-31" gender="M" nation="BRA" license="406953" athleteid="1720" externalid="406953">
              <RESULTS>
                <RESULT eventid="1152" points="255" swimtime="00:05:34.39" resultid="1721" heatid="3497" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.67" />
                    <SPLIT distance="100" swimtime="00:01:17.38" />
                    <SPLIT distance="150" swimtime="00:02:00.70" />
                    <SPLIT distance="200" swimtime="00:02:45.37" />
                    <SPLIT distance="250" swimtime="00:03:30.01" />
                    <SPLIT distance="300" swimtime="00:04:14.13" />
                    <SPLIT distance="350" swimtime="00:04:57.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="365" swimtime="00:00:28.19" resultid="1722" heatid="3540" lane="3" />
                <RESULT eventid="1248" points="328" swimtime="00:01:04.96" resultid="1723" heatid="3573" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vicente" lastname="Bileski" birthdate="2011-06-29" gender="M" nation="BRA" license="406950" athleteid="1710" externalid="406950">
              <RESULTS>
                <RESULT eventid="1216" points="153" swimtime="00:00:37.67" resultid="1711" heatid="3543" lane="5" />
                <RESULT eventid="1312" points="141" swimtime="00:00:47.91" resultid="1712" heatid="3607" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="De Queiroz" birthdate="2007-08-20" gender="M" nation="BRA" license="406949" athleteid="1707" externalid="406949">
              <RESULTS>
                <RESULT eventid="1184" points="197" swimtime="00:00:37.33" resultid="1708" heatid="3517" lane="7" />
                <RESULT eventid="1248" points="179" swimtime="00:01:19.55" resultid="1709" heatid="3574" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernando" lastname="Jun Melo Ogima" birthdate="2006-07-05" gender="M" nation="BRA" license="378332" swrid="5622284" athleteid="1672" externalid="378332">
              <RESULTS>
                <RESULT eventid="1184" points="363" swimtime="00:00:30.48" resultid="1673" heatid="3521" lane="2" entrytime="00:00:32.22" entrycourse="SCM" />
                <RESULT eventid="1216" points="392" swimtime="00:00:27.54" resultid="1674" heatid="3542" lane="2" />
                <RESULT eventid="1232" points="291" swimtime="00:02:45.27" resultid="1675" heatid="3557" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                    <SPLIT distance="100" swimtime="00:01:16.16" />
                    <SPLIT distance="150" swimtime="00:02:05.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="335" swimtime="00:00:35.92" resultid="1676" heatid="3611" lane="8" entrytime="00:00:39.12" entrycourse="SCM" />
                <RESULT eventid="1280" points="281" swimtime="00:00:33.73" resultid="1677" heatid="3592" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thomas" lastname="Gomes" birthdate="2009-06-15" gender="M" nation="BRA" license="406948" athleteid="1703" externalid="406948">
              <RESULTS>
                <RESULT eventid="1312" points="128" swimtime="00:00:49.43" resultid="1704" heatid="3609" lane="3" />
                <RESULT eventid="1280" points="124" reactiontime="+50" swimtime="00:00:44.32" resultid="1705" heatid="3592" lane="1" />
                <RESULT eventid="1248" points="154" swimtime="00:01:23.61" resultid="1706" heatid="3575" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Cavalcante Pierin" birthdate="2012-10-30" gender="F" nation="BRA" license="406952" athleteid="1716" externalid="406952">
              <RESULTS>
                <RESULT eventid="1074" status="DSQ" swimtime="00:00:44.16" resultid="1717" heatid="3407" lane="3" />
                <RESULT eventid="1102" points="174" swimtime="00:01:41.03" resultid="1718" heatid="3445" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1138" points="228" swimtime="00:00:37.52" resultid="1719" heatid="3477" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Vieira Coelho" birthdate="2014-09-28" gender="F" nation="BRA" license="406951" athleteid="1713" externalid="406951">
              <RESULTS>
                <RESULT eventid="1068" points="111" swimtime="00:00:58.90" resultid="1714" heatid="3399" lane="4" />
                <RESULT eventid="1128" points="97" swimtime="00:00:49.84" resultid="1715" heatid="3466" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Cavalcante Pierin" birthdate="2010-12-28" gender="M" nation="BRA" license="391227" swrid="5622269" athleteid="1688" externalid="391227">
              <RESULTS>
                <RESULT eventid="1184" status="DNS" swimtime="00:00:00.00" resultid="1689" heatid="3520" lane="3" />
                <RESULT eventid="1152" points="217" swimtime="00:05:53.02" resultid="1690" heatid="3497" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                    <SPLIT distance="100" swimtime="00:01:20.93" />
                    <SPLIT distance="150" swimtime="00:02:07.30" />
                    <SPLIT distance="200" swimtime="00:02:53.89" />
                    <SPLIT distance="250" swimtime="00:03:40.04" />
                    <SPLIT distance="300" swimtime="00:04:27.05" />
                    <SPLIT distance="350" swimtime="00:05:11.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="142" swimtime="00:00:47.77" resultid="1691" heatid="3607" lane="2" />
                <RESULT eventid="1280" points="173" reactiontime="+66" swimtime="00:00:39.67" resultid="1692" heatid="3591" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Torres Oliveira" birthdate="2008-04-10" gender="M" nation="BRA" license="400274" swrid="5653303" athleteid="1693" externalid="400274">
              <RESULTS>
                <RESULT eventid="1168" points="255" swimtime="00:01:27.13" resultid="1694" heatid="3508" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="327" swimtime="00:00:29.24" resultid="1695" heatid="3541" lane="6" />
                <RESULT eventid="1312" points="297" swimtime="00:00:37.39" resultid="1696" heatid="3607" lane="4" />
                <RESULT eventid="1280" points="218" reactiontime="+61" swimtime="00:00:36.71" resultid="1697" heatid="3591" lane="7" />
                <RESULT eventid="1248" points="290" swimtime="00:01:07.68" resultid="1698" heatid="3573" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Maria Romanelli" birthdate="2011-04-18" gender="F" nation="BRA" license="378335" swrid="5588803" athleteid="1678" externalid="378335">
              <RESULTS>
                <RESULT eventid="1208" points="356" swimtime="00:00:32.35" resultid="1679" heatid="3537" lane="8" entrytime="00:00:33.74" entrycourse="SCM" />
                <RESULT eventid="1304" points="213" swimtime="00:00:47.46" resultid="1680" heatid="3605" lane="3" entrytime="00:00:48.52" entrycourse="SCM" />
                <RESULT eventid="1272" points="249" reactiontime="+77" swimtime="00:00:40.11" resultid="1681" heatid="3588" lane="2" entrytime="00:00:40.89" entrycourse="SCM" />
                <RESULT eventid="1240" points="369" swimtime="00:01:10.00" resultid="1682" heatid="3567" lane="7" entrytime="00:01:12.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Vieira De Macedo Brasil" birthdate="2009-12-19" gender="F" nation="BRA" license="344143" swrid="5622311" athleteid="1668" externalid="344143">
              <RESULTS>
                <RESULT eventid="1144" points="314" swimtime="00:05:40.28" resultid="1669" heatid="3492" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.49" />
                    <SPLIT distance="100" swimtime="00:01:15.19" />
                    <SPLIT distance="150" swimtime="00:01:58.12" />
                    <SPLIT distance="200" swimtime="00:02:41.34" />
                    <SPLIT distance="250" swimtime="00:03:26.33" />
                    <SPLIT distance="300" swimtime="00:04:12.10" />
                    <SPLIT distance="350" swimtime="00:04:58.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="364" swimtime="00:00:32.11" resultid="1670" heatid="3534" lane="1" />
                <RESULT eventid="1304" points="297" swimtime="00:00:42.51" resultid="1671" heatid="3604" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Manocchio" birthdate="2011-07-28" gender="M" nation="BRA" license="384916" swrid="5588573" athleteid="1683" externalid="384916">
              <RESULTS>
                <RESULT eventid="1184" points="197" swimtime="00:00:37.33" resultid="1684" heatid="3520" lane="1" />
                <RESULT eventid="1152" points="318" swimtime="00:05:10.65" resultid="1685" heatid="3498" lane="4" entrytime="00:05:32.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                    <SPLIT distance="100" swimtime="00:01:10.48" />
                    <SPLIT distance="150" swimtime="00:01:50.53" />
                    <SPLIT distance="200" swimtime="00:02:32.45" />
                    <SPLIT distance="250" swimtime="00:03:12.20" />
                    <SPLIT distance="300" swimtime="00:03:52.86" />
                    <SPLIT distance="350" swimtime="00:04:33.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="315" swimtime="00:00:29.60" resultid="1686" heatid="3545" lane="8" entrytime="00:00:32.19" entrycourse="SCM" />
                <RESULT eventid="1248" points="315" swimtime="00:01:05.84" resultid="1687" heatid="3577" lane="1" entrytime="00:01:08.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="2773" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Ribeiro Melo" birthdate="2011-07-01" gender="F" nation="BRA" license="390923" swrid="5602577" athleteid="2801" externalid="390923">
              <RESULTS>
                <RESULT eventid="1208" points="369" swimtime="00:00:31.95" resultid="2802" heatid="3537" lane="6" entrytime="00:00:32.20" entrycourse="SCM" />
                <RESULT eventid="1160" points="274" swimtime="00:01:35.91" resultid="2803" heatid="3503" lane="5" entrytime="00:01:51.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" status="DSQ" swimtime="00:03:02.10" resultid="2804" heatid="3553" lane="2" entrytime="00:03:39.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.64" />
                    <SPLIT distance="100" swimtime="00:01:30.91" />
                    <SPLIT distance="150" swimtime="00:02:23.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1304" points="293" swimtime="00:00:42.69" resultid="2805" heatid="3605" lane="4" entrytime="00:00:44.16" entrycourse="SCM" />
                <RESULT eventid="1240" points="339" swimtime="00:01:12.05" resultid="2806" heatid="3566" lane="4" entrytime="00:01:13.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Schneider Yazbek" birthdate="2013-03-07" gender="F" nation="BRA" license="378329" swrid="5588907" athleteid="2780" externalid="378329">
              <RESULTS>
                <RESULT eventid="1086" points="321" swimtime="00:02:41.08" resultid="2781" heatid="3428" lane="7" entrytime="00:02:44.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                    <SPLIT distance="100" swimtime="00:01:18.10" />
                    <SPLIT distance="150" swimtime="00:02:00.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="217" swimtime="00:00:41.99" resultid="2782" heatid="3409" lane="3" entrytime="00:00:45.83" entrycourse="SCM" />
                <RESULT eventid="1102" points="267" swimtime="00:01:27.72" resultid="2783" heatid="3447" lane="4" entrytime="00:01:33.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1118" points="194" swimtime="00:01:33.25" resultid="2784" heatid="3462" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Zanatta Duda" birthdate="2013-08-28" gender="F" nation="BRA" license="406914" athleteid="2813" externalid="406914">
              <RESULTS>
                <RESULT eventid="1138" points="139" swimtime="00:00:44.22" resultid="2814" heatid="3477" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Ferreira Rais" birthdate="2007-07-04" gender="M" nation="BRA" license="398656" swrid="5697227" athleteid="2791" externalid="398656">
              <RESULTS>
                <RESULT eventid="1184" points="260" swimtime="00:00:34.07" resultid="2792" heatid="3521" lane="7" entrytime="00:00:35.68" entrycourse="SCM" />
                <RESULT eventid="1216" points="331" swimtime="00:00:29.14" resultid="2793" heatid="3546" lane="7" entrytime="00:00:30.20" entrycourse="SCM" />
                <RESULT eventid="1296" status="DNS" swimtime="00:00:00.00" resultid="2794" heatid="3597" lane="4" />
                <RESULT eventid="1280" points="202" reactiontime="+55" swimtime="00:00:37.66" resultid="2795" heatid="3592" lane="3" entrytime="00:00:39.44" entrycourse="SCM" />
                <RESULT eventid="1248" points="294" swimtime="00:01:07.43" resultid="2796" heatid="3575" lane="3" entrytime="00:01:19.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Paes Schemiko" birthdate="2013-02-25" gender="F" nation="BRA" license="406918" athleteid="2820" externalid="406918" />
            <ATHLETE firstname="Rodrigo" lastname="Zanatta Duda" birthdate="2011-09-12" gender="M" nation="BRA" license="406917" athleteid="2815" externalid="406917">
              <RESULTS>
                <RESULT eventid="1200" points="180" reactiontime="+82" swimtime="00:01:25.55" resultid="2816" heatid="3529" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="159" swimtime="00:00:37.14" resultid="2817" heatid="3543" lane="3" />
                <RESULT eventid="1280" points="177" reactiontime="+76" swimtime="00:00:39.35" resultid="2818" heatid="3590" lane="1" />
                <RESULT eventid="1248" points="136" swimtime="00:01:27.05" resultid="2819" heatid="3572" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Ribeiro Melo" birthdate="2013-02-25" gender="M" nation="BRA" license="406921" athleteid="2821" externalid="406921">
              <RESULTS>
                <RESULT eventid="1077" reactiontime="+72" status="DSQ" swimtime="00:00:52.09" resultid="2822" heatid="3413" lane="1" />
                <RESULT eventid="1065" points="88" swimtime="00:02:03.95" resultid="2823" heatid="3395" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="100" swimtime="00:01:45.96" resultid="2824" heatid="3450" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1141" points="134" swimtime="00:00:39.37" resultid="2825" heatid="3482" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aline" lastname="Hirano" birthdate="2007-11-13" gender="F" nation="BRA" license="358898" swrid="5622283" athleteid="2807" externalid="358898">
              <RESULTS>
                <RESULT eventid="1144" points="381" swimtime="00:05:19.02" resultid="2808" heatid="3490" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="100" swimtime="00:01:14.26" />
                    <SPLIT distance="150" swimtime="00:01:54.49" />
                    <SPLIT distance="200" swimtime="00:02:35.91" />
                    <SPLIT distance="250" swimtime="00:03:17.29" />
                    <SPLIT distance="300" swimtime="00:03:59.12" />
                    <SPLIT distance="350" swimtime="00:04:40.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="406" swimtime="00:00:30.96" resultid="2809" heatid="3533" lane="6" />
                <RESULT eventid="1192" points="360" reactiontime="+68" swimtime="00:01:17.16" resultid="2810" heatid="3525" lane="3" entrytime="00:01:24.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1224" points="325" swimtime="00:02:57.08" resultid="2811" heatid="3552" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                    <SPLIT distance="100" swimtime="00:01:25.19" />
                    <SPLIT distance="150" swimtime="00:02:18.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1256" points="357" swimtime="00:21:19.89" resultid="2812" heatid="3582" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:01:18.51" />
                    <SPLIT distance="150" swimtime="00:02:01.43" />
                    <SPLIT distance="200" swimtime="00:02:44.43" />
                    <SPLIT distance="250" swimtime="00:03:28.32" />
                    <SPLIT distance="300" swimtime="00:04:12.08" />
                    <SPLIT distance="350" swimtime="00:04:56.30" />
                    <SPLIT distance="400" swimtime="00:05:39.73" />
                    <SPLIT distance="450" swimtime="00:06:24.00" />
                    <SPLIT distance="500" swimtime="00:07:08.01" />
                    <SPLIT distance="550" swimtime="00:07:50.83" />
                    <SPLIT distance="600" swimtime="00:08:34.64" />
                    <SPLIT distance="650" swimtime="00:09:17.28" />
                    <SPLIT distance="700" swimtime="00:10:00.75" />
                    <SPLIT distance="750" swimtime="00:10:44.08" />
                    <SPLIT distance="800" swimtime="00:11:27.70" />
                    <SPLIT distance="850" swimtime="00:12:11.12" />
                    <SPLIT distance="900" swimtime="00:12:54.84" />
                    <SPLIT distance="950" swimtime="00:13:38.40" />
                    <SPLIT distance="1000" swimtime="00:14:22.48" />
                    <SPLIT distance="1050" swimtime="00:15:04.85" />
                    <SPLIT distance="1100" swimtime="00:15:47.63" />
                    <SPLIT distance="1150" swimtime="00:16:29.92" />
                    <SPLIT distance="1200" swimtime="00:17:13.40" />
                    <SPLIT distance="1250" swimtime="00:17:55.42" />
                    <SPLIT distance="1300" swimtime="00:18:37.57" />
                    <SPLIT distance="1350" swimtime="00:19:19.47" />
                    <SPLIT distance="1400" swimtime="00:20:01.46" />
                    <SPLIT distance="1450" swimtime="00:20:42.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jennifer" lastname="De Abreu" birthdate="2009-11-07" gender="F" nation="BRA" license="356212" swrid="5600144" athleteid="2774" externalid="356212">
              <RESULTS>
                <RESULT eventid="1144" points="479" swimtime="00:04:55.60" resultid="2775" heatid="3490" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.56" />
                    <SPLIT distance="100" swimtime="00:01:11.24" />
                    <SPLIT distance="150" swimtime="00:01:49.50" />
                    <SPLIT distance="200" swimtime="00:02:27.54" />
                    <SPLIT distance="250" swimtime="00:03:05.50" />
                    <SPLIT distance="300" swimtime="00:03:43.95" />
                    <SPLIT distance="350" swimtime="00:04:20.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="464" swimtime="00:00:29.61" resultid="2776" heatid="3539" lane="1" entrytime="00:00:30.18" entrycourse="SCM" />
                <RESULT eventid="1224" status="DSQ" swimtime="00:02:42.71" resultid="2777" heatid="3555" lane="4" entrytime="00:02:49.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.98" />
                    <SPLIT distance="100" swimtime="00:01:18.43" />
                    <SPLIT distance="150" swimtime="00:02:06.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1288" points="357" swimtime="00:01:16.17" resultid="2778" heatid="3594" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1240" points="487" swimtime="00:01:03.83" resultid="2779" heatid="3569" lane="6" entrytime="00:01:06.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Guilherme Ballatka" birthdate="2007-06-24" gender="M" nation="BRA" license="398616" swrid="5697228" athleteid="2785" externalid="398616">
              <RESULTS>
                <RESULT eventid="1200" points="315" reactiontime="+73" swimtime="00:01:10.99" resultid="2786" heatid="3529" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="408" swimtime="00:00:27.17" resultid="2787" heatid="3548" lane="6" entrytime="00:00:27.51" entrycourse="SCM" />
                <RESULT eventid="1312" status="DSQ" swimtime="00:00:38.56" resultid="2788" heatid="3610" lane="4" entrytime="00:00:39.18" entrycourse="SCM" />
                <RESULT eventid="1280" points="367" reactiontime="+64" swimtime="00:00:30.87" resultid="2789" heatid="3593" lane="7" entrytime="00:00:31.71" entrycourse="SCM" />
                <RESULT eventid="1248" points="401" swimtime="00:01:00.76" resultid="2790" heatid="3577" lane="8" entrytime="00:01:09.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Sprengel Betim" birthdate="2012-08-17" gender="F" nation="BRA" license="385011" swrid="5588922" athleteid="2797" externalid="385011">
              <RESULTS>
                <RESULT eventid="1062" points="143" swimtime="00:01:59.17" resultid="2798" heatid="3393" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1102" points="209" swimtime="00:01:35.21" resultid="2799" heatid="3444" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1118" points="145" swimtime="00:01:42.84" resultid="2800" heatid="3461" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
