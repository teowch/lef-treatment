<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.80168">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Curitiba" name="Torneio Regional da 1ª Região (Pré-Mirim/Petiz)" course="LCM" deadline="2024-08-12" entrystartdate="2024-08-06" entrytype="INVITATION" hostclub="Clube Curitibano" hostclub.url="https://clubecuritibano.com.br/" number="38314" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/newInterface/eventos/38314" startmethod="1" timing="AUTOMATIC" touchpad="ONESIDE" masters="F" withdrawuntil="2024-08-14" state="PR" nation="BRA" hytek.courseorder="L">
      <AGEDATE value="2024-01-01" type="YEAR" />
      <POOL name="Parque Aquático do Clube Curitibano" lanemin="1" lanemax="8" />
      <FACILITY city="Curitiba" name="Parque Aquático do Clube Curitibano" nation="BRA" state="PR" street="Avenida Presidente Getúlio Vargas, 2857" street2="Água Verde" zip="80240-040" />
      <POINTTABLE pointtableid="3017" name="AQUA Point Scoring" version="2024" />
      <QUALIFY from="2023-08-18" until="2024-08-16" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-08-17" daytime="09:10" endtime="11:50" number="1" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1060" daytime="09:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1367" />
                    <RANKING order="2" place="2" resultid="1168" />
                    <RANKING order="3" place="3" resultid="1754" />
                    <RANKING order="4" place="4" resultid="1377" />
                    <RANKING order="5" place="5" resultid="1864" />
                    <RANKING order="6" place="6" resultid="1406" />
                    <RANKING order="7" place="7" resultid="1530" />
                    <RANKING order="8" place="8" resultid="1593" />
                    <RANKING order="9" place="9" resultid="1396" />
                    <RANKING order="10" place="10" resultid="1201" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1322" />
                    <RANKING order="2" place="2" resultid="1287" />
                    <RANKING order="3" place="3" resultid="1347" />
                    <RANKING order="4" place="4" resultid="1292" />
                    <RANKING order="5" place="5" resultid="1743" />
                    <RANKING order="6" place="6" resultid="1873" />
                    <RANKING order="7" place="7" resultid="1327" />
                    <RANKING order="8" place="8" resultid="1972" />
                    <RANKING order="9" place="9" resultid="1490" />
                    <RANKING order="10" place="10" resultid="1372" />
                    <RANKING order="11" place="11" resultid="1431" />
                    <RANKING order="12" place="12" resultid="1859" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2129" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2130" daytime="09:15" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2131" daytime="09:15" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1063" daytime="09:20" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1064" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2019" />
                    <RANKING order="2" place="2" resultid="1436" />
                    <RANKING order="3" place="3" resultid="1242" />
                    <RANKING order="4" place="4" resultid="1387" />
                    <RANKING order="5" place="5" resultid="1426" />
                    <RANKING order="6" place="6" resultid="1465" />
                    <RANKING order="7" place="7" resultid="2029" />
                    <RANKING order="8" place="8" resultid="1451" />
                    <RANKING order="9" place="9" resultid="2080" />
                    <RANKING order="10" place="10" resultid="1869" />
                    <RANKING order="11" place="11" resultid="1827" />
                    <RANKING order="12" place="-1" resultid="1818" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1312" />
                    <RANKING order="2" place="2" resultid="1967" />
                    <RANKING order="3" place="3" resultid="1337" />
                    <RANKING order="4" place="4" resultid="1485" />
                    <RANKING order="5" place="5" resultid="1352" />
                    <RANKING order="6" place="6" resultid="1277" />
                    <RANKING order="7" place="7" resultid="1307" />
                    <RANKING order="8" place="8" resultid="1342" />
                    <RANKING order="9" place="9" resultid="1192" />
                    <RANKING order="10" place="10" resultid="1392" />
                    <RANKING order="11" place="11" resultid="2043" />
                    <RANKING order="12" place="12" resultid="1461" />
                    <RANKING order="13" place="13" resultid="2088" />
                    <RANKING order="14" place="14" resultid="2119" />
                    <RANKING order="15" place="-1" resultid="1441" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2132" daytime="09:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2133" daytime="09:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2134" daytime="09:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2135" daytime="09:30" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1066" daytime="09:30" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1067" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1673" />
                    <RANKING order="2" place="2" resultid="1940" />
                    <RANKING order="3" place="3" resultid="1663" />
                    <RANKING order="4" place="4" resultid="1171" />
                    <RANKING order="5" place="5" resultid="1693" />
                    <RANKING order="6" place="6" resultid="1628" />
                    <RANKING order="7" place="7" resultid="1221" />
                    <RANKING order="8" place="8" resultid="1764" />
                    <RANKING order="9" place="9" resultid="1623" />
                    <RANKING order="10" place="10" resultid="1782" />
                    <RANKING order="11" place="11" resultid="1738" />
                    <RANKING order="12" place="-1" resultid="1638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1977" />
                    <RANKING order="2" place="2" resultid="1505" />
                    <RANKING order="3" place="3" resultid="1608" />
                    <RANKING order="4" place="4" resultid="2097" />
                    <RANKING order="5" place="5" resultid="2106" />
                    <RANKING order="6" place="6" resultid="1613" />
                    <RANKING order="7" place="7" resultid="1698" />
                    <RANKING order="8" place="8" resultid="1160" />
                    <RANKING order="9" place="9" resultid="2092" />
                    <RANKING order="10" place="10" resultid="1258" />
                    <RANKING order="11" place="11" resultid="1180" />
                    <RANKING order="12" place="12" resultid="1777" />
                    <RANKING order="13" place="13" resultid="1945" />
                    <RANKING order="14" place="-1" resultid="1583" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2136" daytime="09:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2137" daytime="09:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2138" daytime="09:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2139" daytime="09:40" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1069" daytime="09:40" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1070" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1618" />
                    <RANKING order="2" place="2" resultid="1733" />
                    <RANKING order="3" place="3" resultid="2038" />
                    <RANKING order="4" place="4" resultid="1713" />
                    <RANKING order="5" place="5" resultid="1668" />
                    <RANKING order="6" place="6" resultid="1896" />
                    <RANKING order="7" place="7" resultid="1748" />
                    <RANKING order="8" place="8" resultid="1769" />
                    <RANKING order="9" place="-1" resultid="1773" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1525" />
                    <RANKING order="2" place="2" resultid="1997" />
                    <RANKING order="3" place="3" resultid="1175" />
                    <RANKING order="4" place="4" resultid="1553" />
                    <RANKING order="5" place="5" resultid="1573" />
                    <RANKING order="6" place="6" resultid="1935" />
                    <RANKING order="7" place="7" resultid="1558" />
                    <RANKING order="8" place="8" resultid="1212" />
                    <RANKING order="9" place="9" resultid="2071" />
                    <RANKING order="10" place="10" resultid="1578" />
                    <RANKING order="11" place="11" resultid="1792" />
                    <RANKING order="12" place="12" resultid="2066" />
                    <RANKING order="13" place="13" resultid="2058" />
                    <RANKING order="14" place="14" resultid="1183" />
                    <RANKING order="15" place="15" resultid="1563" />
                    <RANKING order="16" place="-1" resultid="1535" />
                    <RANKING order="17" place="-1" resultid="1540" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2140" daytime="09:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2141" daytime="09:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2142" daytime="09:45" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2143" daytime="09:50" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1072" daytime="09:50" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1073" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1481" />
                    <RANKING order="2" place="2" resultid="1363" />
                    <RANKING order="3" place="3" resultid="1422" />
                    <RANKING order="4" place="4" resultid="1883" />
                    <RANKING order="5" place="5" resultid="1407" />
                    <RANKING order="6" place="6" resultid="1983" />
                    <RANKING order="7" place="7" resultid="1236" />
                    <RANKING order="8" place="8" resultid="1927" />
                    <RANKING order="9" place="9" resultid="1205" />
                    <RANKING order="10" place="10" resultid="1501" />
                    <RANKING order="11" place="11" resultid="2007" />
                    <RANKING order="12" place="12" resultid="2025" />
                    <RANKING order="13" place="13" resultid="1169" />
                    <RANKING order="14" place="14" resultid="1879" />
                    <RANKING order="15" place="15" resultid="1549" />
                    <RANKING order="16" place="16" resultid="1202" />
                    <RANKING order="17" place="17" resultid="1397" />
                    <RANKING order="18" place="18" resultid="1224" />
                    <RANKING order="19" place="19" resultid="2103" />
                    <RANKING order="20" place="-1" resultid="1412" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1074" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1447" />
                    <RANKING order="2" place="2" resultid="1589" />
                    <RANKING order="3" place="3" resultid="1383" />
                    <RANKING order="4" place="4" resultid="2076" />
                    <RANKING order="5" place="5" resultid="1973" />
                    <RANKING order="6" place="6" resultid="1373" />
                    <RANKING order="7" place="7" resultid="1988" />
                    <RANKING order="8" place="8" resultid="1333" />
                    <RANKING order="9" place="9" resultid="1348" />
                    <RANKING order="10" place="10" resultid="1197" />
                    <RANKING order="11" place="11" resultid="1218" />
                    <RANKING order="12" place="12" resultid="1147" />
                    <RANKING order="13" place="13" resultid="1860" />
                    <RANKING order="14" place="14" resultid="1491" />
                    <RANKING order="15" place="15" resultid="1252" />
                    <RANKING order="16" place="-1" resultid="2085" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2144" daytime="09:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2145" daytime="09:55" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2146" daytime="09:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2147" daytime="10:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2148" daytime="10:00" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1075" daytime="10:05" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1076" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1150" />
                    <RANKING order="2" place="2" resultid="1603" />
                    <RANKING order="3" place="3" resultid="2033" />
                    <RANKING order="4" place="4" resultid="1456" />
                    <RANKING order="5" place="5" resultid="1357" />
                    <RANKING order="6" place="6" resultid="1470" />
                    <RANKING order="7" place="7" resultid="1416" />
                    <RANKING order="8" place="8" resultid="2010" />
                    <RANKING order="9" place="9" resultid="1401" />
                    <RANKING order="10" place="10" resultid="1887" />
                    <RANKING order="11" place="11" resultid="1475" />
                    <RANKING order="12" place="12" resultid="1265" />
                    <RANKING order="13" place="13" resultid="2030" />
                    <RANKING order="14" place="14" resultid="1930" />
                    <RANKING order="15" place="15" resultid="1917" />
                    <RANKING order="16" place="16" resultid="1870" />
                    <RANKING order="17" place="17" resultid="1828" />
                    <RANKING order="18" place="-1" resultid="1831" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1077" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1272" />
                    <RANKING order="2" place="2" resultid="1921" />
                    <RANKING order="3" place="3" resultid="1317" />
                    <RANKING order="4" place="4" resultid="1208" />
                    <RANKING order="5" place="5" resultid="1302" />
                    <RANKING order="6" place="6" resultid="1297" />
                    <RANKING order="7" place="7" resultid="1282" />
                    <RANKING order="8" place="8" resultid="1353" />
                    <RANKING order="9" place="9" resultid="2063" />
                    <RANKING order="10" place="10" resultid="1188" />
                    <RANKING order="11" place="11" resultid="1308" />
                    <RANKING order="12" place="12" resultid="1462" />
                    <RANKING order="13" place="13" resultid="1193" />
                    <RANKING order="14" place="14" resultid="2089" />
                    <RANKING order="15" place="15" resultid="1393" />
                    <RANKING order="16" place="16" resultid="2002" />
                    <RANKING order="17" place="17" resultid="1442" />
                    <RANKING order="18" place="18" resultid="1227" />
                    <RANKING order="19" place="19" resultid="2120" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2149" daytime="10:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2150" daytime="10:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2151" daytime="10:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2152" daytime="10:10" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2153" daytime="10:15" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1078" daytime="10:15" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1079" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1950" />
                    <RANKING order="2" place="2" resultid="1688" />
                    <RANKING order="3" place="3" resultid="1648" />
                    <RANKING order="4" place="4" resultid="1718" />
                    <RANKING order="5" place="5" resultid="1629" />
                    <RANKING order="6" place="6" resultid="1683" />
                    <RANKING order="7" place="7" resultid="1823" />
                    <RANKING order="8" place="8" resultid="1624" />
                    <RANKING order="9" place="9" resultid="1664" />
                    <RANKING order="10" place="10" resultid="1783" />
                    <RANKING order="11" place="-1" resultid="1639" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1080" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2048" />
                    <RANKING order="2" place="2" resultid="1653" />
                    <RANKING order="3" place="3" resultid="2053" />
                    <RANKING order="4" place="4" resultid="1155" />
                    <RANKING order="5" place="5" resultid="1598" />
                    <RANKING order="6" place="6" resultid="2098" />
                    <RANKING order="7" place="7" resultid="1510" />
                    <RANKING order="8" place="8" resultid="1609" />
                    <RANKING order="9" place="9" resultid="1568" />
                    <RANKING order="10" place="10" resultid="1900" />
                    <RANKING order="11" place="11" resultid="1614" />
                    <RANKING order="12" place="12" resultid="1161" />
                    <RANKING order="13" place="13" resultid="2093" />
                    <RANKING order="14" place="14" resultid="1778" />
                    <RANKING order="15" place="-1" resultid="1544" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2154" daytime="10:15" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2155" daytime="10:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2156" daytime="10:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2157" daytime="10:25" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1081" daytime="10:25" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1082" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1633" />
                    <RANKING order="2" place="2" resultid="1787" />
                    <RANKING order="3" place="3" resultid="1678" />
                    <RANKING order="4" place="4" resultid="1669" />
                    <RANKING order="5" place="5" resultid="1909" />
                    <RANKING order="6" place="6" resultid="1892" />
                    <RANKING order="7" place="7" resultid="1714" />
                    <RANKING order="8" place="8" resultid="1897" />
                    <RANKING order="9" place="9" resultid="1749" />
                    <RANKING order="10" place="10" resultid="1728" />
                    <RANKING order="11" place="11" resultid="1723" />
                    <RANKING order="12" place="12" resultid="1708" />
                    <RANKING order="13" place="13" resultid="1759" />
                    <RANKING order="14" place="14" resultid="1770" />
                    <RANKING order="15" place="-1" resultid="1774" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1904" />
                    <RANKING order="2" place="2" resultid="1703" />
                    <RANKING order="3" place="3" resultid="1520" />
                    <RANKING order="4" place="4" resultid="1495" />
                    <RANKING order="5" place="5" resultid="1658" />
                    <RANKING order="6" place="6" resultid="1526" />
                    <RANKING order="7" place="7" resultid="1992" />
                    <RANKING order="8" place="8" resultid="1515" />
                    <RANKING order="9" place="9" resultid="1559" />
                    <RANKING order="10" place="10" resultid="2072" />
                    <RANKING order="11" place="11" resultid="1230" />
                    <RANKING order="12" place="12" resultid="2014" />
                    <RANKING order="13" place="13" resultid="1793" />
                    <RANKING order="14" place="14" resultid="1184" />
                    <RANKING order="15" place="-1" resultid="1536" />
                    <RANKING order="16" place="-1" resultid="1643" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2158" daytime="10:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2159" daytime="10:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2160" daytime="10:35" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2161" daytime="10:35" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1084" daytime="10:40" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1085" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1865" />
                    <RANKING order="2" place="2" resultid="1755" />
                    <RANKING order="3" place="3" resultid="1368" />
                    <RANKING order="4" place="4" resultid="1362" />
                    <RANKING order="5" place="5" resultid="1982" />
                    <RANKING order="6" place="6" resultid="1378" />
                    <RANKING order="7" place="7" resultid="2024" />
                    <RANKING order="8" place="8" resultid="1480" />
                    <RANKING order="9" place="9" resultid="1421" />
                    <RANKING order="10" place="10" resultid="2006" />
                    <RANKING order="11" place="11" resultid="1882" />
                    <RANKING order="12" place="12" resultid="1235" />
                    <RANKING order="13" place="13" resultid="1500" />
                    <RANKING order="14" place="14" resultid="1548" />
                    <RANKING order="15" place="15" resultid="1531" />
                    <RANKING order="16" place="16" resultid="1594" />
                    <RANKING order="17" place="17" resultid="1926" />
                    <RANKING order="18" place="18" resultid="1878" />
                    <RANKING order="19" place="19" resultid="2102" />
                    <RANKING order="20" place="-1" resultid="1204" />
                    <RANKING order="21" place="-1" resultid="1411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1288" />
                    <RANKING order="2" place="2" resultid="1446" />
                    <RANKING order="3" place="3" resultid="1293" />
                    <RANKING order="4" place="4" resultid="1382" />
                    <RANKING order="5" place="5" resultid="1328" />
                    <RANKING order="6" place="6" resultid="1588" />
                    <RANKING order="7" place="7" resultid="1332" />
                    <RANKING order="8" place="8" resultid="1744" />
                    <RANKING order="9" place="9" resultid="1245" />
                    <RANKING order="10" place="10" resultid="1987" />
                    <RANKING order="11" place="11" resultid="1146" />
                    <RANKING order="12" place="12" resultid="1874" />
                    <RANKING order="13" place="13" resultid="1196" />
                    <RANKING order="14" place="14" resultid="1323" />
                    <RANKING order="15" place="15" resultid="1959" />
                    <RANKING order="16" place="16" resultid="1432" />
                    <RANKING order="17" place="17" resultid="1217" />
                    <RANKING order="18" place="-1" resultid="2075" />
                    <RANKING order="19" place="-1" resultid="2084" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2162" daytime="10:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2163" daytime="10:45" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2164" daytime="10:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2165" daytime="10:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2166" daytime="10:55" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1087" daytime="11:00" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1088" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1358" />
                    <RANKING order="2" place="2" resultid="1427" />
                    <RANKING order="3" place="3" resultid="2034" />
                    <RANKING order="4" place="4" resultid="1151" />
                    <RANKING order="5" place="5" resultid="1604" />
                    <RANKING order="6" place="6" resultid="1452" />
                    <RANKING order="7" place="7" resultid="1471" />
                    <RANKING order="8" place="8" resultid="1888" />
                    <RANKING order="9" place="9" resultid="1457" />
                    <RANKING order="10" place="10" resultid="2020" />
                    <RANKING order="11" place="11" resultid="1819" />
                    <RANKING order="12" place="12" resultid="1437" />
                    <RANKING order="13" place="13" resultid="1417" />
                    <RANKING order="14" place="14" resultid="1466" />
                    <RANKING order="15" place="15" resultid="1476" />
                    <RANKING order="16" place="16" resultid="2011" />
                    <RANKING order="17" place="17" resultid="1388" />
                    <RANKING order="18" place="18" resultid="1402" />
                    <RANKING order="19" place="19" resultid="2081" />
                    <RANKING order="20" place="20" resultid="1931" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1273" />
                    <RANKING order="2" place="2" resultid="1313" />
                    <RANKING order="3" place="3" resultid="1303" />
                    <RANKING order="4" place="4" resultid="1968" />
                    <RANKING order="5" place="5" resultid="1318" />
                    <RANKING order="6" place="6" resultid="1283" />
                    <RANKING order="7" place="7" resultid="1338" />
                    <RANKING order="8" place="8" resultid="1249" />
                    <RANKING order="9" place="9" resultid="1922" />
                    <RANKING order="10" place="10" resultid="1298" />
                    <RANKING order="11" place="11" resultid="1278" />
                    <RANKING order="12" place="12" resultid="1343" />
                    <RANKING order="13" place="13" resultid="1486" />
                    <RANKING order="14" place="14" resultid="1209" />
                    <RANKING order="15" place="15" resultid="1189" />
                    <RANKING order="16" place="16" resultid="2044" />
                    <RANKING order="17" place="17" resultid="2003" />
                    <RANKING order="18" place="18" resultid="2064" />
                    <RANKING order="19" place="19" resultid="2111" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2167" daytime="11:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2168" daytime="11:05" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2169" daytime="11:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2170" daytime="11:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2171" daytime="11:20" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1090" daytime="11:25" gender="F" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1091" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1941" />
                    <RANKING order="2" place="2" resultid="1694" />
                    <RANKING order="3" place="3" resultid="1649" />
                    <RANKING order="4" place="4" resultid="1951" />
                    <RANKING order="5" place="5" resultid="1674" />
                    <RANKING order="6" place="6" resultid="1689" />
                    <RANKING order="7" place="7" resultid="1172" />
                    <RANKING order="8" place="8" resultid="1222" />
                    <RANKING order="9" place="9" resultid="1739" />
                    <RANKING order="10" place="10" resultid="1684" />
                    <RANKING order="11" place="11" resultid="1765" />
                    <RANKING order="12" place="12" resultid="1824" />
                    <RANKING order="13" place="13" resultid="1719" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1092" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1978" />
                    <RANKING order="2" place="2" resultid="1506" />
                    <RANKING order="3" place="3" resultid="2049" />
                    <RANKING order="4" place="4" resultid="2107" />
                    <RANKING order="5" place="5" resultid="1699" />
                    <RANKING order="6" place="6" resultid="1599" />
                    <RANKING order="7" place="7" resultid="1156" />
                    <RANKING order="8" place="8" resultid="1946" />
                    <RANKING order="9" place="9" resultid="2054" />
                    <RANKING order="10" place="10" resultid="1181" />
                    <RANKING order="11" place="11" resultid="1511" />
                    <RANKING order="12" place="12" resultid="1654" />
                    <RANKING order="13" place="13" resultid="1259" />
                    <RANKING order="14" place="14" resultid="1955" />
                    <RANKING order="15" place="15" resultid="1901" />
                    <RANKING order="16" place="16" resultid="1569" />
                    <RANKING order="17" place="-1" resultid="1545" />
                    <RANKING order="18" place="-1" resultid="1584" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2172" daytime="11:25" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2173" daytime="11:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2174" daytime="11:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2175" daytime="11:30" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1093" daytime="11:35" gender="M" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1094" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1634" />
                    <RANKING order="2" place="2" resultid="2039" />
                    <RANKING order="3" place="3" resultid="1910" />
                    <RANKING order="4" place="4" resultid="1679" />
                    <RANKING order="5" place="5" resultid="1619" />
                    <RANKING order="6" place="6" resultid="1788" />
                    <RANKING order="7" place="7" resultid="1709" />
                    <RANKING order="8" place="8" resultid="1893" />
                    <RANKING order="9" place="9" resultid="1729" />
                    <RANKING order="10" place="10" resultid="1734" />
                    <RANKING order="11" place="11" resultid="1724" />
                    <RANKING order="12" place="12" resultid="1760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1579" />
                    <RANKING order="2" place="2" resultid="1905" />
                    <RANKING order="3" place="3" resultid="1659" />
                    <RANKING order="4" place="4" resultid="1496" />
                    <RANKING order="5" place="5" resultid="1521" />
                    <RANKING order="6" place="6" resultid="1176" />
                    <RANKING order="7" place="7" resultid="1516" />
                    <RANKING order="8" place="8" resultid="1998" />
                    <RANKING order="9" place="9" resultid="1704" />
                    <RANKING order="10" place="10" resultid="1993" />
                    <RANKING order="11" place="11" resultid="1574" />
                    <RANKING order="12" place="12" resultid="2067" />
                    <RANKING order="13" place="13" resultid="1936" />
                    <RANKING order="14" place="14" resultid="2015" />
                    <RANKING order="15" place="15" resultid="2059" />
                    <RANKING order="16" place="16" resultid="1231" />
                    <RANKING order="17" place="17" resultid="1213" />
                    <RANKING order="18" place="18" resultid="1554" />
                    <RANKING order="19" place="19" resultid="1564" />
                    <RANKING order="20" place="-1" resultid="1541" />
                    <RANKING order="21" place="-1" resultid="1644" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2176" daytime="11:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2177" daytime="11:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2178" daytime="11:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2179" daytime="11:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2180" daytime="11:50" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-08-17" daytime="15:40" endtime="22:26" number="2" officialmeeting="15:00" teamleadermeeting="15:30" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1096" daytime="15:40" gender="F" number="13" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1097" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1806" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2181" daytime="15:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1098" daytime="15:40" gender="M" number="14" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2122" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1100" daytime="15:40" gender="F" number="15" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1101" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1866" />
                    <RANKING order="2" place="2" resultid="1364" />
                    <RANKING order="3" place="3" resultid="1369" />
                    <RANKING order="4" place="4" resultid="1756" />
                    <RANKING order="5" place="5" resultid="1408" />
                    <RANKING order="6" place="6" resultid="1379" />
                    <RANKING order="7" place="7" resultid="1482" />
                    <RANKING order="8" place="8" resultid="1884" />
                    <RANKING order="9" place="9" resultid="1423" />
                    <RANKING order="10" place="10" resultid="1502" />
                    <RANKING order="11" place="11" resultid="1595" />
                    <RANKING order="12" place="12" resultid="1398" />
                    <RANKING order="13" place="-1" resultid="1413" />
                    <RANKING order="14" place="-1" resultid="1984" />
                    <RANKING order="15" place="-1" resultid="1532" />
                    <RANKING order="16" place="-1" resultid="1963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1294" />
                    <RANKING order="2" place="2" resultid="1289" />
                    <RANKING order="3" place="3" resultid="1384" />
                    <RANKING order="4" place="4" resultid="1329" />
                    <RANKING order="5" place="5" resultid="1349" />
                    <RANKING order="6" place="6" resultid="1590" />
                    <RANKING order="7" place="7" resultid="1324" />
                    <RANKING order="8" place="8" resultid="1989" />
                    <RANKING order="9" place="9" resultid="1374" />
                    <RANKING order="10" place="10" resultid="1974" />
                    <RANKING order="11" place="11" resultid="2077" />
                    <RANKING order="12" place="12" resultid="1960" />
                    <RANKING order="13" place="13" resultid="1492" />
                    <RANKING order="14" place="14" resultid="1433" />
                    <RANKING order="15" place="-1" resultid="1745" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2182" daytime="15:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2183" daytime="15:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2184" daytime="15:55" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2185" daytime="16:00" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1103" daytime="16:05" gender="M" number="16" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1104" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1428" />
                    <RANKING order="2" place="2" resultid="1359" />
                    <RANKING order="3" place="3" resultid="2035" />
                    <RANKING order="4" place="4" resultid="1820" />
                    <RANKING order="5" place="5" resultid="2021" />
                    <RANKING order="6" place="6" resultid="1605" />
                    <RANKING order="7" place="7" resultid="1438" />
                    <RANKING order="8" place="8" resultid="1453" />
                    <RANKING order="9" place="9" resultid="1458" />
                    <RANKING order="10" place="10" resultid="1467" />
                    <RANKING order="11" place="11" resultid="1477" />
                    <RANKING order="12" place="12" resultid="1418" />
                    <RANKING order="13" place="13" resultid="1889" />
                    <RANKING order="14" place="14" resultid="1403" />
                    <RANKING order="15" place="15" resultid="1266" />
                    <RANKING order="16" place="16" resultid="1932" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1274" />
                    <RANKING order="2" place="2" resultid="1314" />
                    <RANKING order="3" place="3" resultid="1969" />
                    <RANKING order="4" place="4" resultid="1304" />
                    <RANKING order="5" place="5" resultid="1339" />
                    <RANKING order="6" place="6" resultid="1923" />
                    <RANKING order="7" place="7" resultid="1309" />
                    <RANKING order="8" place="8" resultid="1299" />
                    <RANKING order="9" place="9" resultid="1354" />
                    <RANKING order="10" place="10" resultid="2045" />
                    <RANKING order="11" place="11" resultid="1443" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2186" daytime="16:05" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2187" daytime="16:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2188" daytime="16:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2189" daytime="16:15" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1106" daytime="16:20" gender="F" number="17" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1107" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1942" />
                    <RANKING order="2" place="2" resultid="1675" />
                    <RANKING order="3" place="3" resultid="1952" />
                    <RANKING order="4" place="4" resultid="1690" />
                    <RANKING order="5" place="5" resultid="1650" />
                    <RANKING order="6" place="6" resultid="1685" />
                    <RANKING order="7" place="7" resultid="1630" />
                    <RANKING order="8" place="8" resultid="1695" />
                    <RANKING order="9" place="9" resultid="1665" />
                    <RANKING order="10" place="10" resultid="1625" />
                    <RANKING order="11" place="11" resultid="1740" />
                    <RANKING order="12" place="12" resultid="1784" />
                    <RANKING order="13" place="-1" resultid="1766" />
                    <RANKING order="14" place="-1" resultid="1640" />
                    <RANKING order="15" place="-1" resultid="1720" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1108" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1979" />
                    <RANKING order="2" place="2" resultid="1507" />
                    <RANKING order="3" place="3" resultid="1700" />
                    <RANKING order="4" place="4" resultid="2050" />
                    <RANKING order="5" place="5" resultid="1512" />
                    <RANKING order="6" place="6" resultid="2099" />
                    <RANKING order="7" place="7" resultid="1655" />
                    <RANKING order="8" place="8" resultid="1956" />
                    <RANKING order="9" place="9" resultid="2108" />
                    <RANKING order="10" place="10" resultid="1600" />
                    <RANKING order="11" place="11" resultid="1157" />
                    <RANKING order="12" place="12" resultid="1610" />
                    <RANKING order="13" place="13" resultid="1947" />
                    <RANKING order="14" place="14" resultid="2055" />
                    <RANKING order="15" place="15" resultid="1162" />
                    <RANKING order="16" place="16" resultid="2094" />
                    <RANKING order="17" place="17" resultid="1615" />
                    <RANKING order="18" place="18" resultid="1570" />
                    <RANKING order="19" place="19" resultid="1779" />
                    <RANKING order="20" place="-1" resultid="1585" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2190" daytime="16:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2191" daytime="16:25" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2192" daytime="16:25" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2193" daytime="16:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2194" daytime="16:30" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1109" daytime="16:35" gender="M" number="18" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1110" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1636" />
                    <RANKING order="2" place="2" resultid="2041" />
                    <RANKING order="3" place="3" resultid="1681" />
                    <RANKING order="4" place="4" resultid="1621" />
                    <RANKING order="5" place="5" resultid="1671" />
                    <RANKING order="6" place="6" resultid="1736" />
                    <RANKING order="7" place="7" resultid="1790" />
                    <RANKING order="8" place="8" resultid="1711" />
                    <RANKING order="9" place="9" resultid="1716" />
                    <RANKING order="10" place="10" resultid="1912" />
                    <RANKING order="11" place="11" resultid="1751" />
                    <RANKING order="12" place="12" resultid="1731" />
                    <RANKING order="13" place="13" resultid="1762" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1498" />
                    <RANKING order="2" place="2" resultid="1528" />
                    <RANKING order="3" place="3" resultid="1518" />
                    <RANKING order="4" place="4" resultid="1581" />
                    <RANKING order="5" place="5" resultid="1576" />
                    <RANKING order="6" place="6" resultid="1523" />
                    <RANKING order="7" place="7" resultid="1178" />
                    <RANKING order="8" place="8" resultid="1166" />
                    <RANKING order="9" place="9" resultid="1706" />
                    <RANKING order="10" place="10" resultid="1995" />
                    <RANKING order="11" place="11" resultid="1661" />
                    <RANKING order="12" place="12" resultid="1907" />
                    <RANKING order="13" place="13" resultid="2000" />
                    <RANKING order="14" place="13" resultid="2017" />
                    <RANKING order="15" place="15" resultid="1561" />
                    <RANKING order="16" place="16" resultid="1556" />
                    <RANKING order="17" place="17" resultid="2061" />
                    <RANKING order="18" place="18" resultid="1215" />
                    <RANKING order="19" place="19" resultid="2069" />
                    <RANKING order="20" place="20" resultid="1795" />
                    <RANKING order="21" place="21" resultid="1566" />
                    <RANKING order="22" place="-1" resultid="1538" />
                    <RANKING order="23" place="-1" resultid="1646" />
                    <RANKING order="24" place="-1" resultid="1938" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2195" daytime="16:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2196" daytime="16:35" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2197" daytime="16:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2198" daytime="16:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2199" daytime="16:45" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1112" daytime="16:45" gender="F" number="19" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2123" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1840" />
                    <RANKING order="2" place="2" resultid="1834" />
                    <RANKING order="3" place="3" resultid="1809" />
                    <RANKING order="4" place="-1" resultid="1800" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2200" daytime="16:45" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1114" daytime="16:50" gender="M" number="20" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2124" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1846" />
                    <RANKING order="2" place="2" resultid="1849" />
                    <RANKING order="3" place="3" resultid="2114" />
                    <RANKING order="4" place="-1" resultid="1797" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2201" daytime="16:50" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1116" daytime="16:50" gender="F" number="21" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1117" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1867" />
                    <RANKING order="2" place="2" resultid="1409" />
                    <RANKING order="3" place="3" resultid="1550" />
                    <RANKING order="4" place="4" resultid="2026" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1448" />
                    <RANKING order="2" place="2" resultid="1334" />
                    <RANKING order="3" place="3" resultid="1350" />
                    <RANKING order="4" place="4" resultid="1875" />
                    <RANKING order="5" place="5" resultid="1246" />
                    <RANKING order="6" place="6" resultid="1198" />
                    <RANKING order="7" place="7" resultid="1914" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2202" daytime="16:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2203" daytime="16:55" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1119" daytime="16:55" gender="M" number="22" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1120" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1152" />
                    <RANKING order="2" place="2" resultid="1389" />
                    <RANKING order="3" place="3" resultid="1360" />
                    <RANKING order="4" place="4" resultid="1454" />
                    <RANKING order="5" place="5" resultid="1472" />
                    <RANKING order="6" place="6" resultid="1459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1275" />
                    <RANKING order="2" place="2" resultid="1239" />
                    <RANKING order="3" place="3" resultid="1284" />
                    <RANKING order="4" place="4" resultid="1487" />
                    <RANKING order="5" place="5" resultid="1344" />
                    <RANKING order="6" place="6" resultid="1279" />
                    <RANKING order="7" place="7" resultid="1319" />
                    <RANKING order="8" place="8" resultid="2046" />
                    <RANKING order="9" place="-1" resultid="1924" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2204" daytime="16:55" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2205" daytime="17:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1122" daytime="17:00" gender="F" number="23" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2125" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1255" />
                    <RANKING order="2" place="2" resultid="1812" />
                    <RANKING order="3" place="3" resultid="1852" />
                    <RANKING order="4" place="4" resultid="1835" />
                    <RANKING order="5" place="5" resultid="1855" />
                    <RANKING order="6" place="-1" resultid="1815" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2206" daytime="17:00" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1124" daytime="17:05" gender="M" number="24" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2126" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1262" />
                    <RANKING order="2" place="2" resultid="1803" />
                    <RANKING order="3" place="-1" resultid="1837" />
                    <RANKING order="4" place="-1" resultid="1843" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2207" daytime="17:05" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1126" daytime="17:10" gender="F" number="25" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1127" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1943" />
                    <RANKING order="2" place="2" resultid="1696" />
                    <RANKING order="3" place="3" resultid="1651" />
                    <RANKING order="4" place="4" resultid="1173" />
                    <RANKING order="5" place="5" resultid="1676" />
                    <RANKING order="6" place="6" resultid="1953" />
                    <RANKING order="7" place="7" resultid="1691" />
                    <RANKING order="8" place="8" resultid="1825" />
                    <RANKING order="9" place="9" resultid="1767" />
                    <RANKING order="10" place="10" resultid="1741" />
                    <RANKING order="11" place="11" resultid="1631" />
                    <RANKING order="12" place="12" resultid="1666" />
                    <RANKING order="13" place="13" resultid="1686" />
                    <RANKING order="14" place="14" resultid="1626" />
                    <RANKING order="15" place="15" resultid="1785" />
                    <RANKING order="16" place="-1" resultid="1641" />
                    <RANKING order="17" place="-1" resultid="1721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1980" />
                    <RANKING order="2" place="2" resultid="1508" />
                    <RANKING order="3" place="3" resultid="2051" />
                    <RANKING order="4" place="4" resultid="1158" />
                    <RANKING order="5" place="5" resultid="1701" />
                    <RANKING order="6" place="6" resultid="2056" />
                    <RANKING order="7" place="7" resultid="2109" />
                    <RANKING order="8" place="8" resultid="2100" />
                    <RANKING order="9" place="9" resultid="1948" />
                    <RANKING order="10" place="10" resultid="1601" />
                    <RANKING order="11" place="11" resultid="1656" />
                    <RANKING order="12" place="12" resultid="1163" />
                    <RANKING order="13" place="13" resultid="1260" />
                    <RANKING order="14" place="14" resultid="1611" />
                    <RANKING order="15" place="14" resultid="1616" />
                    <RANKING order="16" place="16" resultid="1513" />
                    <RANKING order="17" place="17" resultid="1957" />
                    <RANKING order="18" place="18" resultid="1902" />
                    <RANKING order="19" place="19" resultid="1571" />
                    <RANKING order="20" place="20" resultid="2095" />
                    <RANKING order="21" place="21" resultid="1780" />
                    <RANKING order="22" place="-1" resultid="1546" />
                    <RANKING order="23" place="-1" resultid="1586" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2208" daytime="17:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2209" daytime="17:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2210" daytime="17:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2211" daytime="17:15" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2212" daytime="17:15" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1129" daytime="17:20" gender="M" number="26" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1130" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1635" />
                    <RANKING order="2" place="2" resultid="2040" />
                    <RANKING order="3" place="3" resultid="1620" />
                    <RANKING order="4" place="4" resultid="1680" />
                    <RANKING order="5" place="5" resultid="1911" />
                    <RANKING order="6" place="6" resultid="1894" />
                    <RANKING order="7" place="7" resultid="1789" />
                    <RANKING order="8" place="8" resultid="1670" />
                    <RANKING order="9" place="9" resultid="2117" />
                    <RANKING order="10" place="10" resultid="1715" />
                    <RANKING order="11" place="11" resultid="1710" />
                    <RANKING order="12" place="12" resultid="1898" />
                    <RANKING order="13" place="13" resultid="1730" />
                    <RANKING order="14" place="14" resultid="1725" />
                    <RANKING order="15" place="15" resultid="1771" />
                    <RANKING order="16" place="16" resultid="1761" />
                    <RANKING order="17" place="17" resultid="1750" />
                    <RANKING order="18" place="-1" resultid="1735" />
                    <RANKING order="19" place="-1" resultid="1775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1580" />
                    <RANKING order="2" place="2" resultid="1906" />
                    <RANKING order="3" place="3" resultid="1497" />
                    <RANKING order="4" place="4" resultid="1527" />
                    <RANKING order="5" place="5" resultid="1660" />
                    <RANKING order="6" place="6" resultid="1999" />
                    <RANKING order="7" place="7" resultid="1177" />
                    <RANKING order="8" place="8" resultid="1517" />
                    <RANKING order="9" place="9" resultid="1522" />
                    <RANKING order="10" place="10" resultid="1165" />
                    <RANKING order="11" place="11" resultid="1705" />
                    <RANKING order="12" place="11" resultid="1937" />
                    <RANKING order="13" place="13" resultid="1214" />
                    <RANKING order="14" place="14" resultid="1575" />
                    <RANKING order="15" place="15" resultid="2068" />
                    <RANKING order="16" place="16" resultid="2016" />
                    <RANKING order="17" place="17" resultid="2073" />
                    <RANKING order="18" place="18" resultid="1994" />
                    <RANKING order="19" place="19" resultid="1555" />
                    <RANKING order="20" place="20" resultid="2060" />
                    <RANKING order="21" place="21" resultid="1560" />
                    <RANKING order="22" place="22" resultid="1232" />
                    <RANKING order="23" place="23" resultid="1794" />
                    <RANKING order="24" place="24" resultid="1185" />
                    <RANKING order="25" place="25" resultid="1565" />
                    <RANKING order="26" place="-1" resultid="1537" />
                    <RANKING order="27" place="-1" resultid="1542" />
                    <RANKING order="28" place="-1" resultid="1645" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2213" daytime="17:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2214" daytime="17:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2215" daytime="17:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2216" daytime="17:25" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2217" daytime="17:25" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2218" daytime="17:25" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1132" daytime="17:30" gender="F" number="27" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2127" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1807" />
                    <RANKING order="2" place="2" resultid="1813" />
                    <RANKING order="3" place="3" resultid="1841" />
                    <RANKING order="4" place="4" resultid="1853" />
                    <RANKING order="5" place="5" resultid="1856" />
                    <RANKING order="6" place="6" resultid="1810" />
                    <RANKING order="7" place="-1" resultid="1256" />
                    <RANKING order="8" place="-1" resultid="1801" />
                    <RANKING order="9" place="-1" resultid="1816" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2219" daytime="17:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2220" daytime="17:30" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1134" daytime="17:35" gender="M" number="28" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="2128" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1263" />
                    <RANKING order="2" place="2" resultid="2115" />
                    <RANKING order="3" place="3" resultid="1838" />
                    <RANKING order="4" place="4" resultid="1847" />
                    <RANKING order="5" place="5" resultid="1850" />
                    <RANKING order="6" place="-1" resultid="1798" />
                    <RANKING order="7" place="-1" resultid="1804" />
                    <RANKING order="8" place="-1" resultid="1844" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2221" daytime="17:35" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1136" daytime="17:35" gender="F" number="29" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1137" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1414" />
                    <RANKING order="2" place="2" resultid="1380" />
                    <RANKING order="3" place="3" resultid="1757" />
                    <RANKING order="4" place="4" resultid="1365" />
                    <RANKING order="5" place="5" resultid="1885" />
                    <RANKING order="6" place="6" resultid="1237" />
                    <RANKING order="7" place="7" resultid="1483" />
                    <RANKING order="8" place="8" resultid="1370" />
                    <RANKING order="9" place="9" resultid="2008" />
                    <RANKING order="10" place="10" resultid="1206" />
                    <RANKING order="11" place="11" resultid="1424" />
                    <RANKING order="12" place="12" resultid="2027" />
                    <RANKING order="13" place="13" resultid="1985" />
                    <RANKING order="14" place="14" resultid="1503" />
                    <RANKING order="15" place="15" resultid="1551" />
                    <RANKING order="16" place="16" resultid="1928" />
                    <RANKING order="17" place="17" resultid="1596" />
                    <RANKING order="18" place="18" resultid="1399" />
                    <RANKING order="19" place="19" resultid="1880" />
                    <RANKING order="20" place="20" resultid="1964" />
                    <RANKING order="21" place="21" resultid="1225" />
                    <RANKING order="22" place="22" resultid="2104" />
                    <RANKING order="23" place="-1" resultid="1533" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1449" />
                    <RANKING order="2" place="2" resultid="1385" />
                    <RANKING order="3" place="3" resultid="1295" />
                    <RANKING order="4" place="4" resultid="1290" />
                    <RANKING order="5" place="5" resultid="1591" />
                    <RANKING order="6" place="6" resultid="1335" />
                    <RANKING order="7" place="7" resultid="1975" />
                    <RANKING order="8" place="8" resultid="1330" />
                    <RANKING order="9" place="9" resultid="1746" />
                    <RANKING order="10" place="10" resultid="1990" />
                    <RANKING order="11" place="11" resultid="1375" />
                    <RANKING order="12" place="12" resultid="2078" />
                    <RANKING order="13" place="13" resultid="1325" />
                    <RANKING order="14" place="14" resultid="1915" />
                    <RANKING order="15" place="15" resultid="1199" />
                    <RANKING order="16" place="16" resultid="1247" />
                    <RANKING order="17" place="17" resultid="1148" />
                    <RANKING order="18" place="18" resultid="1961" />
                    <RANKING order="19" place="19" resultid="1861" />
                    <RANKING order="20" place="20" resultid="1876" />
                    <RANKING order="21" place="21" resultid="1219" />
                    <RANKING order="22" place="22" resultid="1434" />
                    <RANKING order="23" place="23" resultid="1493" />
                    <RANKING order="24" place="24" resultid="1253" />
                    <RANKING order="25" place="-1" resultid="2086" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2222" daytime="17:35" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2223" daytime="17:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2224" daytime="17:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2225" daytime="17:45" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2226" daytime="17:45" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2227" daytime="17:45" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1139" daytime="17:50" gender="M" number="30" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="26" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1140" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1243" />
                    <RANKING order="2" place="2" resultid="1153" />
                    <RANKING order="3" place="3" resultid="2036" />
                    <RANKING order="4" place="4" resultid="1606" />
                    <RANKING order="5" place="5" resultid="1429" />
                    <RANKING order="6" place="6" resultid="2022" />
                    <RANKING order="7" place="7" resultid="1821" />
                    <RANKING order="8" place="8" resultid="1439" />
                    <RANKING order="9" place="9" resultid="1473" />
                    <RANKING order="10" place="10" resultid="2012" />
                    <RANKING order="11" place="11" resultid="2031" />
                    <RANKING order="12" place="12" resultid="1390" />
                    <RANKING order="13" place="13" resultid="1404" />
                    <RANKING order="14" place="14" resultid="1890" />
                    <RANKING order="15" place="15" resultid="1419" />
                    <RANKING order="16" place="16" resultid="1468" />
                    <RANKING order="17" place="17" resultid="1478" />
                    <RANKING order="18" place="18" resultid="2082" />
                    <RANKING order="19" place="19" resultid="1267" />
                    <RANKING order="20" place="20" resultid="1933" />
                    <RANKING order="21" place="21" resultid="1871" />
                    <RANKING order="22" place="22" resultid="1918" />
                    <RANKING order="23" place="23" resultid="1829" />
                    <RANKING order="24" place="24" resultid="1832" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1141" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1315" />
                    <RANKING order="2" place="2" resultid="1970" />
                    <RANKING order="3" place="3" resultid="1305" />
                    <RANKING order="4" place="4" resultid="1250" />
                    <RANKING order="5" place="5" resultid="1210" />
                    <RANKING order="6" place="6" resultid="1340" />
                    <RANKING order="7" place="7" resultid="1320" />
                    <RANKING order="8" place="8" resultid="1280" />
                    <RANKING order="9" place="8" resultid="1300" />
                    <RANKING order="10" place="10" resultid="1355" />
                    <RANKING order="11" place="11" resultid="1285" />
                    <RANKING order="12" place="12" resultid="1345" />
                    <RANKING order="13" place="12" resultid="1488" />
                    <RANKING order="14" place="14" resultid="1190" />
                    <RANKING order="15" place="15" resultid="1240" />
                    <RANKING order="16" place="16" resultid="1463" />
                    <RANKING order="17" place="17" resultid="1194" />
                    <RANKING order="18" place="18" resultid="1310" />
                    <RANKING order="19" place="19" resultid="1269" />
                    <RANKING order="20" place="20" resultid="1394" />
                    <RANKING order="21" place="21" resultid="2004" />
                    <RANKING order="22" place="22" resultid="2090" />
                    <RANKING order="23" place="23" resultid="2112" />
                    <RANKING order="24" place="24" resultid="1444" />
                    <RANKING order="25" place="25" resultid="1228" />
                    <RANKING order="26" place="26" resultid="2121" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2228" daytime="17:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2229" daytime="17:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2230" daytime="17:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2231" daytime="17:55" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2232" daytime="17:55" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2233" daytime="17:55" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2234" daytime="18:00" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="263" nation="BRA" region="PR" clubid="1270" swrid="75436" name="Clube Curitibano" shortname="Curitibano">
          <ATHLETES>
            <ATHLETE firstname="Rafael" lastname="Nishimura Ramina" birthdate="2013-11-25" gender="M" nation="BRA" license="376989" swrid="5588831" athleteid="1474" externalid="376989">
              <RESULTS>
                <RESULT eventid="1075" points="132" swimtime="00:00:46.18" resultid="1475" heatid="2151" lane="5" entrytime="00:00:47.09" entrycourse="LCM" />
                <RESULT eventid="1087" points="158" swimtime="00:03:08.46" resultid="1476" heatid="2169" lane="7" entrytime="00:03:07.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="162" swimtime="00:03:28.90" resultid="1477" heatid="2187" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="146" swimtime="00:00:39.66" resultid="1478" heatid="2231" lane="3" entrytime="00:00:38.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Massimo" lastname="Puppi Cardoso" birthdate="2015-03-30" gender="M" nation="BRA" license="406742" swrid="5717290" athleteid="1712" externalid="406742">
              <RESULTS>
                <RESULT eventid="1069" points="92" swimtime="00:00:57.41" resultid="1713" heatid="2142" lane="1" entrytime="00:00:58.44" entrycourse="LCM" />
                <RESULT eventid="1081" points="76" swimtime="00:00:55.49" resultid="1714" heatid="2159" lane="6" entrytime="00:00:59.33" entrycourse="LCM" />
                <RESULT eventid="1129" points="79" swimtime="00:00:48.63" resultid="1715" heatid="2214" lane="1" />
                <RESULT eventid="1109" points="54" swimtime="00:00:58.61" resultid="1716" heatid="2196" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Cavalcanti Breginski" birthdate="2016-04-06" gender="F" nation="BRA" license="415012" athleteid="1839" externalid="415012">
              <RESULTS>
                <RESULT eventid="1112" points="68" swimtime="00:01:05.62" resultid="1840" heatid="2200" lane="4" />
                <RESULT eventid="1132" points="43" swimtime="00:01:07.28" resultid="1841" heatid="2219" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Sieczkowski Pacheco" birthdate="2015-11-20" gender="F" nation="BRA" license="393261" swrid="5616450" athleteid="1627" externalid="393261">
              <RESULTS>
                <RESULT eventid="1066" points="124" swimtime="00:00:58.43" resultid="1628" heatid="2138" lane="3" entrytime="00:00:58.97" entrycourse="LCM" />
                <RESULT eventid="1078" points="128" swimtime="00:00:53.26" resultid="1629" heatid="2155" lane="7" entrytime="00:01:03.89" entrycourse="LCM" />
                <RESULT eventid="1106" points="80" swimtime="00:00:56.60" resultid="1630" heatid="2193" lane="8" entrytime="00:00:57.77" entrycourse="LCM" />
                <RESULT eventid="1126" points="116" swimtime="00:00:48.37" resultid="1631" heatid="2209" lane="4" entrytime="00:00:51.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Henrique Tiboni Araujo" birthdate="2013-06-11" gender="M" nation="BRA" license="376968" swrid="5588747" athleteid="1400" externalid="376968">
              <RESULTS>
                <RESULT eventid="1075" points="148" swimtime="00:00:44.50" resultid="1401" heatid="2151" lane="4" entrytime="00:00:45.70" entrycourse="LCM" />
                <RESULT eventid="1087" points="147" swimtime="00:03:13.18" resultid="1402" heatid="2168" lane="4" entrytime="00:03:30.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="139" swimtime="00:03:39.55" resultid="1403" heatid="2188" lane="2" entrytime="00:03:45.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="186" swimtime="00:00:36.57" resultid="1404" heatid="2231" lane="2" entrytime="00:00:38.57" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Cabrini Vieira" birthdate="2012-02-11" gender="F" nation="BRA" license="376961" swrid="5588571" athleteid="1381" externalid="376961">
              <RESULTS>
                <RESULT eventid="1084" points="421" swimtime="00:02:30.49" resultid="1382" heatid="2166" lane="1" entrytime="00:02:38.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="389" swimtime="00:00:36.77" resultid="1383" heatid="2148" lane="4" entrytime="00:00:35.22" entrycourse="LCM" />
                <RESULT eventid="1100" points="346" swimtime="00:02:59.49" resultid="1384" heatid="2182" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="453" swimtime="00:00:30.73" resultid="1385" heatid="2227" lane="4" entrytime="00:00:29.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="De Moraes" birthdate="2014-09-18" gender="M" nation="BRA" license="391024" swrid="5602529" athleteid="1577" externalid="391024">
              <RESULTS>
                <RESULT eventid="1069" points="116" swimtime="00:00:53.18" resultid="1578" heatid="2143" lane="5" entrytime="00:00:48.38" entrycourse="LCM" />
                <RESULT eventid="1093" points="233" swimtime="00:01:16.06" resultid="1579" heatid="2179" lane="3" entrytime="00:01:31.20" entrycourse="LCM" />
                <RESULT eventid="1129" points="239" swimtime="00:00:33.67" resultid="1580" heatid="2218" lane="5" entrytime="00:00:35.31" entrycourse="LCM" />
                <RESULT eventid="1109" points="151" swimtime="00:00:41.82" resultid="1581" heatid="2199" lane="3" entrytime="00:00:40.53" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Zagonel Krempel" birthdate="2015-07-27" gender="F" nation="BRA" license="406962" swrid="5717305" athleteid="1763" externalid="406962">
              <RESULTS>
                <RESULT eventid="1066" points="99" swimtime="00:01:02.90" resultid="1764" heatid="2137" lane="5" entrytime="00:01:06.98" entrycourse="LCM" />
                <RESULT eventid="1090" points="95" swimtime="00:01:53.28" resultid="1765" heatid="2173" lane="1" entrytime="00:02:15.15" entrycourse="LCM" />
                <RESULT comment="SW 8.3 - Movimento alternado das pernas ou pés.  (Horário: 16:29), Nadou livre." eventid="1106" status="DSQ" swimtime="00:00:48.22" resultid="1766" heatid="2192" lane="7" />
                <RESULT eventid="1126" points="122" swimtime="00:00:47.52" resultid="1767" heatid="2209" lane="7" entrytime="00:00:56.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Paulo Celles" birthdate="2016-09-07" gender="M" nation="BRA" license="411996" swrid="5740017" athleteid="1796" externalid="411996">
              <RESULTS>
                <RESULT eventid="1114" status="DNS" swimtime="00:00:00.00" resultid="1797" heatid="2201" lane="4" />
                <RESULT eventid="1134" status="DNS" swimtime="00:00:00.00" resultid="1798" heatid="2221" lane="5" entrytime="00:01:08.21" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Francia Soares" birthdate="2014-06-01" gender="F" nation="BRA" license="391011" swrid="5602540" athleteid="1543" externalid="391011">
              <RESULTS>
                <RESULT eventid="1078" status="DNS" swimtime="00:00:00.00" resultid="1544" heatid="2155" lane="5" entrytime="00:01:01.16" entrycourse="LCM" />
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="1545" heatid="2174" lane="5" entrytime="00:01:40.41" entrycourse="LCM" />
                <RESULT eventid="1126" status="DNS" swimtime="00:00:00.00" resultid="1546" heatid="2211" lane="2" entrytime="00:00:42.89" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Salomao" birthdate="2012-05-07" gender="M" nation="BRA" license="369261" swrid="5602581" athleteid="1281" externalid="369261">
              <RESULTS>
                <RESULT eventid="1075" points="200" swimtime="00:00:40.22" resultid="1282" heatid="2149" lane="3" />
                <RESULT eventid="1087" points="271" swimtime="00:02:37.54" resultid="1283" heatid="2171" lane="2" entrytime="00:02:37.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="186" swimtime="00:01:26.49" resultid="1284" heatid="2205" lane="2" entrytime="00:01:28.18" entrycourse="LCM" />
                <RESULT eventid="1139" points="254" swimtime="00:00:32.99" resultid="1285" heatid="2233" lane="4" entrytime="00:00:32.53" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Kraemer Geremia" birthdate="2013-08-16" gender="M" nation="BRA" license="377041" swrid="5588762" athleteid="1455" externalid="377041">
              <RESULTS>
                <RESULT eventid="1075" points="217" swimtime="00:00:39.13" resultid="1456" heatid="2153" lane="7" entrytime="00:00:39.11" entrycourse="LCM" />
                <RESULT eventid="1087" points="200" swimtime="00:02:54.15" resultid="1457" heatid="2170" lane="2" entrytime="00:02:50.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="199" swimtime="00:03:14.96" resultid="1458" heatid="2189" lane="8" entrytime="00:03:19.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="96" swimtime="00:01:47.74" resultid="1459" heatid="2204" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Jacob Brunetti" birthdate="2015-11-10" gender="M" nation="BRA" license="406837" swrid="5717274" athleteid="1752" externalid="406837" />
            <ATHLETE firstname="Giuliana" lastname="Sovierzoski Ferreira" birthdate="2015-01-20" gender="F" nation="BRA" license="397168" swrid="5641776" athleteid="1662" externalid="397168">
              <RESULTS>
                <RESULT eventid="1066" points="164" swimtime="00:00:53.18" resultid="1663" heatid="2139" lane="2" entrytime="00:00:53.15" entrycourse="LCM" />
                <RESULT eventid="1078" points="93" swimtime="00:00:59.15" resultid="1664" heatid="2155" lane="2" entrytime="00:01:03.14" entrycourse="LCM" />
                <RESULT eventid="1106" points="52" swimtime="00:01:05.04" resultid="1665" heatid="2191" lane="7" />
                <RESULT eventid="1126" points="102" swimtime="00:00:50.42" resultid="1666" heatid="2209" lane="8" entrytime="00:01:05.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Ribas Luz" birthdate="2015-02-05" gender="F" nation="BRA" license="406743" swrid="5717291" athleteid="1717" externalid="406743">
              <RESULTS>
                <RESULT eventid="1078" points="129" swimtime="00:00:53.10" resultid="1718" heatid="2156" lane="1" entrytime="00:00:57.53" entrycourse="LCM" />
                <RESULT eventid="1090" points="73" swimtime="00:02:03.20" resultid="1719" heatid="2173" lane="7" entrytime="00:02:06.25" entrycourse="LCM" />
                <RESULT eventid="1106" status="DNS" swimtime="00:00:00.00" resultid="1720" heatid="2191" lane="4" />
                <RESULT eventid="1126" status="DNS" swimtime="00:00:00.00" resultid="1721" heatid="2210" lane="8" entrytime="00:00:50.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Antunes Luzzi" birthdate="2014-02-14" gender="M" nation="BRA" license="391019" swrid="5602510" athleteid="1562" externalid="391019">
              <RESULTS>
                <RESULT eventid="1069" points="79" swimtime="00:01:00.39" resultid="1563" heatid="2141" lane="2" entrytime="00:01:02.04" entrycourse="LCM" />
                <RESULT eventid="1093" points="66" swimtime="00:01:55.59" resultid="1564" heatid="2178" lane="1" entrytime="00:01:55.23" entrycourse="LCM" />
                <RESULT eventid="1129" points="79" swimtime="00:00:48.58" resultid="1565" heatid="2214" lane="4" entrytime="00:00:55.78" entrycourse="LCM" />
                <RESULT eventid="1109" points="26" swimtime="00:01:14.38" resultid="1566" heatid="2197" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Cavalca Petraglia" birthdate="2015-08-06" gender="M" nation="BRA" license="397275" swrid="5641757" athleteid="1667" externalid="397275">
              <RESULTS>
                <RESULT eventid="1069" points="89" swimtime="00:00:58.10" resultid="1668" heatid="2141" lane="3" entrytime="00:01:01.63" entrycourse="LCM" />
                <RESULT eventid="1081" points="94" swimtime="00:00:51.74" resultid="1669" heatid="2160" lane="8" entrytime="00:00:53.65" entrycourse="LCM" />
                <RESULT eventid="1129" points="97" swimtime="00:00:45.43" resultid="1670" heatid="2213" lane="2" />
                <RESULT eventid="1109" points="68" swimtime="00:00:54.37" resultid="1671" heatid="2197" lane="5" entrytime="00:01:03.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Portes Fabiane" birthdate="2012-12-28" gender="M" nation="BRA" license="376983" swrid="5588864" athleteid="1440" externalid="376983">
              <RESULTS>
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada.  (Horário: 9:38), Após a volta dos 50m." eventid="1063" status="DSQ" swimtime="00:02:05.77" resultid="1441" heatid="2134" lane="2" entrytime="00:02:09.71" entrycourse="LCM" />
                <RESULT eventid="1075" points="90" swimtime="00:00:52.42" resultid="1442" heatid="2150" lane="4" entrytime="00:00:55.83" entrycourse="LCM" />
                <RESULT eventid="1103" points="109" swimtime="00:03:57.96" resultid="1443" heatid="2188" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:01.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="102" swimtime="00:00:44.68" resultid="1444" heatid="2230" lane="7" entrytime="00:00:44.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Szpak Zraik" birthdate="2015-04-10" gender="M" nation="BRA" license="393259" swrid="5616451" athleteid="1617" externalid="393259">
              <RESULTS>
                <RESULT eventid="1069" points="155" swimtime="00:00:48.23" resultid="1618" heatid="2143" lane="2" entrytime="00:00:50.96" entrycourse="LCM" />
                <RESULT eventid="1093" points="123" swimtime="00:01:34.20" resultid="1619" heatid="2178" lane="4" entrytime="00:01:41.34" entrycourse="LCM" />
                <RESULT eventid="1129" points="135" swimtime="00:00:40.69" resultid="1620" heatid="2215" lane="5" entrytime="00:00:46.28" entrycourse="LCM" />
                <RESULT eventid="1109" points="98" swimtime="00:00:48.16" resultid="1621" heatid="2196" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Cury Abreu" birthdate="2013-05-17" gender="F" nation="BRA" license="376974" swrid="5588614" athleteid="1410" externalid="376974">
              <RESULTS>
                <RESULT eventid="1084" status="DNS" swimtime="00:00:00.00" resultid="1411" heatid="2164" lane="2" entrytime="00:03:07.79" entrycourse="LCM" />
                <RESULT eventid="1072" status="DNS" swimtime="00:00:00.00" resultid="1412" heatid="2148" lane="7" entrytime="00:00:39.41" entrycourse="LCM" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 15:58), Virada dos 150M." eventid="1100" status="DSQ" swimtime="00:03:16.73" resultid="1413" heatid="2184" lane="1" entrytime="00:03:40.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="378" swimtime="00:00:32.65" resultid="1414" heatid="2226" lane="3" entrytime="00:00:33.59" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Alice Silva Gomes Xavier" birthdate="2013-02-25" gender="F" nation="BRA" license="371040" swrid="5717241" athleteid="1753" externalid="371040">
              <RESULTS>
                <RESULT eventid="1060" points="262" swimtime="00:01:40.20" resultid="1754" heatid="2131" lane="7" entrytime="00:01:36.52" entrycourse="LCM" />
                <RESULT eventid="1084" points="334" swimtime="00:02:42.63" resultid="1755" heatid="2165" lane="4" entrytime="00:02:47.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="282" swimtime="00:03:12.23" resultid="1756" heatid="2182" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="364" swimtime="00:00:33.06" resultid="1757" heatid="2227" lane="8" entrytime="00:00:32.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Rampazzo" birthdate="2013-02-18" gender="M" nation="BRA" license="400269" swrid="5748679" athleteid="1817" externalid="400269">
              <RESULTS>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 9:34)" eventid="1063" status="DSQ" swimtime="00:01:36.01" resultid="1818" heatid="2133" lane="6" />
                <RESULT eventid="1087" points="196" swimtime="00:02:55.55" resultid="1819" heatid="2168" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="211" swimtime="00:03:11.32" resultid="1820" heatid="2187" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="237" swimtime="00:00:33.76" resultid="1821" heatid="2229" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="De Lima Cavalcanti" birthdate="2014-10-07" gender="M" nation="BRA" license="385884" swrid="5684550" athleteid="1702" externalid="385884">
              <RESULTS>
                <RESULT eventid="1081" points="194" swimtime="00:00:40.63" resultid="1703" heatid="2161" lane="5" entrytime="00:00:43.07" entrycourse="LCM" />
                <RESULT eventid="1093" points="180" swimtime="00:01:22.99" resultid="1704" heatid="2180" lane="3" entrytime="00:01:24.01" entrycourse="LCM" />
                <RESULT eventid="1129" points="172" swimtime="00:00:37.56" resultid="1705" heatid="2217" lane="4" entrytime="00:00:37.98" entrycourse="LCM" />
                <RESULT eventid="1109" points="134" swimtime="00:00:43.46" resultid="1706" heatid="2199" lane="8" entrytime="00:00:48.94" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Antunes Saboia" birthdate="2012-06-28" gender="M" nation="BRA" license="369278" swrid="5602511" athleteid="1336" externalid="369278">
              <RESULTS>
                <RESULT eventid="1063" points="240" swimtime="00:01:31.43" resultid="1337" heatid="2135" lane="3" entrytime="00:01:30.44" entrycourse="LCM" />
                <RESULT eventid="1087" points="266" swimtime="00:02:38.53" resultid="1338" heatid="2170" lane="4" entrytime="00:02:41.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="240" swimtime="00:03:03.41" resultid="1339" heatid="2189" lane="5" entrytime="00:02:57.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="276" swimtime="00:00:32.09" resultid="1340" heatid="2233" lane="5" entrytime="00:00:32.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olavo" lastname="Valduga Artigas" birthdate="2012-06-26" gender="M" nation="BRA" license="369270" swrid="5588941" athleteid="1306" externalid="369270">
              <RESULTS>
                <RESULT eventid="1063" points="167" swimtime="00:01:43.24" resultid="1307" heatid="2135" lane="1" entrytime="00:01:44.16" entrycourse="LCM" />
                <RESULT eventid="1075" points="150" swimtime="00:00:44.28" resultid="1308" heatid="2152" lane="8" entrytime="00:00:45.41" entrycourse="LCM" />
                <RESULT eventid="1103" points="216" swimtime="00:03:09.83" resultid="1309" heatid="2188" lane="4" entrytime="00:03:21.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="203" swimtime="00:00:35.57" resultid="1310" heatid="2229" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Vian" birthdate="2014-03-25" gender="F" nation="BRA" license="393919" swrid="5641779" athleteid="1652" externalid="393919">
              <RESULTS>
                <RESULT eventid="1078" points="202" swimtime="00:00:45.73" resultid="1653" heatid="2157" lane="6" entrytime="00:00:48.38" entrycourse="LCM" />
                <RESULT eventid="1090" points="154" swimtime="00:01:36.42" resultid="1654" heatid="2174" lane="4" entrytime="00:01:39.69" entrycourse="LCM" />
                <RESULT eventid="1106" points="131" swimtime="00:00:48.00" resultid="1655" heatid="2194" lane="1" entrytime="00:00:50.48" entrycourse="LCM" />
                <RESULT eventid="1126" points="196" swimtime="00:00:40.63" resultid="1656" heatid="2212" lane="8" entrytime="00:00:41.27" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Baptistella" birthdate="2013-01-23" gender="M" nation="BRA" license="391152" swrid="5602545" athleteid="1602" externalid="391152">
              <RESULTS>
                <RESULT eventid="1075" points="231" swimtime="00:00:38.34" resultid="1603" heatid="2152" lane="4" entrytime="00:00:40.34" entrycourse="LCM" />
                <RESULT eventid="1087" points="228" swimtime="00:02:46.93" resultid="1604" heatid="2169" lane="1" entrytime="00:03:12.28" entrycourse="LCM" />
                <RESULT eventid="1103" points="210" swimtime="00:03:11.74" resultid="1605" heatid="2188" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="245" swimtime="00:00:33.39" resultid="1606" heatid="2231" lane="6" entrytime="00:00:38.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Pisani Ferreira" birthdate="2014-01-26" gender="M" nation="BRA" license="391017" swrid="5602570" athleteid="1552" externalid="391017">
              <RESULTS>
                <RESULT eventid="1069" points="134" swimtime="00:00:50.61" resultid="1553" heatid="2142" lane="7" entrytime="00:00:57.70" entrycourse="LCM" />
                <RESULT eventid="1093" points="117" swimtime="00:01:35.60" resultid="1554" heatid="2176" lane="3" />
                <RESULT eventid="1129" points="138" swimtime="00:00:40.45" resultid="1555" heatid="2213" lane="1" />
                <RESULT eventid="1109" points="75" swimtime="00:00:52.70" resultid="1556" heatid="2198" lane="7" entrytime="00:00:59.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Schmidt Wozniaki" birthdate="2012-07-07" gender="M" nation="BRA" license="376963" swrid="5588905" athleteid="1391" externalid="376963">
              <RESULTS>
                <RESULT eventid="1063" points="128" swimtime="00:01:52.82" resultid="1392" heatid="2134" lane="3" entrytime="00:02:00.95" entrycourse="LCM" />
                <RESULT eventid="1075" points="109" swimtime="00:00:49.23" resultid="1393" heatid="2151" lane="2" entrytime="00:00:48.38" entrycourse="LCM" />
                <RESULT eventid="1139" points="181" swimtime="00:00:36.92" resultid="1394" heatid="2231" lane="7" entrytime="00:00:38.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Pisani Ferreira" birthdate="2012-08-06" gender="F" nation="BRA" license="376985" swrid="5588862" athleteid="1489" externalid="376985">
              <RESULTS>
                <RESULT eventid="1060" points="238" swimtime="00:01:43.44" resultid="1490" heatid="2130" lane="3" entrytime="00:01:46.43" entrycourse="LCM" />
                <RESULT eventid="1072" points="153" swimtime="00:00:50.18" resultid="1491" heatid="2145" lane="6" entrytime="00:00:53.56" entrycourse="LCM" />
                <RESULT eventid="1100" points="189" swimtime="00:03:39.41" resultid="1492" heatid="2182" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="231" swimtime="00:00:38.45" resultid="1493" heatid="2224" lane="3" entrytime="00:00:40.19" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Steven" lastname="Matheussi Viana E Silva" birthdate="2012-05-03" gender="M" nation="BRA" license="376986" swrid="5588810" athleteid="1484" externalid="376986">
              <RESULTS>
                <RESULT eventid="1063" points="234" swimtime="00:01:32.19" resultid="1485" heatid="2135" lane="6" entrytime="00:01:33.25" entrycourse="LCM" />
                <RESULT eventid="1087" points="249" swimtime="00:02:42.01" resultid="1486" heatid="2169" lane="4" entrytime="00:02:59.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="183" swimtime="00:01:27.05" resultid="1487" heatid="2205" lane="6" entrytime="00:01:25.23" entrycourse="LCM" />
                <RESULT eventid="1139" points="241" swimtime="00:00:33.57" resultid="1488" heatid="2230" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Ruschka Druszcz" birthdate="2016-05-09" gender="F" nation="BRA" license="412025" swrid="5740018" athleteid="1814" externalid="412025">
              <RESULTS>
                <RESULT eventid="1122" status="DNS" swimtime="00:00:00.00" resultid="1815" heatid="2206" lane="4" entrytime="00:01:06.26" entrycourse="LCM" />
                <RESULT eventid="1132" status="DNS" swimtime="00:00:00.00" resultid="1816" heatid="2220" lane="5" entrytime="00:00:52.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Spadari Soso" birthdate="2012-12-28" gender="F" nation="BRA" license="377313" swrid="5588921" athleteid="1742" externalid="377313">
              <RESULTS>
                <RESULT eventid="1060" points="290" swimtime="00:01:36.88" resultid="1743" heatid="2131" lane="1" entrytime="00:01:37.26" entrycourse="LCM" />
                <RESULT eventid="1084" points="372" swimtime="00:02:36.85" resultid="1744" heatid="2166" lane="2" entrytime="00:02:32.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.94" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 6.2 - Deixou a posição de costas, exceto ao executar uma virada.  (Horário: 15:48)" eventid="1100" status="DSQ" swimtime="00:03:06.41" resultid="1745" heatid="2182" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="374" swimtime="00:00:32.76" resultid="1746" heatid="2227" lane="6" entrytime="00:00:31.53" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Alzamora Calado" birthdate="2013-04-26" gender="F" nation="BRA" license="376960" swrid="5588522" athleteid="1376" externalid="376960">
              <RESULTS>
                <RESULT eventid="1060" points="259" swimtime="00:01:40.49" resultid="1377" heatid="2130" lane="4" entrytime="00:01:43.65" entrycourse="LCM" />
                <RESULT eventid="1084" points="288" swimtime="00:02:50.88" resultid="1378" heatid="2164" lane="4" entrytime="00:03:01.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="260" swimtime="00:03:17.46" resultid="1379" heatid="2184" lane="6" entrytime="00:03:29.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="373" swimtime="00:00:32.78" resultid="1380" heatid="2225" lane="5" entrytime="00:00:35.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia" lastname="Ziliotto Mehl" birthdate="2015-10-09" gender="F" nation="BRA" license="400122" swrid="5652905" athleteid="1692" externalid="400122">
              <RESULTS>
                <RESULT eventid="1066" points="126" swimtime="00:00:58.04" resultid="1693" heatid="2138" lane="6" entrytime="00:00:59.69" entrycourse="LCM" />
                <RESULT eventid="1090" points="174" swimtime="00:01:32.61" resultid="1694" heatid="2172" lane="3" />
                <RESULT eventid="1106" points="64" swimtime="00:01:00.91" resultid="1695" heatid="2192" lane="4" entrytime="00:00:59.52" entrycourse="LCM" />
                <RESULT eventid="1126" points="193" swimtime="00:00:40.85" resultid="1696" heatid="2211" lane="3" entrytime="00:00:42.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Albuquerque" birthdate="2012-11-16" gender="F" nation="BRA" license="369281" swrid="5602506" athleteid="1346" externalid="369281">
              <RESULTS>
                <RESULT eventid="1060" points="313" swimtime="00:01:34.38" resultid="1347" heatid="2131" lane="5" entrytime="00:01:35.21" entrycourse="LCM" />
                <RESULT eventid="1072" points="289" swimtime="00:00:40.59" resultid="1348" heatid="2144" lane="5" />
                <RESULT eventid="1100" points="331" swimtime="00:03:02.27" resultid="1349" heatid="2185" lane="3" entrytime="00:02:59.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="244" swimtime="00:01:28.70" resultid="1350" heatid="2203" lane="3" entrytime="00:01:25.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Hyczy Sarraff" birthdate="2016-12-22" gender="M" nation="BRA" license="415013" athleteid="1842" externalid="415013">
              <RESULTS>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="1843" heatid="2207" lane="6" />
                <RESULT eventid="1134" status="DNS" swimtime="00:00:00.00" resultid="1844" heatid="2221" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Della Villa Yang" birthdate="2015-02-27" gender="F" nation="BRA" license="393283" swrid="5616442" athleteid="1647" externalid="393283">
              <RESULTS>
                <RESULT eventid="1078" points="156" swimtime="00:00:49.86" resultid="1648" heatid="2156" lane="7" entrytime="00:00:56.74" entrycourse="LCM" />
                <RESULT eventid="1090" points="172" swimtime="00:01:32.86" resultid="1649" heatid="2172" lane="2" />
                <RESULT eventid="1106" points="98" swimtime="00:00:52.90" resultid="1650" heatid="2194" lane="8" entrytime="00:00:51.17" entrycourse="LCM" />
                <RESULT eventid="1126" points="177" swimtime="00:00:41.98" resultid="1651" heatid="2211" lane="7" entrytime="00:00:43.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Morais Shibata" birthdate="2014-02-09" gender="M" nation="BRA" license="391018" swrid="5602561" athleteid="1557" externalid="391018">
              <RESULTS>
                <RESULT eventid="1069" points="122" swimtime="00:00:52.29" resultid="1558" heatid="2143" lane="1" entrytime="00:00:53.07" entrycourse="LCM" />
                <RESULT eventid="1081" points="140" swimtime="00:00:45.33" resultid="1559" heatid="2161" lane="2" entrytime="00:00:46.77" entrycourse="LCM" />
                <RESULT eventid="1129" points="133" swimtime="00:00:40.94" resultid="1560" heatid="2216" lane="4" entrytime="00:00:41.57" entrycourse="LCM" />
                <RESULT eventid="1109" points="81" swimtime="00:00:51.43" resultid="1561" heatid="2198" lane="1" entrytime="00:00:59.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Felipe Canalli" birthdate="2015-12-23" gender="M" nation="BRA" license="406749" swrid="5717261" athleteid="1732" externalid="406749">
              <RESULTS>
                <RESULT eventid="1069" points="131" swimtime="00:00:51.04" resultid="1733" heatid="2142" lane="2" entrytime="00:00:55.85" entrycourse="LCM" />
                <RESULT eventid="1093" points="64" swimtime="00:01:56.69" resultid="1734" heatid="2177" lane="5" entrytime="00:02:07.81" entrycourse="LCM" />
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="1735" heatid="2213" lane="7" />
                <RESULT eventid="1109" points="64" swimtime="00:00:55.46" resultid="1736" heatid="2198" lane="2" entrytime="00:00:58.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Moreira Pasqual" birthdate="2014-07-09" gender="M" nation="BRA" license="382125" swrid="5602562" athleteid="1514" externalid="382125">
              <RESULTS>
                <RESULT eventid="1081" points="142" swimtime="00:00:45.06" resultid="1515" heatid="2161" lane="1" entrytime="00:00:47.60" entrycourse="LCM" />
                <RESULT eventid="1093" points="187" swimtime="00:01:21.85" resultid="1516" heatid="2178" lane="5" entrytime="00:01:41.44" entrycourse="LCM" />
                <RESULT eventid="1129" points="183" swimtime="00:00:36.81" resultid="1517" heatid="2216" lane="3" entrytime="00:00:42.35" entrycourse="LCM" />
                <RESULT eventid="1109" points="163" swimtime="00:00:40.70" resultid="1518" heatid="2198" lane="6" entrytime="00:00:55.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Da Cunha Souza" birthdate="2015-05-30" gender="F" nation="BRA" license="400016" swrid="5652883" athleteid="1687" externalid="400016">
              <RESULTS>
                <RESULT eventid="1078" points="202" swimtime="00:00:45.72" resultid="1688" heatid="2157" lane="8" entrytime="00:00:50.51" entrycourse="LCM" />
                <RESULT eventid="1090" points="150" swimtime="00:01:37.30" resultid="1689" heatid="2174" lane="6" entrytime="00:01:44.00" entrycourse="LCM" />
                <RESULT eventid="1106" points="102" swimtime="00:00:52.13" resultid="1690" heatid="2192" lane="3" entrytime="00:01:05.59" entrycourse="LCM" />
                <RESULT eventid="1126" points="153" swimtime="00:00:44.14" resultid="1691" heatid="2211" lane="1" entrytime="00:00:44.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Gonçalves Sperandio" birthdate="2013-05-22" gender="M" nation="BRA" license="376980" swrid="5588851" athleteid="1425" externalid="376980">
              <RESULTS>
                <RESULT eventid="1063" points="176" swimtime="00:01:41.41" resultid="1426" heatid="2132" lane="4" />
                <RESULT eventid="1087" points="246" swimtime="00:02:42.71" resultid="1427" heatid="2170" lane="6" entrytime="00:02:48.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="222" swimtime="00:03:08.03" resultid="1428" heatid="2189" lane="1" entrytime="00:03:16.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="241" swimtime="00:00:33.59" resultid="1429" heatid="2233" lane="8" entrytime="00:00:35.05" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Bernardi Pedrosa" birthdate="2013-03-09" gender="F" nation="BRA" license="376977" swrid="5588551" athleteid="1420" externalid="376977">
              <RESULTS>
                <RESULT eventid="1084" points="255" swimtime="00:02:57.92" resultid="1421" heatid="2163" lane="5" entrytime="00:03:30.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="293" swimtime="00:00:40.43" resultid="1422" heatid="2147" lane="3" entrytime="00:00:42.24" entrycourse="LCM" />
                <RESULT eventid="1100" points="216" swimtime="00:03:29.98" resultid="1423" heatid="2183" lane="5" entrytime="00:04:09.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="303" swimtime="00:00:35.14" resultid="1424" heatid="2225" lane="6" entrytime="00:00:36.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Liam" lastname="Batista Grise" birthdate="2014-03-27" gender="M" nation="BRA" license="391008" swrid="5602514" athleteid="1539" externalid="391008">
              <RESULTS>
                <RESULT eventid="1069" status="DNS" swimtime="00:00:00.00" resultid="1540" heatid="2142" lane="4" entrytime="00:00:54.92" entrycourse="LCM" />
                <RESULT eventid="1093" status="DNS" swimtime="00:00:00.00" resultid="1541" heatid="2178" lane="3" entrytime="00:01:43.84" entrycourse="LCM" />
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="1542" heatid="2216" lane="7" entrytime="00:00:43.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enrico" lastname="Calixto Rauen" birthdate="2016-06-25" gender="M" nation="BRA" license="415011" athleteid="1836" externalid="415011">
              <RESULTS>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="1837" heatid="2207" lane="5" />
                <RESULT eventid="1134" points="36" swimtime="00:01:02.99" resultid="1838" heatid="2221" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Albuquerque" birthdate="2012-08-17" gender="F" nation="BRA" license="369275" swrid="5602507" athleteid="1321" externalid="369275">
              <RESULTS>
                <RESULT eventid="1060" points="431" swimtime="00:01:24.87" resultid="1322" heatid="2131" lane="4" entrytime="00:01:25.83" entrycourse="LCM" />
                <RESULT eventid="1084" points="247" swimtime="00:02:59.66" resultid="1323" heatid="2164" lane="5" entrytime="00:03:02.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="294" swimtime="00:03:09.55" resultid="1324" heatid="2185" lane="2" entrytime="00:03:06.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="344" swimtime="00:00:33.68" resultid="1325" heatid="2226" lane="5" entrytime="00:00:33.21" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Prosdocimo" birthdate="2012-11-30" gender="M" nation="BRA" license="369272" swrid="5602575" athleteid="1316" externalid="369272">
              <RESULTS>
                <RESULT eventid="1075" points="270" swimtime="00:00:36.42" resultid="1317" heatid="2153" lane="6" entrytime="00:00:38.33" entrycourse="LCM" />
                <RESULT eventid="1087" points="272" swimtime="00:02:37.30" resultid="1318" heatid="2171" lane="3" entrytime="00:02:36.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="145" swimtime="00:01:33.99" resultid="1319" heatid="2204" lane="1" />
                <RESULT eventid="1139" points="270" swimtime="00:00:32.35" resultid="1320" heatid="2234" lane="8" entrytime="00:00:32.53" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="De Almeida Dias" birthdate="2012-02-18" gender="F" nation="BRA" license="369262" swrid="5588638" athleteid="1286" externalid="369262">
              <RESULTS>
                <RESULT eventid="1060" points="362" swimtime="00:01:29.96" resultid="1287" heatid="2131" lane="8" entrytime="00:01:37.88" entrycourse="LCM" />
                <RESULT eventid="1084" points="476" swimtime="00:02:24.47" resultid="1288" heatid="2166" lane="5" entrytime="00:02:27.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="377" swimtime="00:02:54.57" resultid="1289" heatid="2185" lane="6" entrytime="00:03:03.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="421" swimtime="00:00:31.48" resultid="1290" heatid="2227" lane="3" entrytime="00:00:30.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Hadad" birthdate="2015-09-09" gender="M" nation="BRA" license="406740" swrid="5717272" athleteid="1707" externalid="406740">
              <RESULTS>
                <RESULT eventid="1081" points="61" swimtime="00:00:59.70" resultid="1708" heatid="2159" lane="1" entrytime="00:01:03.66" entrycourse="LCM" />
                <RESULT eventid="1093" points="90" swimtime="00:01:44.33" resultid="1709" heatid="2178" lane="8" entrytime="00:01:55.31" entrycourse="LCM" />
                <RESULT eventid="1129" points="75" swimtime="00:00:49.42" resultid="1710" heatid="2213" lane="4" />
                <RESULT eventid="1109" points="55" swimtime="00:00:58.39" resultid="1711" heatid="2195" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enrico" lastname="Hallage Bianchini" birthdate="2014-02-27" gender="M" nation="BRA" license="397164" swrid="5661348" athleteid="1657" externalid="397164">
              <RESULTS>
                <RESULT eventid="1081" points="165" swimtime="00:00:42.93" resultid="1658" heatid="2161" lane="7" entrytime="00:00:46.80" entrycourse="LCM" />
                <RESULT eventid="1093" points="224" swimtime="00:01:17.14" resultid="1659" heatid="2180" lane="7" entrytime="00:01:27.47" entrycourse="LCM" />
                <RESULT eventid="1129" points="205" swimtime="00:00:35.44" resultid="1660" heatid="2216" lane="5" entrytime="00:00:41.93" entrycourse="LCM" />
                <RESULT eventid="1109" points="130" swimtime="00:00:43.86" resultid="1661" heatid="2199" lane="1" entrytime="00:00:47.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Saporiti Salvi" birthdate="2013-06-28" gender="M" nation="BRA" license="377032" swrid="5588896" athleteid="1450" externalid="377032">
              <RESULTS>
                <RESULT eventid="1063" points="143" swimtime="00:01:48.69" resultid="1451" heatid="2132" lane="3" />
                <RESULT eventid="1087" points="219" swimtime="00:02:49.12" resultid="1452" heatid="2170" lane="5" entrytime="00:02:45.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="205" swimtime="00:03:13.10" resultid="1453" heatid="2189" lane="3" entrytime="00:03:10.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="147" swimtime="00:01:33.65" resultid="1454" heatid="2205" lane="1" entrytime="00:01:29.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Bittencourt Ribas" birthdate="2013-02-01" gender="F" nation="BRA" license="372682" swrid="5588555" athleteid="1361" externalid="372682">
              <RESULTS>
                <RESULT eventid="1084" points="316" swimtime="00:02:45.58" resultid="1362" heatid="2165" lane="2" entrytime="00:02:52.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="315" swimtime="00:00:39.44" resultid="1363" heatid="2148" lane="8" entrytime="00:00:40.35" entrycourse="LCM" />
                <RESULT eventid="1100" points="311" swimtime="00:03:06.10" resultid="1364" heatid="2184" lane="5" entrytime="00:03:13.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="342" swimtime="00:00:33.75" resultid="1365" heatid="2226" lane="8" entrytime="00:00:34.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Xavier Jardim" birthdate="2012-01-23" gender="M" nation="BRA" license="369259" swrid="5641781" athleteid="1276" externalid="369259">
              <RESULTS>
                <RESULT eventid="1063" points="170" swimtime="00:01:42.62" resultid="1277" heatid="2133" lane="4" />
                <RESULT eventid="1087" points="252" swimtime="00:02:41.48" resultid="1278" heatid="2171" lane="7" entrytime="00:02:38.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="148" swimtime="00:01:33.45" resultid="1279" heatid="2205" lane="8" entrytime="00:01:30.44" entrycourse="LCM" />
                <RESULT eventid="1139" points="259" swimtime="00:00:32.79" resultid="1280" heatid="2234" lane="7" entrytime="00:00:31.86" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ravi" lastname="Osternack Erbe" birthdate="2013-08-10" gender="M" nation="BRA" license="372681" swrid="5588841" athleteid="1356" externalid="372681">
              <RESULTS>
                <RESULT eventid="1075" points="208" swimtime="00:00:39.72" resultid="1357" heatid="2152" lane="2" entrytime="00:00:44.63" entrycourse="LCM" />
                <RESULT eventid="1087" points="249" swimtime="00:02:41.94" resultid="1358" heatid="2170" lane="8" entrytime="00:02:56.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="219" swimtime="00:03:09.11" resultid="1359" heatid="2188" lane="3" entrytime="00:03:25.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="154" swimtime="00:01:32.22" resultid="1360" heatid="2204" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Menezes" birthdate="2015-07-28" gender="F" nation="BRA" license="412898" athleteid="1822" externalid="412898">
              <RESULTS>
                <RESULT eventid="1078" points="102" swimtime="00:00:57.43" resultid="1823" heatid="2154" lane="5" />
                <RESULT eventid="1090" points="91" swimtime="00:01:54.72" resultid="1824" heatid="2172" lane="5" />
                <RESULT eventid="1126" points="125" swimtime="00:00:47.17" resultid="1825" heatid="2208" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Afonso Fowler" birthdate="2014-01-22" gender="M" nation="BRA" license="393264" swrid="5661338" athleteid="1642" externalid="393264">
              <RESULTS>
                <RESULT eventid="1081" status="DNS" swimtime="00:00:00.00" resultid="1643" heatid="2160" lane="5" entrytime="00:00:49.09" entrycourse="LCM" />
                <RESULT eventid="1093" status="DNS" swimtime="00:00:00.00" resultid="1644" heatid="2179" lane="1" entrytime="00:01:36.96" entrycourse="LCM" />
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="1645" heatid="2218" lane="8" entrytime="00:00:37.78" entrycourse="LCM" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="1646" heatid="2198" lane="3" entrytime="00:00:52.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Guimaraes Mesquita" birthdate="2013-12-30" gender="F" nation="BRA" license="391027" swrid="5602544" athleteid="1592" externalid="391027">
              <RESULTS>
                <RESULT eventid="1060" points="168" swimtime="00:01:56.13" resultid="1593" heatid="2130" lane="6" entrytime="00:01:51.97" entrycourse="LCM" />
                <RESULT eventid="1084" points="189" swimtime="00:03:16.38" resultid="1594" heatid="2162" lane="5" />
                <RESULT eventid="1100" points="191" swimtime="00:03:38.73" resultid="1595" heatid="2184" lane="8" entrytime="00:04:06.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:53.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="199" swimtime="00:00:40.40" resultid="1596" heatid="2223" lane="4" entrytime="00:00:42.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Almeida Jorge" birthdate="2015-05-27" gender="M" nation="BRA" license="406836" swrid="5717242" athleteid="1747" externalid="406836">
              <RESULTS>
                <RESULT eventid="1069" points="70" swimtime="00:01:02.73" resultid="1748" heatid="2141" lane="7" entrytime="00:01:04.95" entrycourse="LCM" />
                <RESULT eventid="1081" points="70" swimtime="00:00:56.88" resultid="1749" heatid="2159" lane="3" entrytime="00:00:58.23" entrycourse="LCM" />
                <RESULT eventid="1129" points="38" swimtime="00:01:02.00" resultid="1750" heatid="2214" lane="6" entrytime="00:01:03.14" entrycourse="LCM" />
                <RESULT eventid="1109" points="35" swimtime="00:01:07.45" resultid="1751" heatid="2197" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Simioni Albuquerque" birthdate="2014-12-23" gender="F" nation="BRA" license="401980" swrid="5661355" athleteid="1697" externalid="401980">
              <RESULTS>
                <RESULT eventid="1066" points="150" swimtime="00:00:54.85" resultid="1698" heatid="2138" lane="8" entrytime="00:01:05.71" entrycourse="LCM" />
                <RESULT eventid="1090" points="186" swimtime="00:01:30.45" resultid="1699" heatid="2173" lane="4" entrytime="00:01:52.63" entrycourse="LCM" />
                <RESULT eventid="1106" points="184" swimtime="00:00:42.95" resultid="1700" heatid="2190" lane="5" />
                <RESULT eventid="1126" points="232" swimtime="00:00:38.39" resultid="1701" heatid="2210" lane="2" entrytime="00:00:45.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Fonseca Ribeiro" birthdate="2016-02-25" gender="F" nation="BRA" license="412016" swrid="5740011" athleteid="1811" externalid="412016">
              <RESULTS>
                <RESULT eventid="1122" points="76" swimtime="00:01:08.70" resultid="1812" heatid="2206" lane="3" entrytime="00:01:09.84" entrycourse="LCM" />
                <RESULT eventid="1132" points="84" swimtime="00:00:53.85" resultid="1813" heatid="2220" lane="6" entrytime="00:00:55.56" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Vianna Almeida" birthdate="2014-12-16" gender="M" nation="BRA" license="410292" swrid="5740019" athleteid="1791" externalid="410292">
              <RESULTS>
                <RESULT eventid="1069" points="109" swimtime="00:00:54.16" resultid="1792" heatid="2141" lane="6" entrytime="00:01:01.80" entrycourse="LCM" />
                <RESULT eventid="1081" points="91" swimtime="00:00:52.19" resultid="1793" heatid="2158" lane="1" />
                <RESULT eventid="1129" points="110" swimtime="00:00:43.60" resultid="1794" heatid="2215" lane="8" entrytime="00:00:50.79" entrycourse="LCM" />
                <RESULT eventid="1109" points="48" swimtime="00:01:00.87" resultid="1795" heatid="2197" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Alice Palhano" birthdate="2016-04-06" gender="F" nation="BRA" license="412015" swrid="5740004" athleteid="1808" externalid="412015">
              <RESULTS>
                <RESULT eventid="1112" points="48" swimtime="00:01:13.51" resultid="1809" heatid="2200" lane="5" />
                <RESULT eventid="1132" points="26" swimtime="00:01:18.80" resultid="1810" heatid="2220" lane="7" entrytime="00:01:10.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Schiavo Vianna" birthdate="2013-04-27" gender="F" nation="BRA" license="391005" swrid="5602582" athleteid="1529" externalid="391005">
              <RESULTS>
                <RESULT eventid="1060" points="187" swimtime="00:01:52.14" resultid="1530" heatid="2130" lane="2" entrytime="00:01:54.87" entrycourse="LCM" />
                <RESULT eventid="1084" points="194" swimtime="00:03:14.70" resultid="1531" heatid="2163" lane="7" entrytime="00:04:08.21" entrycourse="LCM" />
                <RESULT comment="SW 8.5 - Totalmente submerso durante o nado.  (Horário: 15:53)" eventid="1100" status="DSQ" swimtime="00:03:54.46" resultid="1532" heatid="2183" lane="6" entrytime="00:04:25.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:59.19" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 17:47)" eventid="1136" status="DSQ" swimtime="00:00:36.63" resultid="1533" heatid="2225" lane="8" entrytime="00:00:37.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Poletto Abrahao" birthdate="2014-10-20" gender="M" nation="BRA" license="382128" swrid="5602571" athleteid="1524" externalid="382128">
              <RESULTS>
                <RESULT eventid="1069" points="191" swimtime="00:00:45.02" resultid="1525" heatid="2143" lane="4" entrytime="00:00:44.75" entrycourse="LCM" />
                <RESULT eventid="1081" points="148" swimtime="00:00:44.51" resultid="1526" heatid="2160" lane="2" entrytime="00:00:50.37" entrycourse="LCM" />
                <RESULT eventid="1129" points="211" swimtime="00:00:35.10" resultid="1527" heatid="2217" lane="3" entrytime="00:00:39.24" entrycourse="LCM" />
                <RESULT eventid="1109" points="170" swimtime="00:00:40.17" resultid="1528" heatid="2199" lane="2" entrytime="00:00:45.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Caron Braga" birthdate="2016-02-01" gender="F" nation="BRA" license="415257" athleteid="1854" externalid="415257">
              <RESULTS>
                <RESULT eventid="1122" points="50" swimtime="00:01:18.72" resultid="1855" heatid="2206" lane="7" />
                <RESULT eventid="1132" points="39" swimtime="00:01:09.32" resultid="1856" heatid="2219" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Trevisan De Paula" birthdate="2014-01-27" gender="M" nation="BRA" license="377152" swrid="5602568" athleteid="1494" externalid="377152">
              <RESULTS>
                <RESULT eventid="1081" points="184" swimtime="00:00:41.35" resultid="1495" heatid="2161" lane="6" entrytime="00:00:43.99" entrycourse="LCM" />
                <RESULT eventid="1093" points="217" swimtime="00:01:17.90" resultid="1496" heatid="2180" lane="4" entrytime="00:01:19.00" entrycourse="LCM" />
                <RESULT eventid="1129" points="214" swimtime="00:00:34.93" resultid="1497" heatid="2218" lane="4" entrytime="00:00:33.59" entrycourse="LCM" />
                <RESULT eventid="1109" points="208" swimtime="00:00:37.55" resultid="1498" heatid="2199" lane="4" entrytime="00:00:39.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Mayer Paludetto" birthdate="2012-10-30" gender="F" nation="BRA" license="369264" swrid="5588811" athleteid="1291" externalid="369264">
              <RESULTS>
                <RESULT eventid="1060" points="309" swimtime="00:01:34.81" resultid="1292" heatid="2131" lane="3" entrytime="00:01:35.77" entrycourse="LCM" />
                <RESULT eventid="1084" points="431" swimtime="00:02:29.30" resultid="1293" heatid="2166" lane="6" entrytime="00:02:32.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="405" swimtime="00:02:50.40" resultid="1294" heatid="2185" lane="4" entrytime="00:02:53.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="435" swimtime="00:00:31.15" resultid="1295" heatid="2222" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Vanzo Assumpcao" birthdate="2012-05-15" gender="M" nation="BRA" license="369258" swrid="5588942" athleteid="1271" externalid="369258">
              <RESULTS>
                <RESULT eventid="1075" points="308" swimtime="00:00:34.85" resultid="1272" heatid="2153" lane="5" entrytime="00:00:36.26" entrycourse="LCM" />
                <RESULT eventid="1087" points="335" swimtime="00:02:26.86" resultid="1273" heatid="2167" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="304" swimtime="00:02:49.45" resultid="1274" heatid="2187" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="281" swimtime="00:01:15.41" resultid="1275" heatid="2205" lane="4" entrytime="00:01:18.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Carcereri Navarro" birthdate="2013-12-19" gender="M" nation="BRA" license="376962" swrid="5588576" athleteid="1386" externalid="376962">
              <RESULTS>
                <RESULT eventid="1063" points="177" swimtime="00:01:41.22" resultid="1387" heatid="2133" lane="2" />
                <RESULT eventid="1087" points="157" swimtime="00:03:08.98" resultid="1388" heatid="2168" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="158" swimtime="00:01:31.42" resultid="1389" heatid="2204" lane="4" entrytime="00:01:33.45" entrycourse="LCM" />
                <RESULT eventid="1139" points="190" swimtime="00:00:36.35" resultid="1390" heatid="2232" lane="6" entrytime="00:00:35.33" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="De Macedo Martynychen" birthdate="2015-06-12" gender="F" nation="BRA" license="399681" swrid="5652885" athleteid="1682" externalid="399681">
              <RESULTS>
                <RESULT eventid="1078" points="105" swimtime="00:00:56.76" resultid="1683" heatid="2155" lane="3" entrytime="00:01:02.12" entrycourse="LCM" />
                <RESULT eventid="1090" points="96" swimtime="00:01:52.64" resultid="1684" heatid="2173" lane="2" entrytime="00:02:05.97" entrycourse="LCM" />
                <RESULT eventid="1106" points="80" swimtime="00:00:56.52" resultid="1685" heatid="2192" lane="5" entrytime="00:00:59.53" entrycourse="LCM" />
                <RESULT eventid="1126" points="101" swimtime="00:00:50.61" resultid="1686" heatid="2208" lane="4" entrytime="00:01:06.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Pens Correa" birthdate="2015-11-27" gender="M" nation="BRA" license="393262" swrid="5616449" athleteid="1632" externalid="393262">
              <RESULTS>
                <RESULT eventid="1081" points="206" swimtime="00:00:39.86" resultid="1633" heatid="2161" lane="4" entrytime="00:00:41.28" entrycourse="LCM" />
                <RESULT eventid="1093" points="199" swimtime="00:01:20.13" resultid="1634" heatid="2177" lane="2" />
                <RESULT eventid="1129" points="213" swimtime="00:00:34.96" resultid="1635" heatid="2217" lane="6" entrytime="00:00:39.55" entrycourse="LCM" />
                <RESULT eventid="1109" points="190" swimtime="00:00:38.70" resultid="1636" heatid="2199" lane="5" entrytime="00:00:40.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Fernandes Tramujas" birthdate="2015-01-15" gender="F" nation="BRA" license="406750" swrid="5717263" athleteid="1737" externalid="406750">
              <RESULTS>
                <RESULT eventid="1066" points="65" swimtime="00:01:12.27" resultid="1738" heatid="2137" lane="7" entrytime="00:01:10.52" entrycourse="LCM" />
                <RESULT eventid="1090" points="103" swimtime="00:01:50.30" resultid="1739" heatid="2173" lane="5" entrytime="00:01:59.16" entrycourse="LCM" />
                <RESULT eventid="1106" points="44" swimtime="00:01:09.18" resultid="1740" heatid="2190" lane="4" />
                <RESULT eventid="1126" points="120" swimtime="00:00:47.76" resultid="1741" heatid="2208" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Betina" lastname="Vieira Pellanda" birthdate="2014-02-16" gender="F" nation="BRA" license="391041" swrid="5602589" athleteid="1597" externalid="391041">
              <RESULTS>
                <RESULT eventid="1078" points="185" swimtime="00:00:47.06" resultid="1598" heatid="2156" lane="4" entrytime="00:00:51.35" entrycourse="LCM" />
                <RESULT eventid="1090" points="186" swimtime="00:01:30.53" resultid="1599" heatid="2174" lane="3" entrytime="00:01:42.52" entrycourse="LCM" />
                <RESULT eventid="1106" points="110" swimtime="00:00:50.90" resultid="1600" heatid="2190" lane="3" />
                <RESULT eventid="1126" points="196" swimtime="00:00:40.60" resultid="1601" heatid="2211" lane="6" entrytime="00:00:42.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Shwetz Clivatti" birthdate="2015-03-05" gender="M" nation="BRA" license="406963" swrid="5717297" athleteid="1768" externalid="406963">
              <RESULTS>
                <RESULT eventid="1069" points="52" swimtime="00:01:09.43" resultid="1769" heatid="2141" lane="1" entrytime="00:01:16.70" entrycourse="LCM" />
                <RESULT eventid="1081" points="53" swimtime="00:01:02.66" resultid="1770" heatid="2158" lane="4" entrytime="00:01:05.36" entrycourse="LCM" />
                <RESULT eventid="1129" points="54" swimtime="00:00:55.30" resultid="1771" heatid="2214" lane="5" entrytime="00:00:58.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Rossi Mattioli" birthdate="2013-05-08" gender="F" nation="BRA" license="376988" swrid="5588892" athleteid="1479" externalid="376988">
              <RESULTS>
                <RESULT eventid="1084" points="255" swimtime="00:02:57.73" resultid="1480" heatid="2165" lane="1" entrytime="00:02:55.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="323" swimtime="00:00:39.12" resultid="1481" heatid="2147" lane="5" entrytime="00:00:40.94" entrycourse="LCM" />
                <RESULT eventid="1100" points="260" swimtime="00:03:17.50" resultid="1482" heatid="2183" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="314" swimtime="00:00:34.73" resultid="1483" heatid="2226" lane="7" entrytime="00:00:33.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Clara Prado Biscaia" birthdate="2013-10-24" gender="F" nation="BRA" license="391015" swrid="5602526" athleteid="1547" externalid="391015">
              <RESULTS>
                <RESULT eventid="1084" points="204" swimtime="00:03:11.44" resultid="1548" heatid="2163" lane="3" entrytime="00:03:33.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="183" swimtime="00:00:47.24" resultid="1549" heatid="2144" lane="4" />
                <RESULT eventid="1116" points="148" swimtime="00:01:44.76" resultid="1550" heatid="2203" lane="8" entrytime="00:01:43.45" entrycourse="LCM" />
                <RESULT eventid="1136" points="217" swimtime="00:00:39.28" resultid="1551" heatid="2224" lane="1" entrytime="00:00:42.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Viera Correa" birthdate="2012-03-07" gender="M" nation="BRA" license="369269" swrid="5602590" athleteid="1301" externalid="369269">
              <RESULTS>
                <RESULT eventid="1075" points="227" swimtime="00:00:38.56" resultid="1302" heatid="2153" lane="8" entrytime="00:00:39.83" entrycourse="LCM" />
                <RESULT eventid="1087" points="292" swimtime="00:02:33.70" resultid="1303" heatid="2171" lane="5" entrytime="00:02:32.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="251" swimtime="00:03:00.68" resultid="1304" heatid="2186" lane="5" />
                <RESULT eventid="1139" points="310" swimtime="00:00:30.87" resultid="1305" heatid="2234" lane="6" entrytime="00:00:31.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Garcia" birthdate="2015-10-26" gender="M" nation="BRA" license="406967" swrid="5717271" athleteid="1772" externalid="406967">
              <RESULTS>
                <RESULT eventid="1069" status="DNS" swimtime="00:00:00.00" resultid="1773" heatid="2140" lane="4" entrytime="00:01:27.24" entrycourse="LCM" />
                <RESULT eventid="1081" status="DNS" swimtime="00:00:00.00" resultid="1774" heatid="2159" lane="7" entrytime="00:01:03.30" entrycourse="LCM" />
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="1775" heatid="2214" lane="2" entrytime="00:01:08.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivia" lastname="Mayer Paludetto" birthdate="2016-04-01" gender="F" nation="BRA" license="412014" swrid="5740014" athleteid="1805" externalid="412014">
              <RESULTS>
                <RESULT eventid="1096" points="33" swimtime="00:01:15.73" resultid="1806" heatid="2181" lane="4" />
                <RESULT eventid="1132" points="86" swimtime="00:00:53.47" resultid="1807" heatid="2220" lane="4" entrytime="00:00:50.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Taborda Ribas" birthdate="2015-12-30" gender="M" nation="BRA" license="406748" swrid="5717299" athleteid="1727" externalid="406748">
              <RESULTS>
                <RESULT eventid="1081" points="67" swimtime="00:00:57.77" resultid="1728" heatid="2158" lane="7" />
                <RESULT eventid="1093" points="73" swimtime="00:01:52.11" resultid="1729" heatid="2178" lane="7" entrytime="00:01:55.17" entrycourse="LCM" />
                <RESULT eventid="1129" points="72" swimtime="00:00:50.21" resultid="1730" heatid="2215" lane="7" entrytime="00:00:49.17" entrycourse="LCM" />
                <RESULT eventid="1109" points="24" swimtime="00:01:16.34" resultid="1731" heatid="2197" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Toscani Kim" birthdate="2015-10-02" gender="F" nation="BRA" license="397276" swrid="5641778" athleteid="1672" externalid="397276">
              <RESULTS>
                <RESULT eventid="1066" points="189" swimtime="00:00:50.80" resultid="1673" heatid="2139" lane="6" entrytime="00:00:52.94" entrycourse="LCM" />
                <RESULT eventid="1090" points="158" swimtime="00:01:35.51" resultid="1674" heatid="2172" lane="7" />
                <RESULT eventid="1106" points="125" swimtime="00:00:48.82" resultid="1675" heatid="2193" lane="6" entrytime="00:00:54.59" entrycourse="LCM" />
                <RESULT eventid="1126" points="159" swimtime="00:00:43.58" resultid="1676" heatid="2210" lane="5" entrytime="00:00:44.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Marie Silva" birthdate="2014-08-24" gender="F" nation="BRA" license="391025" swrid="5602556" athleteid="1582" externalid="391025">
              <RESULTS>
                <RESULT eventid="1066" status="DNS" swimtime="00:00:00.00" resultid="1583" heatid="2138" lane="2" entrytime="00:01:00.06" entrycourse="LCM" />
                <RESULT eventid="1090" status="DNS" swimtime="00:00:00.00" resultid="1584" heatid="2175" lane="6" entrytime="00:01:31.58" entrycourse="LCM" />
                <RESULT eventid="1106" status="DNS" swimtime="00:00:00.00" resultid="1585" heatid="2194" lane="2" entrytime="00:00:49.69" entrycourse="LCM" />
                <RESULT eventid="1126" status="DNS" swimtime="00:00:00.00" resultid="1586" heatid="2208" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Andrade Vosgerau" birthdate="2016-02-16" gender="F" nation="BRA" license="415010" athleteid="1833" externalid="415010">
              <RESULTS>
                <RESULT eventid="1112" points="54" swimtime="00:01:11.06" resultid="1834" heatid="2200" lane="3" />
                <RESULT eventid="1122" points="56" swimtime="00:01:15.80" resultid="1835" heatid="2206" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Hallage Papp" birthdate="2012-07-02" gender="M" nation="BRA" license="377042" swrid="5588736" athleteid="1460" externalid="377042">
              <RESULTS>
                <RESULT eventid="1063" points="122" swimtime="00:01:54.40" resultid="1461" heatid="2134" lane="5" entrytime="00:01:59.69" entrycourse="LCM" />
                <RESULT eventid="1075" points="150" swimtime="00:00:44.32" resultid="1462" heatid="2152" lane="7" entrytime="00:00:44.87" entrycourse="LCM" />
                <RESULT eventid="1139" points="211" swimtime="00:00:35.12" resultid="1463" heatid="2232" lane="4" entrytime="00:00:35.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Guimaraes Mesquita" birthdate="2015-10-05" gender="F" nation="BRA" license="393263" swrid="5616444" athleteid="1637" externalid="393263">
              <RESULTS>
                <RESULT eventid="1066" status="DNS" swimtime="00:00:00.00" resultid="1638" heatid="2137" lane="6" entrytime="00:01:10.17" entrycourse="LCM" />
                <RESULT eventid="1078" status="DNS" swimtime="00:00:00.00" resultid="1639" heatid="2155" lane="6" entrytime="00:01:03.07" entrycourse="LCM" />
                <RESULT eventid="1106" status="DNS" swimtime="00:00:00.00" resultid="1640" heatid="2192" lane="1" />
                <RESULT eventid="1126" status="DNS" swimtime="00:00:00.00" resultid="1641" heatid="2209" lane="1" entrytime="00:00:56.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Pacheco" birthdate="2012-10-13" gender="F" nation="BRA" license="376981" swrid="5602566" athleteid="1430" externalid="376981">
              <RESULTS>
                <RESULT eventid="1060" points="201" swimtime="00:01:49.44" resultid="1431" heatid="2130" lane="7" entrytime="00:01:59.91" entrycourse="LCM" />
                <RESULT eventid="1084" points="206" swimtime="00:03:10.88" resultid="1432" heatid="2163" lane="4" entrytime="00:03:26.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="187" swimtime="00:03:40.47" resultid="1433" heatid="2183" lane="4" entrytime="00:04:06.77" entrycourse="LCM" />
                <RESULT eventid="1136" points="243" swimtime="00:00:37.82" resultid="1434" heatid="2222" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Emilia Abrahao" birthdate="2016-06-14" gender="F" nation="BRA" license="412012" swrid="5740010" athleteid="1799" externalid="412012">
              <RESULTS>
                <RESULT eventid="1112" status="DNS" swimtime="00:00:00.00" resultid="1800" heatid="2200" lane="6" />
                <RESULT eventid="1132" status="DNS" swimtime="00:00:00.00" resultid="1801" heatid="2220" lane="2" entrytime="00:01:01.96" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Cabrera Cirino Dos Santos" birthdate="2013-03-30" gender="M" nation="BRA" license="376990" swrid="5588570" athleteid="1469" externalid="376990">
              <RESULTS>
                <RESULT eventid="1075" points="169" swimtime="00:00:42.58" resultid="1470" heatid="2152" lane="6" entrytime="00:00:44.03" entrycourse="LCM" />
                <RESULT eventid="1087" points="219" swimtime="00:02:49.15" resultid="1471" heatid="2170" lane="1" entrytime="00:02:55.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="125" swimtime="00:01:38.68" resultid="1472" heatid="2204" lane="5" entrytime="00:01:46.33" entrycourse="LCM" />
                <RESULT eventid="1139" points="210" swimtime="00:00:35.14" resultid="1473" heatid="2232" lane="3" entrytime="00:00:35.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Artigas Pinheiro" birthdate="2013-07-31" gender="F" nation="BRA" license="377153" swrid="5588534" athleteid="1499" externalid="377153">
              <RESULTS>
                <RESULT eventid="1084" points="229" swimtime="00:03:04.34" resultid="1500" heatid="2164" lane="1" entrytime="00:03:15.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="231" swimtime="00:00:43.75" resultid="1501" heatid="2146" lane="4" entrytime="00:00:46.98" entrycourse="LCM" />
                <RESULT eventid="1100" points="192" swimtime="00:03:38.43" resultid="1502" heatid="2184" lane="7" entrytime="00:03:37.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="231" swimtime="00:00:38.47" resultid="1503" heatid="2224" lane="2" entrytime="00:00:40.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Fischer Araujo" birthdate="2013-10-14" gender="M" nation="BRA" license="414420" athleteid="1826" externalid="414420">
              <RESULTS>
                <RESULT eventid="1063" points="66" swimtime="00:02:20.58" resultid="1827" heatid="2133" lane="5" />
                <RESULT eventid="1075" points="58" swimtime="00:01:00.68" resultid="1828" heatid="2149" lane="6" />
                <RESULT eventid="1139" points="66" swimtime="00:00:51.66" resultid="1829" heatid="2229" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Della Villa Yang" birthdate="2012-10-08" gender="F" nation="BRA" license="369276" swrid="5588653" athleteid="1326" externalid="369276">
              <RESULTS>
                <RESULT eventid="1060" points="256" swimtime="00:01:40.88" resultid="1327" heatid="2130" lane="5" entrytime="00:01:43.78" entrycourse="LCM" />
                <RESULT eventid="1084" points="418" swimtime="00:02:30.84" resultid="1328" heatid="2166" lane="3" entrytime="00:02:30.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="341" swimtime="00:03:00.39" resultid="1329" heatid="2185" lane="5" entrytime="00:02:57.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="379" swimtime="00:00:32.61" resultid="1330" heatid="2227" lane="7" entrytime="00:00:32.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Da Cunha Souza" birthdate="2013-09-17" gender="M" nation="BRA" license="376975" swrid="5588618" athleteid="1415" externalid="376975">
              <RESULTS>
                <RESULT eventid="1075" points="156" swimtime="00:00:43.71" resultid="1416" heatid="2150" lane="8" />
                <RESULT eventid="1087" points="180" swimtime="00:03:00.39" resultid="1417" heatid="2169" lane="3" entrytime="00:03:01.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="156" swimtime="00:03:31.53" resultid="1418" heatid="2187" lane="1" />
                <RESULT eventid="1139" points="173" swimtime="00:00:37.51" resultid="1419" heatid="2232" lane="2" entrytime="00:00:35.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Livia Bittencourt" birthdate="2015-11-23" gender="F" nation="BRA" license="393260" swrid="5616446" athleteid="1622" externalid="393260">
              <RESULTS>
                <RESULT eventid="1066" points="78" swimtime="00:01:08.05" resultid="1623" heatid="2137" lane="1" entrytime="00:01:22.77" entrycourse="LCM" />
                <RESULT eventid="1078" points="95" swimtime="00:00:58.67" resultid="1624" heatid="2154" lane="4" entrytime="00:01:11.14" entrycourse="LCM" />
                <RESULT eventid="1106" points="50" swimtime="00:01:06.26" resultid="1625" heatid="2192" lane="2" entrytime="00:01:30.10" entrycourse="LCM" />
                <RESULT eventid="1126" points="74" swimtime="00:00:56.08" resultid="1626" heatid="2208" lane="5" entrytime="00:01:16.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Magalhaes Dabul" birthdate="2014-01-05" gender="M" nation="BRA" license="391023" swrid="5602555" athleteid="1572" externalid="391023">
              <RESULTS>
                <RESULT eventid="1069" points="132" swimtime="00:00:50.96" resultid="1573" heatid="2143" lane="7" entrytime="00:00:51.05" entrycourse="LCM" />
                <RESULT eventid="1093" points="150" swimtime="00:01:28.16" resultid="1574" heatid="2179" lane="8" entrytime="00:01:37.53" entrycourse="LCM" />
                <RESULT eventid="1129" points="158" swimtime="00:00:38.67" resultid="1575" heatid="2215" lane="6" entrytime="00:00:47.51" entrycourse="LCM" />
                <RESULT eventid="1109" points="147" swimtime="00:00:42.17" resultid="1576" heatid="2199" lane="6" entrytime="00:00:43.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="De Fortes" birthdate="2015-06-01" gender="M" nation="BRA" license="399680" swrid="5652884" athleteid="1677" externalid="399680">
              <RESULTS>
                <RESULT eventid="1081" points="102" swimtime="00:00:50.38" resultid="1678" heatid="2160" lane="1" entrytime="00:00:52.95" entrycourse="LCM" />
                <RESULT eventid="1093" points="133" swimtime="00:01:31.62" resultid="1679" heatid="2177" lane="6" />
                <RESULT eventid="1129" points="129" swimtime="00:00:41.32" resultid="1680" heatid="2214" lane="8" />
                <RESULT eventid="1109" points="104" swimtime="00:00:47.21" resultid="1681" heatid="2198" lane="5" entrytime="00:00:50.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Brandt Macedo" birthdate="2013-04-19" gender="M" nation="BRA" license="414421" athleteid="1830" externalid="414421">
              <RESULTS>
                <RESULT comment="SW 6.2 - Deixou a posição de costas, exceto ao executar uma virada.  (Horário: 10:17), Antes da chegada." eventid="1075" status="DSQ" swimtime="00:01:02.67" resultid="1831" heatid="2150" lane="2" />
                <RESULT eventid="1139" points="60" swimtime="00:00:53.17" resultid="1832" heatid="2229" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Stramandinoli Zanicotti" birthdate="2013-06-18" gender="F" nation="BRA" license="376967" swrid="5588924" athleteid="1395" externalid="376967">
              <RESULTS>
                <RESULT eventid="1060" points="142" swimtime="00:02:02.65" resultid="1396" heatid="2130" lane="1" entrytime="00:02:06.36" entrycourse="LCM" />
                <RESULT eventid="1072" points="142" swimtime="00:00:51.46" resultid="1397" heatid="2146" lane="7" entrytime="00:00:50.37" entrycourse="LCM" />
                <RESULT eventid="1100" points="136" swimtime="00:04:05.23" resultid="1398" heatid="2183" lane="3" entrytime="00:04:11.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:03.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="181" swimtime="00:00:41.73" resultid="1399" heatid="2223" lane="7" entrytime="00:00:43.05" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gael" lastname="Stramandinoli Zanicotti" birthdate="2015-03-21" gender="M" nation="BRA" license="406954" swrid="5717298" athleteid="1758" externalid="406954">
              <RESULTS>
                <RESULT eventid="1081" points="56" swimtime="00:01:01.23" resultid="1759" heatid="2158" lane="5" entrytime="00:01:05.59" entrycourse="LCM" />
                <RESULT eventid="1093" points="51" swimtime="00:02:06.18" resultid="1760" heatid="2177" lane="3" entrytime="00:02:16.58" entrycourse="LCM" />
                <RESULT eventid="1129" points="50" swimtime="00:00:56.59" resultid="1761" heatid="2214" lane="3" entrytime="00:01:00.21" entrycourse="LCM" />
                <RESULT eventid="1109" points="17" swimtime="00:01:25.97" resultid="1762" heatid="2195" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Dolberth Alcantara" birthdate="2014-09-26" gender="F" nation="BRA" license="382124" swrid="5602532" athleteid="1509" externalid="382124">
              <RESULTS>
                <RESULT eventid="1078" points="168" swimtime="00:00:48.62" resultid="1510" heatid="2156" lane="3" entrytime="00:00:51.88" entrycourse="LCM" />
                <RESULT eventid="1090" points="157" swimtime="00:01:35.76" resultid="1511" heatid="2173" lane="3" entrytime="00:02:02.77" entrycourse="LCM" />
                <RESULT eventid="1106" points="142" swimtime="00:00:46.74" resultid="1512" heatid="2193" lane="4" entrytime="00:00:51.41" entrycourse="LCM" />
                <RESULT eventid="1126" points="168" swimtime="00:00:42.72" resultid="1513" heatid="2209" lane="5" entrytime="00:00:52.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Szpak De Vasconcelos" birthdate="2012-06-29" gender="M" nation="BRA" license="369271" swrid="5588928" athleteid="1311" externalid="369271">
              <RESULTS>
                <RESULT eventid="1063" points="300" swimtime="00:01:24.96" resultid="1312" heatid="2135" lane="4" entrytime="00:01:26.59" entrycourse="LCM" />
                <RESULT eventid="1087" points="313" swimtime="00:02:30.10" resultid="1313" heatid="2171" lane="4" entrytime="00:02:30.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="297" swimtime="00:02:50.83" resultid="1314" heatid="2189" lane="4" entrytime="00:02:56.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="331" swimtime="00:00:30.22" resultid="1315" heatid="2234" lane="4" entrytime="00:00:30.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Coelho Ghignone" birthdate="2015-01-05" gender="M" nation="BRA" license="410201" swrid="5740006" athleteid="1786" externalid="410201">
              <RESULTS>
                <RESULT eventid="1081" points="128" swimtime="00:00:46.72" resultid="1787" heatid="2161" lane="8" entrytime="00:00:48.24" entrycourse="LCM" />
                <RESULT eventid="1093" points="117" swimtime="00:01:35.57" resultid="1788" heatid="2178" lane="2" entrytime="00:01:44.70" entrycourse="LCM" />
                <RESULT eventid="1129" points="109" swimtime="00:00:43.72" resultid="1789" heatid="2216" lane="8" entrytime="00:00:44.92" entrycourse="LCM" />
                <RESULT eventid="1109" points="61" swimtime="00:00:56.47" resultid="1790" heatid="2196" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Toscani Kim" birthdate="2013-02-15" gender="F" nation="BRA" license="372683" swrid="5588939" athleteid="1366" externalid="372683">
              <RESULTS>
                <RESULT eventid="1060" points="312" swimtime="00:01:34.51" resultid="1367" heatid="2131" lane="6" entrytime="00:01:36.12" entrycourse="LCM" />
                <RESULT eventid="1084" points="319" swimtime="00:02:45.01" resultid="1368" heatid="2165" lane="8" entrytime="00:02:57.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="310" swimtime="00:03:06.24" resultid="1369" heatid="2185" lane="8" entrytime="00:03:10.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="311" swimtime="00:00:34.84" resultid="1370" heatid="2225" lane="3" entrytime="00:00:36.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Cipriani Presiazniuk" birthdate="2012-07-03" gender="M" nation="BRA" license="369267" swrid="5588594" athleteid="1296" externalid="369267">
              <RESULTS>
                <RESULT eventid="1075" points="211" swimtime="00:00:39.50" resultid="1297" heatid="2153" lane="1" entrytime="00:00:39.75" entrycourse="LCM" />
                <RESULT eventid="1087" points="254" swimtime="00:02:40.90" resultid="1298" heatid="2170" lane="7" entrytime="00:02:53.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="205" swimtime="00:03:13.15" resultid="1299" heatid="2188" lane="5" entrytime="00:03:23.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="259" swimtime="00:00:32.79" resultid="1300" heatid="2232" lane="7" entrytime="00:00:35.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joana" lastname="Asinelli Casagrande" birthdate="2013-10-26" gender="F" nation="BRA" license="376970" swrid="5588536" athleteid="1405" externalid="376970">
              <RESULTS>
                <RESULT eventid="1060" points="200" swimtime="00:01:49.55" resultid="1406" heatid="2130" lane="8" />
                <RESULT eventid="1072" points="264" swimtime="00:00:41.82" resultid="1407" heatid="2147" lane="2" entrytime="00:00:44.67" entrycourse="LCM" />
                <RESULT eventid="1100" points="276" swimtime="00:03:13.61" resultid="1408" heatid="2184" lane="3" entrytime="00:03:14.43" entrycourse="LCM" />
                <RESULT eventid="1116" points="198" swimtime="00:01:35.16" resultid="1409" heatid="2203" lane="6" entrytime="00:01:33.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Gois Nogueira" birthdate="2014-03-11" gender="F" nation="BRA" license="393258" swrid="5616443" athleteid="1612" externalid="393258">
              <RESULTS>
                <RESULT eventid="1066" points="164" swimtime="00:00:53.22" resultid="1613" heatid="2138" lane="4" entrytime="00:00:56.26" entrycourse="LCM" />
                <RESULT eventid="1078" points="146" swimtime="00:00:50.99" resultid="1614" heatid="2156" lane="5" entrytime="00:00:51.82" entrycourse="LCM" />
                <RESULT eventid="1106" points="78" swimtime="00:00:56.96" resultid="1615" heatid="2193" lane="1" entrytime="00:00:57.36" entrycourse="LCM" />
                <RESULT eventid="1126" points="176" swimtime="00:00:42.10" resultid="1616" heatid="2211" lane="5" entrytime="00:00:42.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Lauand Lorenci" birthdate="2013-03-06" gender="M" nation="BRA" license="376982" swrid="5588764" athleteid="1435" externalid="376982">
              <RESULTS>
                <RESULT eventid="1063" points="206" swimtime="00:01:36.16" resultid="1436" heatid="2133" lane="8" />
                <RESULT eventid="1087" points="183" swimtime="00:02:59.63" resultid="1437" heatid="2167" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="209" swimtime="00:03:11.99" resultid="1438" heatid="2189" lane="6" entrytime="00:03:10.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="228" swimtime="00:00:34.22" resultid="1439" heatid="2233" lane="1" entrytime="00:00:34.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cecilia Carvalho" birthdate="2014-10-30" gender="F" nation="BRA" license="391021" swrid="5602525" athleteid="1567" externalid="391021">
              <RESULTS>
                <RESULT eventid="1078" points="151" swimtime="00:00:50.41" resultid="1568" heatid="2155" lane="4" entrytime="00:01:00.22" entrycourse="LCM" />
                <RESULT eventid="1090" points="140" swimtime="00:01:39.53" resultid="1569" heatid="2173" lane="6" entrytime="00:02:05.11" entrycourse="LCM" />
                <RESULT eventid="1106" points="77" swimtime="00:00:57.32" resultid="1570" heatid="2191" lane="1" />
                <RESULT eventid="1126" points="152" swimtime="00:00:44.16" resultid="1571" heatid="2209" lane="3" entrytime="00:00:52.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Caron Braga" birthdate="2016-02-01" gender="F" nation="BRA" license="415256" athleteid="1851" externalid="415256">
              <RESULTS>
                <RESULT eventid="1122" points="66" swimtime="00:01:11.99" resultid="1852" heatid="2206" lane="2" />
                <RESULT eventid="1132" points="41" swimtime="00:01:08.36" resultid="1853" heatid="2219" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Weber Boguszewski" birthdate="2016-10-07" gender="M" nation="BRA" license="415255" athleteid="1848" externalid="415255">
              <RESULTS>
                <RESULT eventid="1114" points="52" swimtime="00:01:03.08" resultid="1849" heatid="2201" lane="3" />
                <RESULT eventid="1134" points="25" swimtime="00:01:10.83" resultid="1850" heatid="2221" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Petraglia" birthdate="2012-03-28" gender="M" nation="BRA" license="369282" swrid="5602569" athleteid="1351" externalid="369282">
              <RESULTS>
                <RESULT eventid="1063" points="184" swimtime="00:01:39.98" resultid="1352" heatid="2135" lane="2" entrytime="00:01:39.37" entrycourse="LCM" />
                <RESULT eventid="1075" points="199" swimtime="00:00:40.33" resultid="1353" heatid="2153" lane="2" entrytime="00:00:38.88" entrycourse="LCM" />
                <RESULT eventid="1103" points="197" swimtime="00:03:15.85" resultid="1354" heatid="2187" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="259" swimtime="00:00:32.80" resultid="1355" heatid="2228" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Jarenko Gomes" birthdate="2014-05-17" gender="F" nation="BRA" license="407692" swrid="5725992" athleteid="1776" externalid="407692">
              <RESULTS>
                <RESULT eventid="1066" points="105" swimtime="00:01:01.64" resultid="1777" heatid="2136" lane="4" />
                <RESULT eventid="1078" points="99" swimtime="00:00:57.92" resultid="1778" heatid="2154" lane="3" />
                <RESULT eventid="1106" points="45" swimtime="00:01:08.23" resultid="1779" heatid="2192" lane="8" />
                <RESULT eventid="1126" points="98" swimtime="00:00:51.11" resultid="1780" heatid="2209" lane="6" entrytime="00:00:53.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alan" lastname="Batista Grise" birthdate="2014-03-27" gender="M" nation="BRA" license="391007" swrid="5602513" athleteid="1534" externalid="391007">
              <RESULTS>
                <RESULT eventid="1069" status="DNS" swimtime="00:00:00.00" resultid="1535" heatid="2141" lane="4" entrytime="00:01:00.33" entrycourse="LCM" />
                <RESULT eventid="1081" status="DNS" swimtime="00:00:00.00" resultid="1536" heatid="2159" lane="5" entrytime="00:00:56.30" entrycourse="LCM" />
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="1537" heatid="2215" lane="2" entrytime="00:00:48.74" entrycourse="LCM" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="1538" heatid="2196" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Wolf Macedo" birthdate="2012-01-27" gender="F" nation="BRA" license="369277" swrid="5602592" athleteid="1331" externalid="369277">
              <RESULTS>
                <RESULT eventid="1084" points="372" swimtime="00:02:36.80" resultid="1332" heatid="2166" lane="7" entrytime="00:02:36.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="317" swimtime="00:00:39.38" resultid="1333" heatid="2145" lane="8" />
                <RESULT eventid="1116" points="247" swimtime="00:01:28.33" resultid="1334" heatid="2203" lane="5" entrytime="00:01:23.68" entrycourse="LCM" />
                <RESULT eventid="1136" points="389" swimtime="00:00:32.34" resultid="1335" heatid="2222" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Azevedo Alanis" birthdate="2013-12-07" gender="M" nation="BRA" license="376991" swrid="5588540" athleteid="1464" externalid="376991">
              <RESULTS>
                <RESULT eventid="1063" points="164" swimtime="00:01:43.87" resultid="1465" heatid="2135" lane="8" entrytime="00:01:49.20" entrycourse="LCM" />
                <RESULT eventid="1087" points="162" swimtime="00:03:07.05" resultid="1466" heatid="2167" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="179" swimtime="00:03:22.14" resultid="1467" heatid="2188" lane="6" entrytime="00:03:35.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="155" swimtime="00:00:38.90" resultid="1468" heatid="2230" lane="3" entrytime="00:00:42.22" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Tallao Benke" birthdate="2012-01-02" gender="F" nation="BRA" license="376984" swrid="5588931" athleteid="1445" externalid="376984">
              <RESULTS>
                <RESULT eventid="1084" points="476" swimtime="00:02:24.48" resultid="1446" heatid="2166" lane="4" entrytime="00:02:25.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="456" swimtime="00:00:34.88" resultid="1447" heatid="2148" lane="5" entrytime="00:00:35.31" entrycourse="LCM" />
                <RESULT eventid="1116" points="416" swimtime="00:01:14.29" resultid="1448" heatid="2203" lane="4" entrytime="00:01:14.85" entrycourse="LCM" />
                <RESULT eventid="1136" points="505" swimtime="00:00:29.64" resultid="1449" heatid="2227" lane="5" entrytime="00:00:30.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Wolff Contin" birthdate="2015-10-10" gender="M" nation="BRA" license="406745" swrid="5717303" athleteid="1722" externalid="406745">
              <RESULTS>
                <RESULT eventid="1081" points="63" swimtime="00:00:59.13" resultid="1723" heatid="2159" lane="8" entrytime="00:01:04.76" entrycourse="LCM" />
                <RESULT eventid="1093" points="59" swimtime="00:02:00.28" resultid="1724" heatid="2177" lane="4" entrytime="00:02:00.58" entrycourse="LCM" />
                <RESULT eventid="1129" points="62" swimtime="00:00:52.77" resultid="1725" heatid="2215" lane="1" entrytime="00:00:50.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Corte Flor" birthdate="2016-12-03" gender="M" nation="BRA" license="412013" swrid="5740007" athleteid="1802" externalid="412013">
              <RESULTS>
                <RESULT eventid="1124" points="50" swimtime="00:01:10.17" resultid="1803" heatid="2207" lane="3" />
                <RESULT eventid="1134" status="DNS" swimtime="00:00:00.00" resultid="1804" heatid="2221" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Saber" birthdate="2014-06-04" gender="F" nation="BRA" license="392141" swrid="5602554" athleteid="1607" externalid="392141">
              <RESULTS>
                <RESULT eventid="1066" points="206" swimtime="00:00:49.34" resultid="1608" heatid="2139" lane="3" entrytime="00:00:51.88" entrycourse="LCM" />
                <RESULT eventid="1078" points="165" swimtime="00:00:48.94" resultid="1609" heatid="2156" lane="6" entrytime="00:00:52.79" entrycourse="LCM" />
                <RESULT eventid="1106" points="99" swimtime="00:00:52.71" resultid="1610" heatid="2192" lane="6" entrytime="00:01:11.88" entrycourse="LCM" />
                <RESULT eventid="1126" points="176" swimtime="00:00:42.10" resultid="1611" heatid="2208" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luigi" lastname="Antoniuk Paganini" birthdate="2014-11-13" gender="M" nation="BRA" license="382127" swrid="5602509" athleteid="1519" externalid="382127">
              <RESULTS>
                <RESULT eventid="1081" points="190" swimtime="00:00:40.90" resultid="1520" heatid="2160" lane="3" entrytime="00:00:50.05" entrycourse="LCM" />
                <RESULT eventid="1093" points="209" swimtime="00:01:18.92" resultid="1521" heatid="2180" lane="8" entrytime="00:01:29.15" entrycourse="LCM" />
                <RESULT eventid="1129" points="183" swimtime="00:00:36.82" resultid="1522" heatid="2216" lane="1" entrytime="00:00:44.80" entrycourse="LCM" />
                <RESULT eventid="1109" points="144" swimtime="00:00:42.45" resultid="1523" heatid="2198" lane="8" entrytime="00:00:59.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Lazzarotti Matias" birthdate="2012-03-19" gender="F" nation="BRA" license="391026" swrid="5602552" athleteid="1587" externalid="391026">
              <RESULTS>
                <RESULT eventid="1084" points="375" swimtime="00:02:36.41" resultid="1588" heatid="2162" lane="6" />
                <RESULT eventid="1072" points="423" swimtime="00:00:35.78" resultid="1589" heatid="2148" lane="3" entrytime="00:00:35.63" entrycourse="LCM" />
                <RESULT eventid="1100" points="318" swimtime="00:03:04.64" resultid="1590" heatid="2184" lane="4" entrytime="00:03:11.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="394" swimtime="00:00:32.19" resultid="1591" heatid="2227" lane="2" entrytime="00:00:31.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elisa" lastname="Osternack Almeida" birthdate="2015-04-14" gender="F" nation="BRA" license="406747" swrid="5717286" athleteid="1726" externalid="406747" />
            <ATHLETE firstname="Miguel" lastname="Fernandes  Dos Reis" birthdate="2012-09-18" gender="M" nation="BRA" license="369279" swrid="5588696" athleteid="1341" externalid="369279">
              <RESULTS>
                <RESULT eventid="1063" points="156" swimtime="00:01:45.48" resultid="1342" heatid="2134" lane="8" />
                <RESULT eventid="1087" points="250" swimtime="00:02:41.78" resultid="1343" heatid="2171" lane="6" entrytime="00:02:36.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="161" swimtime="00:01:30.76" resultid="1344" heatid="2205" lane="5" entrytime="00:01:19.97" entrycourse="LCM" />
                <RESULT eventid="1139" points="241" swimtime="00:00:33.57" resultid="1345" heatid="2234" lane="1" entrytime="00:00:32.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Miranda Carvalho" birthdate="2015-07-07" gender="F" nation="BRA" license="410200" swrid="5740015" athleteid="1781" externalid="410200">
              <RESULTS>
                <RESULT eventid="1066" points="72" swimtime="00:01:10.05" resultid="1782" heatid="2137" lane="3" entrytime="00:01:09.01" entrycourse="LCM" />
                <RESULT eventid="1078" points="79" swimtime="00:01:02.39" resultid="1783" heatid="2155" lane="1" entrytime="00:01:04.00" entrycourse="LCM" />
                <RESULT eventid="1106" points="41" swimtime="00:01:10.83" resultid="1784" heatid="2191" lane="5" />
                <RESULT eventid="1126" points="58" swimtime="00:01:00.77" resultid="1785" heatid="2209" lane="2" entrytime="00:00:56.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Karam Barbosa Lima" birthdate="2012-12-11" gender="F" nation="BRA" license="376956" swrid="5588758" athleteid="1371" externalid="376956">
              <RESULTS>
                <RESULT eventid="1060" points="217" swimtime="00:01:46.60" resultid="1372" heatid="2129" lane="3" />
                <RESULT eventid="1072" points="335" swimtime="00:00:38.67" resultid="1373" heatid="2148" lane="2" entrytime="00:00:38.73" entrycourse="LCM" />
                <RESULT eventid="1100" points="285" swimtime="00:03:11.51" resultid="1374" heatid="2183" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="364" swimtime="00:00:33.04" resultid="1375" heatid="2226" lane="2" entrytime="00:00:33.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Calvo Ribas" birthdate="2016-01-09" gender="M" nation="BRA" license="415014" athleteid="1845" externalid="415014">
              <RESULTS>
                <RESULT eventid="1114" points="77" swimtime="00:00:55.21" resultid="1846" heatid="2201" lane="6" />
                <RESULT eventid="1134" points="33" swimtime="00:01:05.06" resultid="1847" heatid="2221" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcela" lastname="Tallao Benke" birthdate="2014-10-07" gender="F" nation="BRA" license="382075" swrid="5602586" athleteid="1504" externalid="382075">
              <RESULTS>
                <RESULT eventid="1066" points="228" swimtime="00:00:47.67" resultid="1505" heatid="2139" lane="5" entrytime="00:00:48.43" entrycourse="LCM" />
                <RESULT eventid="1090" points="321" swimtime="00:01:15.48" resultid="1506" heatid="2175" lane="5" entrytime="00:01:26.53" entrycourse="LCM" />
                <RESULT eventid="1106" points="228" swimtime="00:00:39.97" resultid="1507" heatid="2194" lane="4" entrytime="00:00:41.31" entrycourse="LCM" />
                <RESULT eventid="1126" points="310" swimtime="00:00:34.88" resultid="1508" heatid="2212" lane="5" entrytime="00:00:36.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2864" nation="BRA" region="PR" clubid="1144" swrid="93756" name="Associacao De Pais E Amigos Da Natacao De Ponta Gr" shortname="Apan Ponta Grossa">
          <ATHLETES>
            <ATHLETE firstname="Gustavo" lastname="Hilgenberg Lievore" birthdate="2014-04-23" gender="M" nation="BRA" license="391167" swrid="5602546" athleteid="1164" externalid="391167">
              <RESULTS>
                <RESULT eventid="1129" points="180" swimtime="00:00:36.99" resultid="1165" heatid="2218" lane="2" entrytime="00:00:36.84" entrycourse="LCM" />
                <RESULT eventid="1109" points="140" swimtime="00:00:42.86" resultid="1166" heatid="2199" lane="7" entrytime="00:00:47.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariana" lastname="Brunetti Silva" birthdate="2014-03-24" gender="F" nation="BRA" license="390878" swrid="5602517" athleteid="1159" externalid="390878">
              <RESULTS>
                <RESULT eventid="1066" points="148" swimtime="00:00:55.06" resultid="1160" heatid="2139" lane="8" entrytime="00:00:54.91" entrycourse="LCM" />
                <RESULT eventid="1078" points="133" swimtime="00:00:52.58" resultid="1161" heatid="2157" lane="1" entrytime="00:00:50.19" entrycourse="LCM" />
                <RESULT eventid="1106" points="84" swimtime="00:00:55.64" resultid="1162" heatid="2193" lane="5" entrytime="00:00:53.21" entrycourse="LCM" />
                <RESULT eventid="1126" points="187" swimtime="00:00:41.24" resultid="1163" heatid="2212" lane="2" entrytime="00:00:40.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Clara Domingues" birthdate="2012-01-19" gender="F" nation="BRA" license="377291" swrid="5588599" athleteid="1145" externalid="377291">
              <RESULTS>
                <RESULT eventid="1084" points="296" swimtime="00:02:49.15" resultid="1146" heatid="2164" lane="6" entrytime="00:03:06.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="231" swimtime="00:00:43.76" resultid="1147" heatid="2145" lane="4" entrytime="00:00:51.97" entrycourse="LCM" />
                <RESULT eventid="1136" points="279" swimtime="00:00:36.11" resultid="1148" heatid="2224" lane="8" entrytime="00:00:42.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Campagnoli" birthdate="2013-03-13" gender="M" nation="BRA" license="370651" swrid="5602519" athleteid="1149" externalid="370651">
              <RESULTS>
                <RESULT eventid="1075" points="280" swimtime="00:00:35.97" resultid="1150" heatid="2153" lane="3" entrytime="00:00:37.08" entrycourse="LCM" />
                <RESULT eventid="1087" points="241" swimtime="00:02:43.79" resultid="1151" heatid="2171" lane="8" entrytime="00:02:40.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="205" swimtime="00:01:23.86" resultid="1152" heatid="2205" lane="3" entrytime="00:01:21.92" entrycourse="LCM" />
                <RESULT eventid="1139" points="264" swimtime="00:00:32.58" resultid="1153" heatid="2234" lane="2" entrytime="00:00:31.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Miretzki" birthdate="2014-09-17" gender="F" nation="BRA" license="414996" athleteid="1179" externalid="414996">
              <RESULTS>
                <RESULT eventid="1066" points="115" swimtime="00:00:59.88" resultid="1180" heatid="2136" lane="3" />
                <RESULT eventid="1090" points="170" swimtime="00:01:33.18" resultid="1181" heatid="2172" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolly" lastname="Victoria Souza" birthdate="2015-11-15" gender="F" nation="BRA" license="400091" swrid="5652902" athleteid="1170" externalid="400091">
              <RESULTS>
                <RESULT eventid="1066" points="153" swimtime="00:00:54.46" resultid="1171" heatid="2138" lane="5" entrytime="00:00:57.94" entrycourse="LCM" />
                <RESULT eventid="1090" points="128" swimtime="00:01:42.52" resultid="1172" heatid="2174" lane="8" entrytime="00:01:51.62" entrycourse="LCM" />
                <RESULT eventid="1126" points="175" swimtime="00:00:42.17" resultid="1173" heatid="2210" lane="3" entrytime="00:00:45.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Bischof Rogoski" birthdate="2014-10-03" gender="M" nation="BRA" license="401860" swrid="5661341" athleteid="1174" externalid="401860">
              <RESULTS>
                <RESULT eventid="1069" points="137" swimtime="00:00:50.23" resultid="1175" heatid="2142" lane="3" entrytime="00:00:55.28" entrycourse="LCM" />
                <RESULT eventid="1093" points="189" swimtime="00:01:21.64" resultid="1176" heatid="2180" lane="1" entrytime="00:01:28.73" entrycourse="LCM" />
                <RESULT eventid="1129" points="189" swimtime="00:00:36.39" resultid="1177" heatid="2218" lane="7" entrytime="00:00:36.97" entrycourse="LCM" />
                <RESULT eventid="1109" points="140" swimtime="00:00:42.79" resultid="1178" heatid="2196" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Clara Rigailo" birthdate="2013-04-06" gender="F" nation="BRA" license="396828" swrid="5641758" athleteid="1167" externalid="396828">
              <RESULTS>
                <RESULT eventid="1060" points="300" swimtime="00:01:35.73" resultid="1168" heatid="2131" lane="2" entrytime="00:01:36.33" entrycourse="LCM" />
                <RESULT eventid="1072" points="202" swimtime="00:00:45.73" resultid="1169" heatid="2147" lane="8" entrytime="00:00:46.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emanuel" lastname="Lucas Ribeiro" birthdate="2014-03-28" gender="M" nation="BRA" license="414997" athleteid="1182" externalid="414997">
              <RESULTS>
                <RESULT eventid="1069" points="99" swimtime="00:00:56.03" resultid="1183" heatid="2140" lane="3" />
                <RESULT eventid="1081" points="76" swimtime="00:00:55.42" resultid="1184" heatid="2158" lane="2" />
                <RESULT eventid="1129" points="96" swimtime="00:00:45.56" resultid="1185" heatid="2213" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Victoria Borges" birthdate="2014-01-16" gender="F" nation="BRA" license="376737" swrid="5602587" athleteid="1154" externalid="376737">
              <RESULTS>
                <RESULT eventid="1078" points="194" swimtime="00:00:46.32" resultid="1155" heatid="2157" lane="7" entrytime="00:00:48.84" entrycourse="LCM" />
                <RESULT eventid="1090" points="186" swimtime="00:01:30.58" resultid="1156" heatid="2175" lane="1" entrytime="00:01:34.92" entrycourse="LCM" />
                <RESULT eventid="1106" points="100" swimtime="00:00:52.55" resultid="1157" heatid="2191" lane="8" />
                <RESULT eventid="1126" points="245" swimtime="00:00:37.71" resultid="1158" heatid="2212" lane="6" entrytime="00:00:40.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13068" nation="BRA" region="PR" clubid="1919" swrid="93787" name="Sociedade Morgenau" shortname="Morgenau">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Fernanda De Lima" birthdate="2013-09-26" gender="F" nation="BRA" license="378290" swrid="5588693" athleteid="1925" externalid="378290">
              <RESULTS>
                <RESULT eventid="1084" points="184" swimtime="00:03:18.13" resultid="1926" heatid="2163" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="247" swimtime="00:00:42.78" resultid="1927" heatid="2146" lane="5" entrytime="00:00:47.12" entrycourse="LCM" />
                <RESULT eventid="1136" points="212" swimtime="00:00:39.56" resultid="1928" heatid="2223" lane="1" entrytime="00:00:43.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Nitz Costa" birthdate="2015-02-09" gender="F" nation="BRA" license="397328" swrid="5641773" athleteid="1939" externalid="397328">
              <RESULTS>
                <RESULT eventid="1066" points="180" swimtime="00:00:51.56" resultid="1940" heatid="2137" lane="4" entrytime="00:01:06.57" entrycourse="LCM" />
                <RESULT eventid="1090" points="252" swimtime="00:01:21.86" resultid="1941" heatid="2175" lane="7" entrytime="00:01:32.45" entrycourse="LCM" />
                <RESULT eventid="1106" points="182" swimtime="00:00:43.07" resultid="1942" heatid="2194" lane="3" entrytime="00:00:47.00" entrycourse="LCM" />
                <RESULT eventid="1126" points="244" swimtime="00:00:37.75" resultid="1943" heatid="2212" lane="7" entrytime="00:00:40.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Paes Pereira" birthdate="2013-03-11" gender="M" nation="BRA" license="391137" swrid="5602567" athleteid="1929" externalid="391137">
              <RESULTS>
                <RESULT eventid="1075" points="114" swimtime="00:00:48.43" resultid="1930" heatid="2151" lane="8" entrytime="00:00:51.05" entrycourse="LCM" />
                <RESULT eventid="1087" points="120" swimtime="00:03:26.56" resultid="1931" heatid="2168" lane="3" entrytime="00:03:46.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="95" swimtime="00:04:09.38" resultid="1932" heatid="2187" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:56.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="128" swimtime="00:00:41.45" resultid="1933" heatid="2230" lane="2" entrytime="00:00:43.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cecilia Carstens" birthdate="2014-02-22" gender="F" nation="BRA" license="406721" swrid="5717251" athleteid="1954" externalid="406721">
              <RESULTS>
                <RESULT eventid="1090" points="149" swimtime="00:01:37.42" resultid="1955" heatid="2174" lane="2" entrytime="00:01:46.50" entrycourse="LCM" />
                <RESULT eventid="1106" points="121" swimtime="00:00:49.35" resultid="1956" heatid="2193" lane="7" entrytime="00:00:56.35" entrycourse="LCM" />
                <RESULT eventid="1126" points="165" swimtime="00:00:42.96" resultid="1957" heatid="2208" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Tomaz Zmievski" birthdate="2012-09-20" gender="F" nation="BRA" license="406725" swrid="5717300" athleteid="1958" externalid="406725">
              <RESULTS>
                <RESULT eventid="1084" points="227" swimtime="00:03:04.99" resultid="1959" heatid="2164" lane="8" entrytime="00:03:22.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="201" swimtime="00:03:35.15" resultid="1960" heatid="2182" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:46.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="278" swimtime="00:00:36.17" resultid="1961" heatid="2222" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Lara" birthdate="2014-09-02" gender="F" nation="BRA" license="406686" swrid="5717259" athleteid="1944" externalid="406686">
              <RESULTS>
                <RESULT eventid="1066" points="98" swimtime="00:01:03.13" resultid="1945" heatid="2136" lane="5" />
                <RESULT eventid="1090" points="184" swimtime="00:01:30.77" resultid="1946" heatid="2172" lane="6" />
                <RESULT eventid="1106" points="94" swimtime="00:00:53.72" resultid="1947" heatid="2191" lane="2" />
                <RESULT eventid="1126" points="199" swimtime="00:00:40.41" resultid="1948" heatid="2211" lane="8" entrytime="00:00:44.24" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Felipe Kuhn" birthdate="2014-03-22" gender="M" nation="BRA" license="392121" swrid="5602536" athleteid="1934" externalid="392121">
              <RESULTS>
                <RESULT eventid="1069" points="131" swimtime="00:00:51.00" resultid="1935" heatid="2143" lane="6" entrytime="00:00:50.20" entrycourse="LCM" />
                <RESULT eventid="1093" points="143" swimtime="00:01:29.47" resultid="1936" heatid="2176" lane="5" />
                <RESULT eventid="1129" points="172" swimtime="00:00:37.56" resultid="1937" heatid="2217" lane="2" entrytime="00:00:39.93" entrycourse="LCM" />
                <RESULT eventid="1109" status="DNS" swimtime="00:00:00.00" resultid="1938" heatid="2195" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Seiffert Mafra" birthdate="2013-01-11" gender="F" nation="BRA" license="406729" swrid="5717296" athleteid="1962" externalid="406729">
              <RESULTS>
                <RESULT comment="SW 8.5 - Totalmente submerso durante o nado.  (Horário: 15:48)" eventid="1100" status="DSQ" swimtime="00:04:03.51" resultid="1963" heatid="2182" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:58.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="158" swimtime="00:00:43.64" resultid="1964" heatid="2222" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Alves" birthdate="2012-10-12" gender="M" nation="BRA" license="369324" swrid="5588674" athleteid="1920" externalid="369324">
              <RESULTS>
                <RESULT eventid="1075" points="283" swimtime="00:00:35.83" resultid="1921" heatid="2153" lane="4" entrytime="00:00:35.95" entrycourse="LCM" />
                <RESULT eventid="1087" points="255" swimtime="00:02:40.64" resultid="1922" heatid="2169" lane="6" entrytime="00:03:02.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="233" swimtime="00:03:05.09" resultid="1923" heatid="2189" lane="2" entrytime="00:03:11.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.90" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 8.5 - Totalmente submerso durante o nado.  (Horário: 17:03)" eventid="1119" status="DSQ" swimtime="00:01:40.24" resultid="1924" heatid="2204" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Melo" birthdate="2015-02-07" gender="F" nation="BRA" license="406717" swrid="5717280" athleteid="1949" externalid="406717">
              <RESULTS>
                <RESULT eventid="1078" points="227" swimtime="00:00:43.99" resultid="1950" heatid="2157" lane="2" entrytime="00:00:48.72" entrycourse="LCM" />
                <RESULT eventid="1090" points="165" swimtime="00:01:34.14" resultid="1951" heatid="2172" lane="1" />
                <RESULT eventid="1106" points="106" swimtime="00:00:51.46" resultid="1952" heatid="2194" lane="7" entrytime="00:00:50.43" entrycourse="LCM" />
                <RESULT eventid="1126" points="158" swimtime="00:00:43.66" resultid="1953" heatid="2210" lane="4" entrytime="00:00:44.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1007" nation="BRA" region="PR" clubid="1965" swrid="93785" name="Santa Mônica Clube De Campo" shortname="Santa Mônica">
          <ATHLETES>
            <ATHLETE firstname="Cleverson" lastname="Cardoso" birthdate="2013-07-20" gender="M" nation="BRA" license="387382" swrid="5588577" athleteid="2028" externalid="387382">
              <RESULTS>
                <RESULT eventid="1063" points="157" swimtime="00:01:45.34" resultid="2029" heatid="2133" lane="3" />
                <RESULT eventid="1075" points="124" swimtime="00:00:47.22" resultid="2030" heatid="2151" lane="7" entrytime="00:00:48.90" entrycourse="LCM" />
                <RESULT eventid="1139" points="190" swimtime="00:00:36.34" resultid="2031" heatid="2231" lane="8" entrytime="00:00:39.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="Cirilo Da Cunha" birthdate="2013-05-26" gender="F" nation="BRA" license="377316" swrid="5588595" athleteid="1981" externalid="377316">
              <RESULTS>
                <RESULT eventid="1084" points="295" swimtime="00:02:49.34" resultid="1982" heatid="2165" lane="5" entrytime="00:02:49.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="253" swimtime="00:00:42.46" resultid="1983" heatid="2147" lane="1" entrytime="00:00:45.94" entrycourse="LCM" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 15:58), Virada dos 150M." eventid="1100" status="DSQ" swimtime="00:03:23.28" resultid="1984" heatid="2184" lane="2" entrytime="00:03:29.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="249" swimtime="00:00:37.51" resultid="1985" heatid="2225" lane="1" entrytime="00:00:37.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Vieira Coelho" birthdate="2014-09-28" gender="F" nation="BRA" license="406951" swrid="5717301" athleteid="2105" externalid="406951">
              <RESULTS>
                <RESULT eventid="1066" points="175" swimtime="00:00:52.06" resultid="2106" heatid="2139" lane="1" entrytime="00:00:53.92" entrycourse="LCM" />
                <RESULT eventid="1090" points="208" swimtime="00:01:27.24" resultid="2107" heatid="2175" lane="2" entrytime="00:01:31.81" entrycourse="LCM" />
                <RESULT eventid="1106" points="115" swimtime="00:00:50.21" resultid="2108" heatid="2193" lane="3" entrytime="00:00:53.23" entrycourse="LCM" />
                <RESULT eventid="1126" points="227" swimtime="00:00:38.67" resultid="2109" heatid="2208" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Luiz Cruz" birthdate="2012-10-13" gender="M" nation="BRA" license="393209" swrid="5616447" athleteid="2042" externalid="393209">
              <RESULTS>
                <RESULT eventid="1063" points="126" swimtime="00:01:53.16" resultid="2043" heatid="2134" lane="4" entrytime="00:01:54.59" entrycourse="LCM" />
                <RESULT eventid="1087" points="171" swimtime="00:03:03.64" resultid="2044" heatid="2169" lane="2" entrytime="00:03:06.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="133" swimtime="00:03:42.84" resultid="2045" heatid="2188" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1119" points="90" swimtime="00:01:50.13" resultid="2046" heatid="2204" lane="3" entrytime="00:01:48.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Fachini Kovalski" birthdate="2012-05-15" gender="M" nation="BRA" license="403404" swrid="5676297" athleteid="2087" externalid="403404">
              <RESULTS>
                <RESULT eventid="1063" points="121" swimtime="00:01:54.75" resultid="2088" heatid="2133" lane="7" />
                <RESULT eventid="1075" points="137" swimtime="00:00:45.61" resultid="2089" heatid="2151" lane="1" entrytime="00:00:50.08" entrycourse="LCM" />
                <RESULT eventid="1139" points="153" swimtime="00:00:39.08" resultid="2090" heatid="2230" lane="5" entrytime="00:00:41.87" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Vicente Lopes" birthdate="2012-03-27" gender="M" nation="BRA" license="415248" athleteid="2118" externalid="415248">
              <RESULTS>
                <RESULT eventid="1063" points="102" swimtime="00:02:01.72" resultid="2119" heatid="2133" lane="1" />
                <RESULT eventid="1075" points="66" swimtime="00:00:58.23" resultid="2120" heatid="2150" lane="3" />
                <RESULT eventid="1139" points="78" swimtime="00:00:48.90" resultid="2121" heatid="2229" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Julia Rocha" birthdate="2014-02-10" gender="F" nation="BRA" license="397158" swrid="5641767" athleteid="2047" externalid="397158">
              <RESULTS>
                <RESULT eventid="1078" points="248" swimtime="00:00:42.70" resultid="2048" heatid="2157" lane="4" entrytime="00:00:44.14" entrycourse="LCM" />
                <RESULT eventid="1090" points="223" swimtime="00:01:25.24" resultid="2049" heatid="2175" lane="3" entrytime="00:01:26.92" entrycourse="LCM" />
                <RESULT eventid="1106" points="183" swimtime="00:00:43.01" resultid="2050" heatid="2194" lane="5" entrytime="00:00:43.44" entrycourse="LCM" />
                <RESULT eventid="1126" points="281" swimtime="00:00:36.02" resultid="2051" heatid="2212" lane="3" entrytime="00:00:37.41" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Victoria De Medeiros" birthdate="2014-08-14" gender="F" nation="BRA" license="403782" swrid="5684611" athleteid="2091" externalid="403782">
              <RESULTS>
                <RESULT eventid="1066" points="126" swimtime="00:00:58.11" resultid="2092" heatid="2138" lane="1" entrytime="00:01:01.71" entrycourse="LCM" />
                <RESULT eventid="1078" points="104" swimtime="00:00:56.99" resultid="2093" heatid="2156" lane="8" entrytime="00:00:57.93" entrycourse="LCM" />
                <RESULT eventid="1106" points="82" swimtime="00:00:56.12" resultid="2094" heatid="2193" lane="2" entrytime="00:00:55.20" entrycourse="LCM" />
                <RESULT eventid="1126" points="133" swimtime="00:00:46.23" resultid="2095" heatid="2210" lane="1" entrytime="00:00:47.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Zattar" birthdate="2012-04-19" gender="F" nation="BRA" license="401736" swrid="5661351" athleteid="2074" externalid="401736">
              <RESULTS>
                <RESULT eventid="1084" status="DNS" swimtime="00:00:00.00" resultid="2075" heatid="2162" lane="4" />
                <RESULT eventid="1072" points="366" swimtime="00:00:37.53" resultid="2076" heatid="2148" lane="6" entrytime="00:00:38.62" entrycourse="LCM" />
                <RESULT eventid="1100" points="254" swimtime="00:03:18.93" resultid="2077" heatid="2183" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="350" swimtime="00:00:33.50" resultid="2078" heatid="2226" lane="4" entrytime="00:00:32.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Zanotto De Souza" birthdate="2013-08-24" gender="M" nation="BRA" license="388361" swrid="5588974" athleteid="2032" externalid="388361">
              <RESULTS>
                <RESULT eventid="1075" points="230" swimtime="00:00:38.41" resultid="2033" heatid="2152" lane="5" entrytime="00:00:40.93" entrycourse="LCM" />
                <RESULT eventid="1087" points="245" swimtime="00:02:42.84" resultid="2034" heatid="2170" lane="3" entrytime="00:02:47.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="218" swimtime="00:03:09.15" resultid="2035" heatid="2189" lane="7" entrytime="00:03:12.87" entrycourse="LCM" />
                <RESULT eventid="1139" points="246" swimtime="00:00:33.33" resultid="2036" heatid="2233" lane="2" entrytime="00:00:34.53" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Prestes Alves Pinto" birthdate="2012-01-19" gender="F" nation="BRA" license="377324" swrid="5588867" athleteid="1986" externalid="377324">
              <RESULTS>
                <RESULT eventid="1084" points="311" swimtime="00:02:46.55" resultid="1987" heatid="2165" lane="6" entrytime="00:02:50.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="327" swimtime="00:00:38.98" resultid="1988" heatid="2148" lane="1" entrytime="00:00:39.84" entrycourse="LCM" />
                <RESULT eventid="1100" points="290" swimtime="00:03:10.48" resultid="1989" heatid="2185" lane="7" entrytime="00:03:07.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="371" swimtime="00:00:32.83" resultid="1990" heatid="2226" lane="6" entrytime="00:00:33.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helloisa" lastname="De Bassani" birthdate="2012-09-23" gender="F" nation="BRA" license="403403" swrid="5676296" athleteid="2083" externalid="403403">
              <RESULTS>
                <RESULT eventid="1084" status="DNS" swimtime="00:00:00.00" resultid="2084" heatid="2163" lane="8" />
                <RESULT eventid="1072" status="DNS" swimtime="00:00:00.00" resultid="2085" heatid="2145" lane="3" entrytime="00:00:53.54" entrycourse="LCM" />
                <RESULT eventid="1136" status="DNS" swimtime="00:00:00.00" resultid="2086" heatid="2223" lane="5" entrytime="00:00:42.44" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Marini" birthdate="2014-04-09" gender="M" nation="BRA" license="382247" swrid="5684582" athleteid="1991" externalid="382247">
              <RESULTS>
                <RESULT eventid="1081" points="147" swimtime="00:00:44.54" resultid="1992" heatid="2160" lane="4" entrytime="00:00:48.54" entrycourse="LCM" />
                <RESULT eventid="1093" points="153" swimtime="00:01:27.56" resultid="1993" heatid="2179" lane="5" entrytime="00:01:31.13" entrycourse="LCM" />
                <RESULT eventid="1129" points="138" swimtime="00:00:40.41" resultid="1994" heatid="2217" lane="8" entrytime="00:00:40.52" entrycourse="LCM" />
                <RESULT eventid="1109" points="131" swimtime="00:00:43.78" resultid="1995" heatid="2196" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Gouvea" birthdate="2013-04-19" gender="M" nation="BRA" license="387378" swrid="5588729" athleteid="2018" externalid="387378">
              <RESULTS>
                <RESULT eventid="1063" points="222" swimtime="00:01:33.82" resultid="2019" heatid="2135" lane="7" entrytime="00:01:42.34" entrycourse="LCM" />
                <RESULT eventid="1087" points="198" swimtime="00:02:54.94" resultid="2020" heatid="2168" lane="1" />
                <RESULT eventid="1103" points="211" swimtime="00:03:11.34" resultid="2021" heatid="2187" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="240" swimtime="00:00:33.62" resultid="2022" heatid="2233" lane="7" entrytime="00:00:34.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="De Siqueira Machado" birthdate="2012-05-25" gender="F" nation="BRA" license="377312" swrid="5588649" athleteid="1971" externalid="377312">
              <RESULTS>
                <RESULT eventid="1060" points="254" swimtime="00:01:41.23" resultid="1972" heatid="2129" lane="6" />
                <RESULT eventid="1072" points="348" swimtime="00:00:38.18" resultid="1973" heatid="2147" lane="4" entrytime="00:00:40.85" entrycourse="LCM" />
                <RESULT eventid="1100" points="267" swimtime="00:03:15.72" resultid="1974" heatid="2182" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="385" swimtime="00:00:32.43" resultid="1975" heatid="2227" lane="1" entrytime="00:00:32.29" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Andrade Guarido" birthdate="2014-05-17" gender="M" nation="BRA" license="400031" swrid="5652873" athleteid="2065" externalid="400031">
              <RESULTS>
                <RESULT eventid="1069" points="107" swimtime="00:00:54.51" resultid="2066" heatid="2143" lane="8" entrytime="00:00:54.04" entrycourse="LCM" />
                <RESULT eventid="1093" points="144" swimtime="00:01:29.20" resultid="2067" heatid="2179" lane="6" entrytime="00:01:32.52" entrycourse="LCM" />
                <RESULT eventid="1129" points="151" swimtime="00:00:39.19" resultid="2068" heatid="2217" lane="7" entrytime="00:00:40.07" entrycourse="LCM" />
                <RESULT eventid="1109" points="53" swimtime="00:00:59.26" resultid="2069" heatid="2197" lane="3" entrytime="00:01:15.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Luiza Rocha Batista" birthdate="2013-11-24" gender="F" nation="BRA" license="387379" swrid="5588784" athleteid="2023" externalid="387379">
              <RESULTS>
                <RESULT eventid="1084" points="270" swimtime="00:02:54.46" resultid="2024" heatid="2163" lane="6" entrytime="00:03:43.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="206" swimtime="00:00:45.44" resultid="2025" heatid="2146" lane="1" entrytime="00:00:51.69" entrycourse="LCM" />
                <RESULT eventid="1116" points="129" swimtime="00:01:49.71" resultid="2026" heatid="2202" lane="4" entrytime="00:01:48.88" entrycourse="LCM" />
                <RESULT eventid="1136" points="262" swimtime="00:00:36.87" resultid="2027" heatid="2224" lane="5" entrytime="00:00:38.32" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Hugo Dos Santos" birthdate="2014-07-25" gender="M" nation="BRA" license="397420" swrid="5641766" athleteid="2057" externalid="397420">
              <RESULTS>
                <RESULT eventid="1069" points="101" swimtime="00:00:55.67" resultid="2058" heatid="2141" lane="5" entrytime="00:01:00.69" entrycourse="LCM" />
                <RESULT eventid="1093" points="130" swimtime="00:01:32.27" resultid="2059" heatid="2179" lane="2" entrytime="00:01:36.32" entrycourse="LCM" />
                <RESULT eventid="1129" points="135" swimtime="00:00:40.70" resultid="2060" heatid="2216" lane="6" entrytime="00:00:42.38" entrycourse="LCM" />
                <RESULT eventid="1109" points="62" swimtime="00:00:56.06" resultid="2061" heatid="2196" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Zanotto Souza" birthdate="2015-07-01" gender="M" nation="BRA" license="415249" athleteid="2116" externalid="415249">
              <RESULTS>
                <RESULT eventid="1129" points="92" swimtime="00:00:46.23" resultid="2117" heatid="2213" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Vitor Vicente" birthdate="2012-09-20" gender="M" nation="BRA" license="415246" athleteid="2110" externalid="415246">
              <RESULTS>
                <RESULT eventid="1087" points="99" swimtime="00:03:39.94" resultid="2111" heatid="2167" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:44.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="114" swimtime="00:00:43.09" resultid="2112" heatid="2229" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Coelho De Oliveira" birthdate="2012-11-11" gender="M" nation="BRA" license="385198" swrid="5588600" athleteid="2001" externalid="385198">
              <RESULTS>
                <RESULT eventid="1075" points="100" swimtime="00:00:50.72" resultid="2002" heatid="2150" lane="5" entrytime="00:00:57.15" entrycourse="LCM" />
                <RESULT eventid="1087" points="138" swimtime="00:03:17.00" resultid="2003" heatid="2168" lane="5" entrytime="00:03:35.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="162" swimtime="00:00:38.30" resultid="2004" heatid="2230" lane="6" entrytime="00:00:42.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Aparecida Lourenço Alves" birthdate="2013-11-06" gender="F" nation="BRA" license="387374" swrid="5588530" athleteid="2005" externalid="387374">
              <RESULTS>
                <RESULT eventid="1084" points="254" swimtime="00:02:58.10" resultid="2006" heatid="2163" lane="2" entrytime="00:03:52.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="224" swimtime="00:00:44.21" resultid="2007" heatid="2146" lane="2" entrytime="00:00:48.90" entrycourse="LCM" />
                <RESULT eventid="1136" points="306" swimtime="00:00:35.00" resultid="2008" heatid="2223" lane="2" entrytime="00:00:43.03" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Borges Piekarzievicz" birthdate="2013-09-10" gender="M" nation="BRA" license="403142" swrid="5676294" athleteid="2079" externalid="403142">
              <RESULTS>
                <RESULT eventid="1063" points="117" swimtime="00:01:56.06" resultid="2080" heatid="2134" lane="6" entrytime="00:02:02.11" entrycourse="LCM" />
                <RESULT eventid="1087" points="128" swimtime="00:03:22.32" resultid="2081" heatid="2167" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="142" swimtime="00:00:40.04" resultid="2082" heatid="2230" lane="4" entrytime="00:00:40.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Camily Moraes" birthdate="2014-07-13" gender="F" nation="BRA" license="397159" swrid="5641755" athleteid="2052" externalid="397159">
              <RESULTS>
                <RESULT eventid="1078" points="196" swimtime="00:00:46.24" resultid="2053" heatid="2157" lane="5" entrytime="00:00:47.16" entrycourse="LCM" />
                <RESULT eventid="1090" points="173" swimtime="00:01:32.70" resultid="2054" heatid="2175" lane="8" entrytime="00:01:37.93" entrycourse="LCM" />
                <RESULT eventid="1106" points="90" swimtime="00:00:54.48" resultid="2055" heatid="2191" lane="3" />
                <RESULT eventid="1126" points="229" swimtime="00:00:38.59" resultid="2056" heatid="2211" lane="4" entrytime="00:00:41.86" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Hoffmann Zoschke" birthdate="2015-03-22" gender="M" nation="BRA" license="390917" swrid="5602547" athleteid="2037" externalid="390917">
              <RESULTS>
                <RESULT eventid="1069" points="126" swimtime="00:00:51.70" resultid="2038" heatid="2142" lane="8" entrytime="00:00:59.34" entrycourse="LCM" />
                <RESULT eventid="1093" points="191" swimtime="00:01:21.32" resultid="2039" heatid="2180" lane="6" entrytime="00:01:25.11" entrycourse="LCM" />
                <RESULT eventid="1129" points="171" swimtime="00:00:37.65" resultid="2040" heatid="2218" lane="1" entrytime="00:00:37.50" entrycourse="LCM" />
                <RESULT eventid="1109" points="141" swimtime="00:00:42.69" resultid="2041" heatid="2198" lane="4" entrytime="00:00:49.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauren" lastname="Kurecki" birthdate="2014-03-06" gender="F" nation="BRA" license="377314" swrid="5602549" athleteid="1976" externalid="377314">
              <RESULTS>
                <RESULT eventid="1066" points="271" swimtime="00:00:45.01" resultid="1977" heatid="2139" lane="4" entrytime="00:00:44.66" entrycourse="LCM" />
                <RESULT eventid="1090" points="323" swimtime="00:01:15.31" resultid="1978" heatid="2175" lane="4" entrytime="00:01:18.18" entrycourse="LCM" />
                <RESULT eventid="1106" points="266" swimtime="00:00:37.95" resultid="1979" heatid="2194" lane="6" entrytime="00:00:47.50" entrycourse="LCM" />
                <RESULT eventid="1126" points="333" swimtime="00:00:34.05" resultid="1980" heatid="2212" lane="4" entrytime="00:00:33.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tais" lastname="Feltrin Martins" birthdate="2013-01-17" gender="F" nation="BRA" license="406840" swrid="5717262" athleteid="2101" externalid="406840">
              <RESULTS>
                <RESULT eventid="1084" points="86" swimtime="00:04:14.70" resultid="2102" heatid="2162" lane="1" />
                <RESULT eventid="1072" points="105" swimtime="00:00:56.87" resultid="2103" heatid="2145" lane="2" entrytime="00:01:01.05" entrycourse="LCM" />
                <RESULT eventid="1136" points="130" swimtime="00:00:46.58" resultid="2104" heatid="2222" lane="4" entrytime="00:00:46.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Soul Santos" birthdate="2016-05-11" gender="M" nation="BRA" license="415247" athleteid="2113" externalid="415247">
              <RESULTS>
                <RESULT eventid="1114" points="49" swimtime="00:01:03.93" resultid="2114" heatid="2201" lane="5" />
                <RESULT eventid="1134" points="46" swimtime="00:00:58.06" resultid="2115" heatid="2221" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Rodrigues Bortoluzzi" birthdate="2013-10-07" gender="M" nation="BRA" license="387375" swrid="5652897" athleteid="2009" externalid="387375">
              <RESULTS>
                <RESULT eventid="1075" points="153" swimtime="00:00:44.03" resultid="2010" heatid="2152" lane="1" entrytime="00:00:45.11" entrycourse="LCM" />
                <RESULT eventid="1087" points="158" swimtime="00:03:08.67" resultid="2011" heatid="2168" lane="6" entrytime="00:03:50.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="195" swimtime="00:00:36.02" resultid="2012" heatid="2232" lane="8" entrytime="00:00:37.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Strapasson" birthdate="2012-03-01" gender="M" nation="BRA" license="371377" swrid="5602585" athleteid="1966" externalid="371377">
              <RESULTS>
                <RESULT eventid="1063" points="273" swimtime="00:01:27.63" resultid="1967" heatid="2135" lane="5" entrytime="00:01:29.35" entrycourse="LCM" />
                <RESULT eventid="1087" points="278" swimtime="00:02:36.21" resultid="1968" heatid="2167" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="267" swimtime="00:02:56.92" resultid="1969" heatid="2187" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="330" swimtime="00:00:30.24" resultid="1970" heatid="2234" lane="3" entrytime="00:00:31.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mathias" lastname="Bernardo" birthdate="2014-05-17" gender="M" nation="BRA" license="387376" swrid="5652880" athleteid="2013" externalid="387376">
              <RESULTS>
                <RESULT eventid="1081" points="98" swimtime="00:00:51.01" resultid="2014" heatid="2159" lane="2" entrytime="00:00:59.85" entrycourse="LCM" />
                <RESULT eventid="1093" points="131" swimtime="00:01:32.26" resultid="2015" heatid="2179" lane="4" entrytime="00:01:30.30" entrycourse="LCM" />
                <RESULT eventid="1129" points="145" swimtime="00:00:39.79" resultid="2016" heatid="2217" lane="5" entrytime="00:00:38.12" entrycourse="LCM" />
                <RESULT eventid="1109" points="83" swimtime="00:00:50.94" resultid="2017" heatid="2195" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Ryan Rosa" birthdate="2014-01-14" gender="M" nation="BRA" license="400032" swrid="5652898" athleteid="2070" externalid="400032">
              <RESULTS>
                <RESULT eventid="1069" points="118" swimtime="00:00:52.88" resultid="2071" heatid="2142" lane="5" entrytime="00:00:55.09" entrycourse="LCM" />
                <RESULT eventid="1081" points="116" swimtime="00:00:48.27" resultid="2072" heatid="2160" lane="6" entrytime="00:00:50.32" entrycourse="LCM" />
                <RESULT eventid="1129" points="142" swimtime="00:00:40.06" resultid="2073" heatid="2215" lane="4" entrytime="00:00:45.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mathias" lastname="Lopes Batista" birthdate="2012-08-22" gender="M" nation="BRA" license="399740" swrid="5652889" athleteid="2062" externalid="399740">
              <RESULTS>
                <RESULT eventid="1075" points="185" swimtime="00:00:41.28" resultid="2063" heatid="2152" lane="3" entrytime="00:00:40.97" entrycourse="LCM" />
                <RESULT eventid="1087" points="130" swimtime="00:03:21.04" resultid="2064" heatid="2169" lane="8" entrytime="00:03:23.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Prestes" birthdate="2014-01-16" gender="M" nation="BRA" license="382249" swrid="5602574" athleteid="1996" externalid="382249">
              <RESULTS>
                <RESULT eventid="1069" points="161" swimtime="00:00:47.63" resultid="1997" heatid="2143" lane="3" entrytime="00:00:50.15" entrycourse="LCM" />
                <RESULT eventid="1093" points="180" swimtime="00:01:22.87" resultid="1998" heatid="2180" lane="2" entrytime="00:01:25.37" entrycourse="LCM" />
                <RESULT eventid="1129" points="191" swimtime="00:00:36.25" resultid="1999" heatid="2218" lane="6" entrytime="00:00:36.70" entrycourse="LCM" />
                <RESULT eventid="1109" points="83" swimtime="00:00:50.94" resultid="2000" heatid="2197" lane="4" entrytime="00:01:02.86" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lis" lastname="Cristini Harmatiuk" birthdate="2014-07-19" gender="F" nation="BRA" license="396830" swrid="5641759" athleteid="2096" externalid="396830">
              <RESULTS>
                <RESULT eventid="1066" points="194" swimtime="00:00:50.37" resultid="2097" heatid="2139" lane="7" entrytime="00:00:53.47" entrycourse="LCM" />
                <RESULT eventid="1078" points="178" swimtime="00:00:47.68" resultid="2098" heatid="2157" lane="3" entrytime="00:00:48.00" entrycourse="LCM" />
                <RESULT eventid="1106" points="136" swimtime="00:00:47.43" resultid="2099" heatid="2191" lane="6" />
                <RESULT eventid="1126" points="210" swimtime="00:00:39.67" resultid="2100" heatid="2212" lane="1" entrytime="00:00:41.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11303" nation="BRA" region="PR" clubid="1233" swrid="93760" name="Associação De Talentos Da Natação" shortname="Atn/Curitiba">
          <ATHLETES>
            <ATHLETE firstname="Arthur" lastname="Lemes Luis" birthdate="2013-10-14" gender="M" nation="BRA" license="410105" swrid="5740012" athleteid="1264" externalid="410105">
              <RESULTS>
                <RESULT eventid="1075" points="128" swimtime="00:00:46.66" resultid="1265" heatid="2151" lane="6" entrytime="00:00:47.37" entrycourse="LCM" />
                <RESULT eventid="1103" points="129" swimtime="00:03:45.57" resultid="1266" heatid="2186" lane="4" />
                <RESULT eventid="1139" points="140" swimtime="00:00:40.19" resultid="1267" heatid="2231" lane="1" entrytime="00:00:39.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Guedes Braga" birthdate="2013-04-09" gender="F" nation="BRA" license="385009" swrid="5602534" athleteid="1234" externalid="385009">
              <RESULTS>
                <RESULT eventid="1084" points="247" swimtime="00:02:59.74" resultid="1235" heatid="2165" lane="7" entrytime="00:02:54.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="252" swimtime="00:00:42.48" resultid="1236" heatid="2144" lane="3" />
                <RESULT eventid="1136" points="331" swimtime="00:00:34.11" resultid="1237" heatid="2226" lane="1" entrytime="00:00:34.05" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isaac" lastname="Zonta" birthdate="2012-11-14" gender="M" nation="BRA" license="414857" athleteid="1268" externalid="414857">
              <RESULTS>
                <RESULT eventid="1139" points="186" swimtime="00:00:36.57" resultid="1269" heatid="2228" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Leal Kuss" birthdate="2012-10-20" gender="M" nation="BRA" license="385085" swrid="5588768" athleteid="1238" externalid="385085">
              <RESULTS>
                <RESULT eventid="1119" points="190" swimtime="00:01:25.93" resultid="1239" heatid="2205" lane="7" entrytime="00:01:29.41" entrycourse="LCM" />
                <RESULT eventid="1139" points="236" swimtime="00:00:33.81" resultid="1240" heatid="2233" lane="6" entrytime="00:00:34.42" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yohanna" lastname="Vitoria Sena" birthdate="2012-01-20" gender="F" nation="BRA" license="406710" swrid="5717302" athleteid="1251" externalid="406710">
              <RESULTS>
                <RESULT eventid="1072" points="133" swimtime="00:00:52.55" resultid="1252" heatid="2146" lane="8" entrytime="00:00:51.74" entrycourse="LCM" />
                <RESULT eventid="1136" points="200" swimtime="00:00:40.34" resultid="1253" heatid="2223" lane="3" entrytime="00:00:42.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Goncalves Ghion" birthdate="2014-10-15" gender="F" nation="BRA" license="406912" swrid="5717269" athleteid="1257" externalid="406912">
              <RESULTS>
                <RESULT eventid="1066" points="124" swimtime="00:00:58.47" resultid="1258" heatid="2138" lane="7" entrytime="00:01:00.28" entrycourse="LCM" />
                <RESULT eventid="1090" points="153" swimtime="00:01:36.59" resultid="1259" heatid="2174" lane="7" entrytime="00:01:47.71" entrycourse="LCM" />
                <RESULT eventid="1126" points="182" swimtime="00:00:41.59" resultid="1260" heatid="2210" lane="7" entrytime="00:00:47.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maximilian" lastname="Hock" birthdate="2016-11-20" gender="M" nation="DEU" license="408352" athleteid="1261" externalid="408352">
              <RESULTS>
                <RESULT eventid="1124" points="71" swimtime="00:01:02.48" resultid="1262" heatid="2207" lane="4" entrytime="00:01:02.48" entrycourse="LCM" />
                <RESULT eventid="1134" points="84" swimtime="00:00:47.58" resultid="1263" heatid="2221" lane="4" entrytime="00:00:49.13" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isis" lastname="De Miranda" birthdate="2012-01-10" gender="F" nation="BRA" license="397278" swrid="5652886" athleteid="1244" externalid="397278">
              <RESULTS>
                <RESULT eventid="1084" points="311" swimtime="00:02:46.51" resultid="1245" heatid="2165" lane="3" entrytime="00:02:50.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="203" swimtime="00:01:34.31" resultid="1246" heatid="2203" lane="1" entrytime="00:01:42.30" entrycourse="LCM" />
                <RESULT eventid="1136" points="287" swimtime="00:00:35.79" resultid="1247" heatid="2225" lane="4" entrytime="00:00:34.96" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Vinicius Zonta" birthdate="2012-11-14" gender="M" nation="BRA" license="399517" swrid="5652903" athleteid="1248" externalid="399517">
              <RESULTS>
                <RESULT eventid="1087" points="256" swimtime="00:02:40.50" resultid="1249" heatid="2171" lane="1" entrytime="00:02:40.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="297" swimtime="00:00:31.32" resultid="1250" heatid="2234" lane="5" entrytime="00:00:30.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Manuela Souza" birthdate="2016-07-07" gender="F" nation="BRA" license="406759" swrid="5717282" athleteid="1254" externalid="406759">
              <RESULTS>
                <RESULT eventid="1122" points="121" swimtime="00:00:58.92" resultid="1255" heatid="2206" lane="5" entrytime="00:01:06.88" entrycourse="LCM" />
                <RESULT eventid="1132" status="DNS" swimtime="00:00:00.00" resultid="1256" heatid="2220" lane="3" entrytime="00:00:53.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Duarte De Almeida" birthdate="2013-12-09" gender="M" nation="BRA" license="385711" swrid="5588666" athleteid="1241" externalid="385711">
              <RESULTS>
                <RESULT eventid="1063" points="186" swimtime="00:01:39.58" resultid="1242" heatid="2134" lane="7" />
                <RESULT eventid="1139" points="273" swimtime="00:00:32.22" resultid="1243" heatid="2233" lane="3" entrytime="00:00:32.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16131" nation="BRA" region="PR" clubid="1857" swrid="93766" name="Associação Nadar Colombo" shortname="Equipe Nadar">
          <ATHLETES>
            <ATHLETE firstname="Tayna" lastname="Macedo Gabardo" birthdate="2012-12-01" gender="F" nation="BRA" license="406704" swrid="5717281" athleteid="1858" externalid="406704">
              <RESULTS>
                <RESULT eventid="1060" points="149" swimtime="00:02:00.70" resultid="1859" heatid="2129" lane="5" />
                <RESULT eventid="1072" points="209" swimtime="00:00:45.19" resultid="1860" heatid="2144" lane="6" />
                <RESULT eventid="1136" points="277" swimtime="00:00:36.20" resultid="1861" heatid="2225" lane="7" entrytime="00:00:37.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="1862" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Marina" lastname="Paes Schemiko" birthdate="2013-02-25" gender="F" nation="BRA" license="406918" swrid="5725995" athleteid="1881" externalid="406918">
              <RESULTS>
                <RESULT eventid="1084" points="249" swimtime="00:02:59.36" resultid="1882" heatid="2162" lane="3" />
                <RESULT eventid="1072" points="289" swimtime="00:00:40.60" resultid="1883" heatid="2145" lane="7" />
                <RESULT eventid="1100" points="257" swimtime="00:03:18.23" resultid="1884" heatid="2183" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="332" swimtime="00:00:34.09" resultid="1885" heatid="2225" lane="2" entrytime="00:00:37.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Siqueira Lopes" birthdate="2012-04-28" gender="F" nation="BRA" license="414671" athleteid="1913" externalid="414671">
              <RESULTS>
                <RESULT eventid="1116" points="173" swimtime="00:01:39.44" resultid="1914" heatid="2202" lane="3" />
                <RESULT eventid="1136" points="317" swimtime="00:00:34.60" resultid="1915" heatid="2222" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Henrique Ballatka" birthdate="2013-08-26" gender="M" nation="BRA" license="405839" swrid="5697229" athleteid="1868" externalid="405839">
              <RESULTS>
                <RESULT eventid="1063" points="89" swimtime="00:02:07.18" resultid="1869" heatid="2134" lane="1" />
                <RESULT eventid="1075" points="63" swimtime="00:00:59.13" resultid="1870" heatid="2149" lane="2" />
                <RESULT eventid="1139" points="111" swimtime="00:00:43.46" resultid="1871" heatid="2229" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Borges Duarte" birthdate="2014-02-10" gender="F" nation="BRA" license="408688" swrid="5725985" athleteid="1899" externalid="408688">
              <RESULTS>
                <RESULT eventid="1078" points="150" swimtime="00:00:50.47" resultid="1900" heatid="2156" lane="2" entrytime="00:00:54.40" entrycourse="LCM" />
                <RESULT eventid="1090" points="142" swimtime="00:01:38.93" resultid="1901" heatid="2173" lane="8" />
                <RESULT eventid="1126" points="162" swimtime="00:00:43.25" resultid="1902" heatid="2210" lane="6" entrytime="00:00:45.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Ribeiro Melo" birthdate="2013-02-25" gender="M" nation="BRA" license="406921" swrid="5717293" athleteid="1886" externalid="406921">
              <RESULTS>
                <RESULT eventid="1075" points="147" swimtime="00:00:44.57" resultid="1887" heatid="2150" lane="7" />
                <RESULT eventid="1087" points="206" swimtime="00:02:52.58" resultid="1888" heatid="2169" lane="5" entrytime="00:02:59.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="156" swimtime="00:03:31.55" resultid="1889" heatid="2186" lane="3" />
                <RESULT eventid="1139" points="180" swimtime="00:00:36.98" resultid="1890" heatid="2232" lane="1" entrytime="00:00:36.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Sprengel Betim" birthdate="2012-08-17" gender="F" nation="BRA" license="385011" swrid="5588922" athleteid="1872" externalid="385011">
              <RESULTS>
                <RESULT eventid="1060" points="262" swimtime="00:01:40.11" resultid="1873" heatid="2129" lane="7" />
                <RESULT eventid="1084" points="293" swimtime="00:02:49.87" resultid="1874" heatid="2164" lane="7" entrytime="00:03:13.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="213" swimtime="00:01:32.83" resultid="1875" heatid="2202" lane="5" />
                <RESULT eventid="1136" points="277" swimtime="00:00:36.21" resultid="1876" heatid="2224" lane="4" entrytime="00:00:37.96" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Cavalcante Pierin" birthdate="2015-03-31" gender="M" nation="BRA" license="408082" swrid="5725986" athleteid="1908" externalid="408082">
              <RESULTS>
                <RESULT eventid="1081" points="93" swimtime="00:00:51.91" resultid="1909" heatid="2160" lane="7" entrytime="00:00:50.92" entrycourse="LCM" />
                <RESULT eventid="1093" points="137" swimtime="00:01:30.80" resultid="1910" heatid="2176" lane="4" />
                <RESULT eventid="1129" points="121" swimtime="00:00:42.26" resultid="1911" heatid="2216" lane="2" entrytime="00:00:43.57" entrycourse="LCM" />
                <RESULT eventid="1109" points="43" swimtime="00:01:03.42" resultid="1912" heatid="2195" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Schneider Yazbek" birthdate="2013-03-07" gender="F" nation="BRA" license="378329" swrid="5588907" athleteid="1863" externalid="378329">
              <RESULTS>
                <RESULT eventid="1060" points="244" swimtime="00:01:42.62" resultid="1864" heatid="2129" lane="2" />
                <RESULT eventid="1084" points="367" swimtime="00:02:37.49" resultid="1865" heatid="2166" lane="8" entrytime="00:02:42.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1100" points="319" swimtime="00:03:04.58" resultid="1866" heatid="2185" lane="1" entrytime="00:03:09.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1116" points="223" swimtime="00:01:31.41" resultid="1867" heatid="2203" lane="2" entrytime="00:01:36.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Samuel" lastname="Melo Lima" birthdate="2015-10-30" gender="M" nation="BRA" license="406933" swrid="5725994" athleteid="1895" externalid="406933">
              <RESULTS>
                <RESULT eventid="1069" points="73" swimtime="00:01:02.06" resultid="1896" heatid="2140" lane="5" />
                <RESULT eventid="1081" points="75" swimtime="00:00:55.81" resultid="1897" heatid="2158" lane="6" />
                <RESULT eventid="1129" points="72" swimtime="00:00:50.19" resultid="1898" heatid="2214" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Manoel Forte" birthdate="2013-01-13" gender="M" nation="BRA" license="414859" athleteid="1916" externalid="414859">
              <RESULTS>
                <RESULT eventid="1075" points="96" swimtime="00:00:51.42" resultid="1917" heatid="2150" lane="6" />
                <RESULT eventid="1139" points="86" swimtime="00:00:47.34" resultid="1918" heatid="2228" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Zanatta Duda" birthdate="2013-08-28" gender="F" nation="BRA" license="406914" swrid="5717306" athleteid="1877" externalid="406914">
              <RESULTS>
                <RESULT eventid="1084" points="154" swimtime="00:03:30.42" resultid="1878" heatid="2162" lane="8" />
                <RESULT eventid="1072" points="188" swimtime="00:00:46.87" resultid="1879" heatid="2146" lane="3" entrytime="00:00:47.26" entrycourse="LCM" />
                <RESULT eventid="1136" points="178" swimtime="00:00:41.94" resultid="1880" heatid="2223" lane="6" entrytime="00:00:42.89" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="De Ormeno" birthdate="2014-04-02" gender="M" nation="BRA" license="408702" swrid="5740009" athleteid="1903" externalid="408702">
              <RESULTS>
                <RESULT eventid="1081" points="201" swimtime="00:00:40.16" resultid="1904" heatid="2161" lane="3" entrytime="00:00:43.94" entrycourse="LCM" />
                <RESULT eventid="1093" points="229" swimtime="00:01:16.58" resultid="1905" heatid="2180" lane="5" entrytime="00:01:21.54" entrycourse="LCM" />
                <RESULT eventid="1129" points="223" swimtime="00:00:34.47" resultid="1906" heatid="2218" lane="3" entrytime="00:00:36.20" entrycourse="LCM" />
                <RESULT eventid="1109" points="121" swimtime="00:00:44.96" resultid="1907" heatid="2197" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="De Andrade" birthdate="2015-12-24" gender="M" nation="BRA" license="406922" swrid="5740008" athleteid="1891" externalid="406922">
              <RESULTS>
                <RESULT eventid="1081" points="87" swimtime="00:00:53.03" resultid="1892" heatid="2159" lane="4" entrytime="00:00:54.51" entrycourse="LCM" />
                <RESULT eventid="1093" points="87" swimtime="00:01:45.39" resultid="1893" heatid="2178" lane="6" entrytime="00:01:44.50" entrycourse="LCM" />
                <RESULT eventid="1129" points="109" swimtime="00:00:43.71" resultid="1894" heatid="2215" lane="3" entrytime="00:00:46.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13038" nation="BRA" region="PR" clubid="1186" swrid="93759" name="Associação De Pais E Atletas De Natação Ws/Crb" shortname="Apan/Ws">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Dos Santos" birthdate="2013-06-26" gender="F" nation="BRA" license="387512" swrid="5588662" athleteid="1203" externalid="387512">
              <RESULTS>
                <RESULT eventid="1084" status="DNS" swimtime="00:00:00.00" resultid="1204" heatid="2164" lane="3" entrytime="00:03:05.03" entrycourse="LCM" />
                <RESULT eventid="1072" points="245" swimtime="00:00:42.92" resultid="1205" heatid="2147" lane="6" entrytime="00:00:44.32" entrycourse="LCM" />
                <RESULT eventid="1136" points="305" swimtime="00:00:35.07" resultid="1206" heatid="2223" lane="8" entrytime="00:00:44.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Bernardi Iurk" birthdate="2012-04-14" gender="M" nation="BRA" license="408687" swrid="5725984" athleteid="1191" externalid="408687">
              <RESULTS>
                <RESULT eventid="1063" points="130" swimtime="00:01:52.11" resultid="1192" heatid="2132" lane="5" />
                <RESULT eventid="1075" points="147" swimtime="00:00:44.58" resultid="1193" heatid="2149" lane="5" />
                <RESULT eventid="1139" points="205" swimtime="00:00:35.42" resultid="1194" heatid="2231" lane="5" entrytime="00:00:38.11" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leon" lastname="Bernardo Bello" birthdate="2014-11-23" gender="M" nation="BRA" license="400324" swrid="5717246" athleteid="1211" externalid="400324">
              <RESULTS>
                <RESULT eventid="1069" points="118" swimtime="00:00:52.84" resultid="1212" heatid="2142" lane="6" entrytime="00:00:55.43" entrycourse="LCM" />
                <RESULT eventid="1093" points="123" swimtime="00:01:34.02" resultid="1213" heatid="2179" lane="7" entrytime="00:01:36.77" entrycourse="LCM" />
                <RESULT eventid="1129" points="166" swimtime="00:00:37.98" resultid="1214" heatid="2217" lane="1" entrytime="00:00:40.45" entrycourse="LCM" />
                <RESULT eventid="1109" points="55" swimtime="00:00:58.24" resultid="1215" heatid="2196" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Bobko Ganacim" birthdate="2013-08-02" gender="F" nation="BRA" license="397332" swrid="5641754" athleteid="1200" externalid="397332">
              <RESULTS>
                <RESULT eventid="1060" points="136" swimtime="00:02:04.47" resultid="1201" heatid="2129" lane="4" />
                <RESULT eventid="1072" points="148" swimtime="00:00:50.77" resultid="1202" heatid="2145" lane="5" entrytime="00:00:52.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Gabriel Cabral" birthdate="2014-02-11" gender="M" nation="BRA" license="415259" athleteid="1229" externalid="415259">
              <RESULTS>
                <RESULT eventid="1081" points="107" swimtime="00:00:49.57" resultid="1230" heatid="2158" lane="3" />
                <RESULT eventid="1093" points="130" swimtime="00:01:32.40" resultid="1231" heatid="2177" lane="7" />
                <RESULT eventid="1129" points="125" swimtime="00:00:41.76" resultid="1232" heatid="2213" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Bernardi Iurk" birthdate="2012-04-14" gender="M" nation="BRA" license="406940" swrid="5717245" athleteid="1187" externalid="406940">
              <RESULTS>
                <RESULT eventid="1075" points="156" swimtime="00:00:43.71" resultid="1188" heatid="2151" lane="3" entrytime="00:00:47.12" entrycourse="LCM" />
                <RESULT eventid="1087" points="227" swimtime="00:02:47.20" resultid="1189" heatid="2167" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="238" swimtime="00:00:33.74" resultid="1190" heatid="2231" lane="4" entrytime="00:00:37.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Cravcenco Marcondes" birthdate="2012-06-23" gender="F" nation="BRA" license="406866" swrid="5725987" athleteid="1216" externalid="406866">
              <RESULTS>
                <RESULT eventid="1084" points="191" swimtime="00:03:15.75" resultid="1217" heatid="2162" lane="2" />
                <RESULT eventid="1072" points="253" swimtime="00:00:42.42" resultid="1218" heatid="2147" lane="7" entrytime="00:00:44.79" entrycourse="LCM" />
                <RESULT eventid="1136" points="266" swimtime="00:00:36.67" resultid="1219" heatid="2224" lane="6" entrytime="00:00:40.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Gramms Dallarosa" birthdate="2015-01-14" gender="F" nation="BRA" license="406868" swrid="5717270" athleteid="1220" externalid="406868">
              <RESULTS>
                <RESULT eventid="1066" points="102" swimtime="00:01:02.28" resultid="1221" heatid="2137" lane="2" entrytime="00:01:10.36" entrycourse="LCM" />
                <RESULT eventid="1090" points="126" swimtime="00:01:42.91" resultid="1222" heatid="2174" lane="1" entrytime="00:01:49.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Da Reginalda" birthdate="2012-11-09" gender="M" nation="BRA" license="400275" swrid="5717253" athleteid="1207" externalid="400275">
              <RESULTS>
                <RESULT eventid="1075" points="259" swimtime="00:00:36.91" resultid="1208" heatid="2150" lane="1" />
                <RESULT eventid="1087" points="235" swimtime="00:02:45.06" resultid="1209" heatid="2168" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="280" swimtime="00:00:31.93" resultid="1210" heatid="2232" lane="5" entrytime="00:00:35.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Ferreira" birthdate="2012-12-29" gender="F" nation="BRA" license="382235" swrid="5602538" athleteid="1195" externalid="382235">
              <RESULTS>
                <RESULT eventid="1084" points="278" swimtime="00:02:52.90" resultid="1196" heatid="2162" lane="7" />
                <RESULT eventid="1072" points="274" swimtime="00:00:41.32" resultid="1197" heatid="2146" lane="6" entrytime="00:00:48.31" entrycourse="LCM" />
                <RESULT eventid="1116" points="195" swimtime="00:01:35.54" resultid="1198" heatid="2203" lane="7" entrytime="00:01:41.46" entrycourse="LCM" />
                <RESULT eventid="1136" points="307" swimtime="00:00:34.99" resultid="1199" heatid="2224" lane="7" entrytime="00:00:40.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Ancai Freire" birthdate="2012-08-11" gender="M" nation="BRA" license="415258" athleteid="1226" externalid="415258">
              <RESULTS>
                <RESULT eventid="1075" points="71" swimtime="00:00:56.78" resultid="1227" heatid="2149" lane="4" />
                <RESULT eventid="1139" points="90" swimtime="00:00:46.55" resultid="1228" heatid="2230" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Iasmim" lastname="Ferenczuk" birthdate="2013-06-06" gender="F" nation="BRA" license="414654" athleteid="1223" externalid="414654">
              <RESULTS>
                <RESULT eventid="1072" points="116" swimtime="00:00:54.92" resultid="1224" heatid="2145" lane="1" />
                <RESULT eventid="1136" points="151" swimtime="00:00:44.32" resultid="1225" heatid="2222" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="UNATTACHED">
          <OFFICIALS>
            <OFFICIAL officialid="2316" firstname="Felipe" gender="M" lastname="Oliveira Mendonça" />
          </OFFICIALS>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
