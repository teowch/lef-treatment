<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.78979">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Curitiba" name="Torneio Regional da 1ª Região (Infantil/Sênior)" course="LCM" deadline="2024-03-17" entrystartdate="2024-03-12" entrytype="INVITATION" hostclub="Clube Curitibano" hostclub.url="https://clubecuritibano.com.br/" number="38302" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/evento/natacao/38302/" startmethod="1" timing="AUTOMATIC" masters="F" withdrawuntil="2024-03-20" state="PR" nation="BRA">
      <AGEDATE value="2024-03-23" type="YEAR" />
      <POOL name="Parque Aquático do Clube Curitibano" lanemin="1" lanemax="8" />
      <FACILITY city="Curitiba" name="Parque Aquático do Clube Curitibano" nation="BRA" state="PR" street="Avenida Presidente Getúlio Vargas, 2857" street2="Água Verde" zip="80240-040" />
      <POINTTABLE pointtableid="3017" name="FINA Point Scoring" version="2024" />
      <QUALIFY from="2023-03-23" until="2024-03-22" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-03-23" daytime="09:10" endtime="12:17" number="1" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1060" daytime="09:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1778" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1063" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1064" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1065" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1066" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1067" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1821" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2246" daytime="09:10" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1068" daytime="09:16" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1069" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1731" />
                    <RANKING order="2" place="2" resultid="1749" />
                    <RANKING order="3" place="3" resultid="1714" />
                    <RANKING order="4" place="4" resultid="1737" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1070" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1374" />
                    <RANKING order="2" place="2" resultid="1658" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1230" />
                    <RANKING order="2" place="2" resultid="1339" />
                    <RANKING order="3" place="3" resultid="1960" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1073" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1074" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1496" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2247" daytime="09:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2248" daytime="09:24" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1076" daytime="09:30" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1077" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1742" />
                    <RANKING order="2" place="2" resultid="1725" />
                    <RANKING order="3" place="3" resultid="1698" />
                    <RANKING order="4" place="4" resultid="1720" />
                    <RANKING order="5" place="5" resultid="1917" />
                    <RANKING order="6" place="6" resultid="1770" />
                    <RANKING order="7" place="7" resultid="1830" />
                    <RANKING order="8" place="8" resultid="1825" />
                    <RANKING order="9" place="9" resultid="1982" />
                    <RANKING order="10" place="10" resultid="1709" />
                    <RANKING order="11" place="11" resultid="2186" />
                    <RANKING order="12" place="12" resultid="1426" />
                    <RANKING order="13" place="-1" resultid="2145" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1609" />
                    <RANKING order="2" place="2" resultid="1653" />
                    <RANKING order="3" place="3" resultid="1615" />
                    <RANKING order="4" place="4" resultid="1621" />
                    <RANKING order="5" place="5" resultid="1641" />
                    <RANKING order="6" place="6" resultid="1525" />
                    <RANKING order="7" place="7" resultid="2194" />
                    <RANKING order="8" place="8" resultid="1804" />
                    <RANKING order="9" place="9" resultid="2226" />
                    <RANKING order="10" place="10" resultid="1996" />
                    <RANKING order="11" place="11" resultid="1865" />
                    <RANKING order="12" place="12" resultid="1663" />
                    <RANKING order="13" place="13" resultid="2241" />
                    <RANKING order="14" place="14" resultid="1289" />
                    <RANKING order="15" place="15" resultid="2237" />
                    <RANKING order="16" place="16" resultid="2047" />
                    <RANKING order="17" place="17" resultid="2042" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1521" />
                    <RANKING order="2" place="2" resultid="1493" />
                    <RANKING order="3" place="3" resultid="2098" />
                    <RANKING order="4" place="4" resultid="1245" />
                    <RANKING order="5" place="5" resultid="2182" />
                    <RANKING order="6" place="6" resultid="1577" />
                    <RANKING order="7" place="7" resultid="1902" />
                    <RANKING order="8" place="8" resultid="2130" />
                    <RANKING order="9" place="9" resultid="2141" />
                    <RANKING order="10" place="10" resultid="1385" />
                    <RANKING order="11" place="11" resultid="2124" />
                    <RANKING order="12" place="12" resultid="1447" />
                    <RANKING order="13" place="-1" resultid="1487" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1080" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2017" />
                    <RANKING order="2" place="2" resultid="2063" />
                    <RANKING order="3" place="3" resultid="1293" />
                    <RANKING order="4" place="4" resultid="1950" />
                    <RANKING order="5" place="5" resultid="2052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1532" />
                    <RANKING order="2" place="2" resultid="1515" />
                    <RANKING order="3" place="3" resultid="1922" />
                    <RANKING order="4" place="4" resultid="1403" />
                    <RANKING order="5" place="5" resultid="1398" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2108" />
                    <RANKING order="2" place="2" resultid="2027" />
                    <RANKING order="3" place="-1" resultid="1879" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1083" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2037" />
                    <RANKING order="2" place="2" resultid="2013" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2249" daytime="09:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2250" daytime="09:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2251" daytime="09:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2252" daytime="09:44" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2253" daytime="09:48" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2254" daytime="09:52" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2255" daytime="09:56" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="2256" daytime="09:58" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1084" daytime="10:04" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1085" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1759" />
                    <RANKING order="2" place="2" resultid="1683" />
                    <RANKING order="3" place="3" resultid="1677" />
                    <RANKING order="4" place="4" resultid="1688" />
                    <RANKING order="5" place="5" resultid="1748" />
                    <RANKING order="6" place="6" resultid="1459" />
                    <RANKING order="7" place="7" resultid="1693" />
                    <RANKING order="8" place="8" resultid="2161" />
                    <RANKING order="9" place="9" resultid="2178" />
                    <RANKING order="10" place="10" resultid="2025" />
                    <RANKING order="11" place="11" resultid="1796" />
                    <RANKING order="12" place="12" resultid="1787" />
                    <RANKING order="13" place="13" resultid="2189" />
                    <RANKING order="14" place="14" resultid="2078" />
                    <RANKING order="15" place="15" resultid="2212" />
                    <RANKING order="16" place="16" resultid="1704" />
                    <RANKING order="17" place="17" resultid="1369" />
                    <RANKING order="18" place="18" resultid="2220" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1086" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1626" />
                    <RANKING order="2" place="2" resultid="1754" />
                    <RANKING order="3" place="3" resultid="1813" />
                    <RANKING order="4" place="4" resultid="1668" />
                    <RANKING order="5" place="5" resultid="1636" />
                    <RANKING order="6" place="6" resultid="1631" />
                    <RANKING order="7" place="7" resultid="1595" />
                    <RANKING order="8" place="8" resultid="2152" />
                    <RANKING order="9" place="9" resultid="1646" />
                    <RANKING order="10" place="10" resultid="2201" />
                    <RANKING order="11" place="11" resultid="2164" />
                    <RANKING order="12" place="12" resultid="1435" />
                    <RANKING order="13" place="13" resultid="1965" />
                    <RANKING order="14" place="14" resultid="1390" />
                    <RANKING order="15" place="15" resultid="2209" />
                    <RANKING order="16" place="16" resultid="1930" />
                    <RANKING order="17" place="17" resultid="1443" />
                    <RANKING order="18" place="18" resultid="2082" />
                    <RANKING order="19" place="19" resultid="1970" />
                    <RANKING order="20" place="20" resultid="1411" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1224" />
                    <RANKING order="2" place="2" resultid="1504" />
                    <RANKING order="3" place="3" resultid="1529" />
                    <RANKING order="4" place="4" resultid="1959" />
                    <RANKING order="5" place="5" resultid="2118" />
                    <RANKING order="6" place="6" resultid="1259" />
                    <RANKING order="7" place="7" resultid="2205" />
                    <RANKING order="8" place="8" resultid="2134" />
                    <RANKING order="9" place="9" resultid="1871" />
                    <RANKING order="10" place="10" resultid="1406" />
                    <RANKING order="11" place="11" resultid="2010" />
                    <RANKING order="12" place="12" resultid="2230" />
                    <RANKING order="13" place="13" resultid="1430" />
                    <RANKING order="14" place="14" resultid="1473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1501" />
                    <RANKING order="2" place="2" resultid="2127" />
                    <RANKING order="3" place="3" resultid="1800" />
                    <RANKING order="4" place="4" resultid="1860" />
                    <RANKING order="5" place="5" resultid="1886" />
                    <RANKING order="6" place="6" resultid="2112" />
                    <RANKING order="7" place="7" resultid="1992" />
                    <RANKING order="8" place="8" resultid="2093" />
                    <RANKING order="9" place="9" resultid="1414" />
                    <RANKING order="10" place="10" resultid="1480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1089" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1536" />
                    <RANKING order="2" place="2" resultid="2104" />
                    <RANKING order="3" place="3" resultid="2058" />
                    <RANKING order="4" place="4" resultid="2233" />
                    <RANKING order="5" place="5" resultid="1907" />
                    <RANKING order="6" place="6" resultid="2073" />
                    <RANKING order="7" place="7" resultid="1912" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1846" />
                    <RANKING order="2" place="2" resultid="2137" />
                    <RANKING order="3" place="3" resultid="1856" />
                    <RANKING order="4" place="4" resultid="2000" />
                    <RANKING order="5" place="5" resultid="2175" />
                    <RANKING order="6" place="6" resultid="1351" />
                    <RANKING order="7" place="7" resultid="1451" />
                    <RANKING order="8" place="8" resultid="2032" />
                    <RANKING order="9" place="9" resultid="1543" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1808" />
                    <RANKING order="2" place="2" resultid="2005" />
                    <RANKING order="3" place="3" resultid="1347" />
                    <RANKING order="4" place="4" resultid="1356" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2257" daytime="10:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2258" daytime="10:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2259" daytime="10:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2260" daytime="10:14" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2261" daytime="10:18" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2262" daytime="10:22" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2263" daytime="10:26" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="2264" daytime="10:30" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="2265" daytime="10:34" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="2266" daytime="10:36" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="2267" daytime="10:40" number="11" order="11" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1092" daytime="10:44" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1093" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1652" />
                    <RANKING order="2" place="2" resultid="2168" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1095" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1096" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1097" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1098" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1099" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1820" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2268" daytime="10:44" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1100" daytime="10:48" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1101" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1713" />
                    <RANKING order="2" place="2" resultid="1682" />
                    <RANKING order="3" place="3" resultid="1786" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1103" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1229" />
                    <RANKING order="2" place="2" resultid="1840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1104" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1553" />
                    <RANKING order="2" place="2" resultid="1421" />
                    <RANKING order="3" place="-1" resultid="1817" />
                    <RANKING order="4" place="-1" resultid="2092" />
                    <RANKING order="5" place="-1" resultid="1508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1105" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1954" />
                    <RANKING order="2" place="-1" resultid="1518" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1107" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1362" />
                    <RANKING order="2" place="2" resultid="2004" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2269" daytime="10:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2270" daytime="10:54" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1108" daytime="10:58" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1109" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1741" />
                    <RANKING order="2" place="2" resultid="1724" />
                    <RANKING order="3" place="3" resultid="1278" />
                    <RANKING order="4" place="4" resultid="1769" />
                    <RANKING order="5" place="5" resultid="1824" />
                    <RANKING order="6" place="6" resultid="1916" />
                    <RANKING order="7" place="7" resultid="1719" />
                    <RANKING order="8" place="8" resultid="1425" />
                    <RANKING order="9" place="9" resultid="1981" />
                    <RANKING order="10" place="10" resultid="1455" />
                    <RANKING order="11" place="11" resultid="1330" />
                    <RANKING order="12" place="12" resultid="2223" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1110" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1614" />
                    <RANKING order="2" place="2" resultid="1605" />
                    <RANKING order="3" place="3" resultid="1305" />
                    <RANKING order="4" place="4" resultid="1620" />
                    <RANKING order="5" place="5" resultid="1864" />
                    <RANKING order="6" place="6" resultid="1640" />
                    <RANKING order="7" place="7" resultid="1995" />
                    <RANKING order="8" place="8" resultid="2236" />
                    <RANKING order="9" place="9" resultid="1765" />
                    <RANKING order="10" place="10" resultid="2240" />
                    <RANKING order="11" place="11" resultid="1662" />
                    <RANKING order="12" place="12" resultid="2041" />
                    <RANKING order="13" place="13" resultid="1939" />
                    <RANKING order="14" place="14" resultid="1926" />
                    <RANKING order="15" place="15" resultid="2046" />
                    <RANKING order="16" place="16" resultid="1324" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1111" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1334" />
                    <RANKING order="2" place="2" resultid="1244" />
                    <RANKING order="3" place="3" resultid="1384" />
                    <RANKING order="4" place="4" resultid="1253" />
                    <RANKING order="5" place="5" resultid="2140" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1112" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1837" />
                    <RANKING order="2" place="2" resultid="1490" />
                    <RANKING order="3" place="3" resultid="2016" />
                    <RANKING order="4" place="4" resultid="1292" />
                    <RANKING order="5" place="5" resultid="1949" />
                    <RANKING order="6" place="6" resultid="2051" />
                    <RANKING order="7" place="7" resultid="1312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2101" />
                    <RANKING order="2" place="2" resultid="1249" />
                    <RANKING order="3" place="3" resultid="1921" />
                    <RANKING order="4" place="4" resultid="1402" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1114" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1286" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1115" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2036" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2271" daytime="10:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2272" daytime="11:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2273" daytime="11:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2274" daytime="11:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2275" daytime="11:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2276" daytime="11:14" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1116" daytime="11:16" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1117" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1758" />
                    <RANKING order="2" place="2" resultid="2148" />
                    <RANKING order="3" place="3" resultid="1321" />
                    <RANKING order="4" place="4" resultid="1268" />
                    <RANKING order="5" place="5" resultid="1736" />
                    <RANKING order="6" place="6" resultid="1692" />
                    <RANKING order="7" place="7" resultid="2024" />
                    <RANKING order="8" place="8" resultid="1676" />
                    <RANKING order="9" place="9" resultid="1935" />
                    <RANKING order="10" place="10" resultid="1703" />
                    <RANKING order="11" place="11" resultid="2077" />
                    <RANKING order="12" place="12" resultid="1795" />
                    <RANKING order="13" place="13" resultid="1327" />
                    <RANKING order="14" place="14" resultid="1477" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1118" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1812" />
                    <RANKING order="2" place="2" resultid="1630" />
                    <RANKING order="3" place="3" resultid="1600" />
                    <RANKING order="4" place="4" resultid="1625" />
                    <RANKING order="5" place="5" resultid="1753" />
                    <RANKING order="6" place="6" resultid="1635" />
                    <RANKING order="7" place="7" resultid="1389" />
                    <RANKING order="8" place="8" resultid="2208" />
                    <RANKING order="9" place="9" resultid="1929" />
                    <RANKING order="10" place="10" resultid="1410" />
                    <RANKING order="11" place="11" resultid="1462" />
                    <RANKING order="12" place="12" resultid="1442" />
                    <RANKING order="13" place="13" resultid="1434" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1338" />
                    <RANKING order="2" place="2" resultid="1223" />
                    <RANKING order="3" place="3" resultid="1853" />
                    <RANKING order="4" place="4" resultid="2121" />
                    <RANKING order="5" place="5" resultid="1583" />
                    <RANKING order="6" place="6" resultid="1958" />
                    <RANKING order="7" place="7" resultid="1870" />
                    <RANKING order="8" place="8" resultid="1562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1120" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1500" />
                    <RANKING order="2" place="2" resultid="1587" />
                    <RANKING order="3" place="3" resultid="1559" />
                    <RANKING order="4" place="4" resultid="1550" />
                    <RANKING order="5" place="5" resultid="1302" />
                    <RANKING order="6" place="6" resultid="1547" />
                    <RANKING order="7" place="-1" resultid="1420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1121" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1850" />
                    <RANKING order="2" place="2" resultid="2244" />
                    <RANKING order="3" place="3" resultid="1906" />
                    <RANKING order="4" place="4" resultid="1911" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1123" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2277" daytime="11:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2278" daytime="11:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2279" daytime="11:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2280" daytime="11:26" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2281" daytime="11:30" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2282" daytime="11:32" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1124" daytime="11:36" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1125" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1718" />
                    <RANKING order="2" place="2" resultid="1697" />
                    <RANKING order="3" place="3" resultid="1829" />
                    <RANKING order="4" place="4" resultid="2185" />
                    <RANKING order="5" place="5" resultid="1708" />
                    <RANKING order="6" place="6" resultid="1893" />
                    <RANKING order="7" place="7" resultid="1318" />
                    <RANKING order="8" place="8" resultid="2216" />
                    <RANKING order="9" place="-1" resultid="2144" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1973" />
                    <RANKING order="2" place="2" resultid="1803" />
                    <RANKING order="3" place="3" resultid="1524" />
                    <RANKING order="4" place="4" resultid="2193" />
                    <RANKING order="5" place="5" resultid="2197" />
                    <RANKING order="6" place="6" resultid="1863" />
                    <RANKING order="7" place="7" resultid="1651" />
                    <RANKING order="8" place="8" resultid="1764" />
                    <RANKING order="9" place="9" resultid="1604" />
                    <RANKING order="10" place="10" resultid="1271" />
                    <RANKING order="11" place="11" resultid="2086" />
                    <RANKING order="12" place="12" resultid="1897" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1127" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1568" />
                    <RANKING order="2" place="2" resultid="1571" />
                    <RANKING order="3" place="3" resultid="1381" />
                    <RANKING order="4" place="4" resultid="1901" />
                    <RANKING order="5" place="5" resultid="1889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1484" />
                    <RANKING order="2" place="2" resultid="1774" />
                    <RANKING order="3" place="3" resultid="2062" />
                    <RANKING order="4" place="4" resultid="1296" />
                    <RANKING order="5" place="5" resultid="2115" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1514" />
                    <RANKING order="2" place="2" resultid="1299" />
                    <RANKING order="3" place="3" resultid="1397" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1130" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1843" />
                    <RANKING order="2" place="2" resultid="1240" />
                    <RANKING order="3" place="-1" resultid="1878" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2283" daytime="11:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2284" daytime="11:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2285" daytime="11:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2286" daytime="11:44" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2287" daytime="11:46" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1132" daytime="11:50" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1133" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1730" />
                    <RANKING order="2" place="2" resultid="1687" />
                    <RANKING order="3" place="3" resultid="1747" />
                    <RANKING order="4" place="4" resultid="2160" />
                    <RANKING order="5" place="5" resultid="1267" />
                    <RANKING order="6" place="6" resultid="2156" />
                    <RANKING order="7" place="7" resultid="1458" />
                    <RANKING order="8" place="8" resultid="1393" />
                    <RANKING order="9" place="9" resultid="2076" />
                    <RANKING order="10" place="10" resultid="2023" />
                    <RANKING order="11" place="11" resultid="1794" />
                    <RANKING order="12" place="12" resultid="1702" />
                    <RANKING order="13" place="13" resultid="1476" />
                    <RANKING order="14" place="14" resultid="2219" />
                    <RANKING order="15" place="-1" resultid="1934" />
                    <RANKING order="16" place="-1" resultid="1785" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1134" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1373" />
                    <RANKING order="2" place="2" resultid="1645" />
                    <RANKING order="3" place="3" resultid="1594" />
                    <RANKING order="4" place="4" resultid="1667" />
                    <RANKING order="5" place="5" resultid="1388" />
                    <RANKING order="6" place="6" resultid="1657" />
                    <RANKING order="7" place="7" resultid="1964" />
                    <RANKING order="8" place="8" resultid="1438" />
                    <RANKING order="9" place="9" resultid="2081" />
                    <RANKING order="10" place="10" resultid="1599" />
                    <RANKING order="11" place="11" resultid="1441" />
                    <RANKING order="12" place="12" resultid="1969" />
                    <RANKING order="13" place="-1" resultid="1433" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1228" />
                    <RANKING order="2" place="2" resultid="1574" />
                    <RANKING order="3" place="3" resultid="1365" />
                    <RANKING order="4" place="4" resultid="1377" />
                    <RANKING order="5" place="5" resultid="2133" />
                    <RANKING order="6" place="6" resultid="1405" />
                    <RANKING order="7" place="7" resultid="2009" />
                    <RANKING order="8" place="-1" resultid="1565" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1511" />
                    <RANKING order="2" place="2" resultid="1834" />
                    <RANKING order="3" place="3" resultid="1782" />
                    <RANKING order="4" place="4" resultid="1791" />
                    <RANKING order="5" place="5" resultid="1875" />
                    <RANKING order="6" place="6" resultid="1991" />
                    <RANKING order="7" place="7" resultid="1466" />
                    <RANKING order="8" place="8" resultid="1309" />
                    <RANKING order="9" place="-1" resultid="1556" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1137" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1539" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1263" />
                    <RANKING order="2" place="2" resultid="1986" />
                    <RANKING order="3" place="3" resultid="1275" />
                    <RANKING order="4" place="4" resultid="1450" />
                    <RANKING order="5" place="5" resultid="1282" />
                    <RANKING order="6" place="6" resultid="2031" />
                    <RANKING order="7" place="-1" resultid="2172" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1139" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1590" />
                    <RANKING order="2" place="2" resultid="1234" />
                    <RANKING order="3" place="3" resultid="1359" />
                    <RANKING order="4" place="4" resultid="1237" />
                    <RANKING order="5" place="5" resultid="1355" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2288" daytime="11:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2289" daytime="11:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2290" daytime="11:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2291" daytime="11:58" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2292" daytime="12:02" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2293" daytime="12:04" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2294" daytime="12:06" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="2295" daytime="12:10" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-03-23" daytime="16:40" endtime="20:35" number="2" officialmeeting="16:00" warmupfrom="15:30" warmupuntil="16:30">
          <EVENTS>
            <EVENT eventid="1140" daytime="16:40" gender="F" number="11" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1141" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1745" />
                    <RANKING order="2" place="2" resultid="1728" />
                    <RANKING order="3" place="3" resultid="1280" />
                    <RANKING order="4" place="4" resultid="1700" />
                    <RANKING order="5" place="5" resultid="1722" />
                    <RANKING order="6" place="6" resultid="1772" />
                    <RANKING order="7" place="7" resultid="1456" />
                    <RANKING order="8" place="8" resultid="1984" />
                    <RANKING order="9" place="9" resultid="1895" />
                    <RANKING order="10" place="10" resultid="1331" />
                    <RANKING order="11" place="11" resultid="2224" />
                    <RANKING order="12" place="12" resultid="1316" />
                    <RANKING order="13" place="-1" resultid="1428" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1612" />
                    <RANKING order="2" place="2" resultid="1618" />
                    <RANKING order="3" place="3" resultid="2228" />
                    <RANKING order="4" place="4" resultid="1623" />
                    <RANKING order="5" place="5" resultid="1806" />
                    <RANKING order="6" place="6" resultid="1307" />
                    <RANKING order="7" place="7" resultid="1607" />
                    <RANKING order="8" place="8" resultid="1998" />
                    <RANKING order="9" place="9" resultid="1767" />
                    <RANKING order="10" place="10" resultid="1273" />
                    <RANKING order="11" place="11" resultid="2049" />
                    <RANKING order="12" place="12" resultid="1940" />
                    <RANKING order="13" place="13" resultid="1325" />
                    <RANKING order="14" place="14" resultid="1898" />
                    <RANKING order="15" place="-1" resultid="1927" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1143" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1494" />
                    <RANKING order="2" place="2" resultid="2183" />
                    <RANKING order="3" place="3" resultid="1247" />
                    <RANKING order="4" place="4" resultid="1904" />
                    <RANKING order="5" place="5" resultid="1336" />
                    <RANKING order="6" place="6" resultid="1386" />
                    <RANKING order="7" place="7" resultid="2131" />
                    <RANKING order="8" place="8" resultid="2142" />
                    <RANKING order="9" place="9" resultid="2068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1144" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2064" />
                    <RANKING order="2" place="2" resultid="2019" />
                    <RANKING order="3" place="3" resultid="1418" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1534" />
                    <RANKING order="2" place="2" resultid="2102" />
                    <RANKING order="3" place="3" resultid="1251" />
                    <RANKING order="4" place="4" resultid="1924" />
                    <RANKING order="5" place="-1" resultid="1400" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1146" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1287" />
                    <RANKING order="2" place="2" resultid="2110" />
                    <RANKING order="3" place="3" resultid="1881" />
                    <RANKING order="4" place="4" resultid="2029" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1822" />
                    <RANKING order="2" place="2" resultid="2014" />
                    <RANKING order="3" place="3" resultid="2039" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2296" daytime="16:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2297" daytime="16:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2298" daytime="16:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2299" daytime="16:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2300" daytime="16:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2301" daytime="16:52" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2302" daytime="16:54" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1148" daytime="16:58" gender="M" number="12" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1149" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1762" />
                    <RANKING order="2" place="2" resultid="1734" />
                    <RANKING order="3" place="3" resultid="1680" />
                    <RANKING order="4" place="4" resultid="2180" />
                    <RANKING order="5" place="5" resultid="1690" />
                    <RANKING order="6" place="6" resultid="1460" />
                    <RANKING order="7" place="7" resultid="1751" />
                    <RANKING order="8" place="8" resultid="1322" />
                    <RANKING order="9" place="9" resultid="1798" />
                    <RANKING order="10" place="10" resultid="2150" />
                    <RANKING order="11" place="11" resultid="1269" />
                    <RANKING order="12" place="12" resultid="2214" />
                    <RANKING order="13" place="13" resultid="2191" />
                    <RANKING order="14" place="14" resultid="2079" />
                    <RANKING order="15" place="15" resultid="1395" />
                    <RANKING order="16" place="16" resultid="1371" />
                    <RANKING order="17" place="17" resultid="1706" />
                    <RANKING order="18" place="18" resultid="1328" />
                    <RANKING order="19" place="19" resultid="1478" />
                    <RANKING order="20" place="20" resultid="1937" />
                    <RANKING order="21" place="21" resultid="2056" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1815" />
                    <RANKING order="2" place="2" resultid="1756" />
                    <RANKING order="3" place="3" resultid="1628" />
                    <RANKING order="4" place="4" resultid="1649" />
                    <RANKING order="5" place="5" resultid="1633" />
                    <RANKING order="6" place="6" resultid="1597" />
                    <RANKING order="7" place="7" resultid="1670" />
                    <RANKING order="8" place="8" resultid="1638" />
                    <RANKING order="9" place="9" resultid="2154" />
                    <RANKING order="10" place="10" resultid="1660" />
                    <RANKING order="11" place="11" resultid="2203" />
                    <RANKING order="12" place="12" resultid="1602" />
                    <RANKING order="13" place="13" resultid="1391" />
                    <RANKING order="14" place="14" resultid="1436" />
                    <RANKING order="15" place="15" resultid="1967" />
                    <RANKING order="16" place="16" resultid="1444" />
                    <RANKING order="17" place="17" resultid="2084" />
                    <RANKING order="18" place="18" resultid="1932" />
                    <RANKING order="19" place="19" resultid="1464" />
                    <RANKING order="20" place="20" resultid="1412" />
                    <RANKING order="21" place="21" resultid="1439" />
                    <RANKING order="22" place="22" resultid="1971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1151" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1506" />
                    <RANKING order="2" place="2" resultid="1226" />
                    <RANKING order="3" place="3" resultid="1379" />
                    <RANKING order="4" place="4" resultid="1979" />
                    <RANKING order="5" place="5" resultid="2135" />
                    <RANKING order="6" place="6" resultid="1257" />
                    <RANKING order="7" place="7" resultid="1872" />
                    <RANKING order="8" place="8" resultid="1408" />
                    <RANKING order="9" place="9" resultid="1261" />
                    <RANKING order="10" place="10" resultid="2011" />
                    <RANKING order="11" place="11" resultid="2231" />
                    <RANKING order="12" place="12" resultid="1581" />
                    <RANKING order="13" place="13" resultid="1431" />
                    <RANKING order="14" place="14" resultid="2071" />
                    <RANKING order="15" place="15" resultid="1474" />
                    <RANKING order="16" place="-1" resultid="1566" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1152" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1835" />
                    <RANKING order="2" place="2" resultid="2128" />
                    <RANKING order="3" place="3" resultid="1801" />
                    <RANKING order="4" place="4" resultid="2113" />
                    <RANKING order="5" place="5" resultid="1423" />
                    <RANKING order="6" place="6" resultid="1481" />
                    <RANKING order="7" place="7" resultid="2095" />
                    <RANKING order="8" place="8" resultid="1415" />
                    <RANKING order="9" place="9" resultid="1876" />
                    <RANKING order="10" place="10" resultid="1468" />
                    <RANKING order="11" place="11" resultid="1310" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1537" />
                    <RANKING order="2" place="2" resultid="2106" />
                    <RANKING order="3" place="3" resultid="2060" />
                    <RANKING order="4" place="4" resultid="1956" />
                    <RANKING order="5" place="5" resultid="2245" />
                    <RANKING order="6" place="6" resultid="1909" />
                    <RANKING order="7" place="7" resultid="2234" />
                    <RANKING order="8" place="8" resultid="2074" />
                    <RANKING order="9" place="9" resultid="1914" />
                    <RANKING order="10" place="-1" resultid="2090" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1154" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1848" />
                    <RANKING order="2" place="2" resultid="2138" />
                    <RANKING order="3" place="3" resultid="1342" />
                    <RANKING order="4" place="3" resultid="1858" />
                    <RANKING order="5" place="5" resultid="1674" />
                    <RANKING order="6" place="6" resultid="2002" />
                    <RANKING order="7" place="7" resultid="1353" />
                    <RANKING order="8" place="8" resultid="1947" />
                    <RANKING order="9" place="9" resultid="1265" />
                    <RANKING order="10" place="10" resultid="1453" />
                    <RANKING order="11" place="11" resultid="1471" />
                    <RANKING order="12" place="12" resultid="1884" />
                    <RANKING order="13" place="13" resultid="1944" />
                    <RANKING order="14" place="14" resultid="1276" />
                    <RANKING order="15" place="15" resultid="1545" />
                    <RANKING order="16" place="16" resultid="2034" />
                    <RANKING order="17" place="17" resultid="1283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1155" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1592" />
                    <RANKING order="2" place="2" resultid="1810" />
                    <RANKING order="3" place="3" resultid="1349" />
                    <RANKING order="4" place="4" resultid="1238" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2303" daytime="16:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2304" daytime="17:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2305" daytime="17:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2306" daytime="17:06" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2307" daytime="17:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2308" daytime="17:12" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2309" daytime="17:14" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="2310" daytime="17:16" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="2311" daytime="17:18" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="2312" daytime="17:20" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="2313" daytime="17:22" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="2314" daytime="17:24" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="2315" daytime="17:26" number="13" order="13" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1156" daytime="17:28" gender="F" number="13" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1157" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1780" />
                    <RANKING order="2" place="2" resultid="1721" />
                    <RANKING order="3" place="3" resultid="1699" />
                    <RANKING order="4" place="4" resultid="1832" />
                    <RANKING order="5" place="5" resultid="1711" />
                    <RANKING order="6" place="6" resultid="2187" />
                    <RANKING order="7" place="7" resultid="1919" />
                    <RANKING order="8" place="8" resultid="1319" />
                    <RANKING order="9" place="9" resultid="2217" />
                    <RANKING order="10" place="-1" resultid="2146" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2195" />
                    <RANKING order="2" place="2" resultid="1527" />
                    <RANKING order="3" place="3" resultid="1975" />
                    <RANKING order="4" place="4" resultid="2199" />
                    <RANKING order="5" place="5" resultid="1805" />
                    <RANKING order="6" place="6" resultid="1867" />
                    <RANKING order="7" place="7" resultid="1766" />
                    <RANKING order="8" place="8" resultid="1272" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1569" />
                    <RANKING order="2" place="2" resultid="1382" />
                    <RANKING order="3" place="3" resultid="1572" />
                    <RANKING order="4" place="4" resultid="1254" />
                    <RANKING order="5" place="5" resultid="1448" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1160" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1485" />
                    <RANKING order="2" place="2" resultid="1775" />
                    <RANKING order="3" place="3" resultid="1297" />
                    <RANKING order="4" place="4" resultid="2116" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1161" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1516" />
                    <RANKING order="2" place="2" resultid="1300" />
                    <RANKING order="3" place="-1" resultid="1399" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1162" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1242" />
                    <RANKING order="2" place="2" resultid="1880" />
                    <RANKING order="3" place="-1" resultid="1844" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1163" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2316" daytime="17:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2317" daytime="17:34" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2318" daytime="17:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2319" daytime="17:44" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2320" daytime="17:48" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1164" daytime="17:52" gender="M" number="14" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1165" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1689" />
                    <RANKING order="2" place="2" resultid="1733" />
                    <RANKING order="3" place="3" resultid="1750" />
                    <RANKING order="4" place="4" resultid="1789" />
                    <RANKING order="5" place="5" resultid="2158" />
                    <RANKING order="6" place="6" resultid="2162" />
                    <RANKING order="7" place="7" resultid="1705" />
                    <RANKING order="8" place="8" resultid="1394" />
                    <RANKING order="9" place="9" resultid="2221" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1648" />
                    <RANKING order="2" place="2" resultid="1596" />
                    <RANKING order="3" place="3" resultid="2166" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1232" />
                    <RANKING order="2" place="2" resultid="1978" />
                    <RANKING order="3" place="3" resultid="1575" />
                    <RANKING order="4" place="4" resultid="1367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1168" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1512" />
                    <RANKING order="2" place="2" resultid="1792" />
                    <RANKING order="3" place="3" resultid="1783" />
                    <RANKING order="4" place="4" resultid="1993" />
                    <RANKING order="5" place="5" resultid="1467" />
                    <RANKING order="6" place="-1" resultid="1557" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1541" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1170" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1498" />
                    <RANKING order="2" place="2" resultid="2173" />
                    <RANKING order="3" place="3" resultid="1943" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1171" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1235" />
                    <RANKING order="2" place="2" resultid="1345" />
                    <RANKING order="3" place="3" resultid="1360" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2321" daytime="17:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2322" daytime="17:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2323" daytime="18:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2324" daytime="18:06" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1172" daytime="18:12" gender="F" number="15" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1173" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1744" />
                    <RANKING order="2" place="2" resultid="1727" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1174" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1655" />
                    <RANKING order="2" place="2" resultid="1643" />
                    <RANKING order="3" place="3" resultid="1617" />
                    <RANKING order="4" place="4" resultid="2170" />
                    <RANKING order="5" place="5" resultid="1665" />
                    <RANKING order="6" place="6" resultid="1997" />
                    <RANKING order="7" place="7" resultid="1974" />
                    <RANKING order="8" place="8" resultid="1290" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1522" />
                    <RANKING order="2" place="2" resultid="2125" />
                    <RANKING order="3" place="3" resultid="1891" />
                    <RANKING order="4" place="-1" resultid="1488" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1176" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2018" />
                    <RANKING order="2" place="2" resultid="1952" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1177" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1533" />
                    <RANKING order="2" place="2" resultid="1923" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1178" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1179" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2325" daytime="18:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2326" daytime="18:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2327" daytime="18:38" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1180" daytime="18:50" gender="M" number="16" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1181" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1685" />
                    <RANKING order="2" place="2" resultid="1679" />
                    <RANKING order="3" place="3" resultid="1695" />
                    <RANKING order="4" place="4" resultid="1732" />
                    <RANKING order="5" place="5" resultid="1716" />
                    <RANKING order="6" place="6" resultid="1797" />
                    <RANKING order="7" place="7" resultid="1739" />
                    <RANKING order="8" place="8" resultid="2190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1627" />
                    <RANKING order="2" place="2" resultid="1637" />
                    <RANKING order="3" place="3" resultid="1669" />
                    <RANKING order="4" place="4" resultid="1755" />
                    <RANKING order="5" place="5" resultid="1966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1183" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1962" />
                    <RANKING order="2" place="2" resultid="1530" />
                    <RANKING order="3" place="3" resultid="1585" />
                    <RANKING order="4" place="4" resultid="1260" />
                    <RANKING order="5" place="5" resultid="1505" />
                    <RANKING order="6" place="6" resultid="1563" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1184" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1861" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2059" />
                    <RANKING order="2" place="2" resultid="2021" />
                    <RANKING order="3" place="3" resultid="2089" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1186" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1946" />
                    <RANKING order="2" place="2" resultid="1987" />
                    <RANKING order="3" place="3" resultid="1544" />
                    <RANKING order="4" place="4" resultid="2033" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1187" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2007" />
                    <RANKING order="2" place="2" resultid="1357" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2328" daytime="18:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2329" daytime="19:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2330" daytime="19:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2331" daytime="19:32" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1188" daytime="19:44" gender="F" number="17" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1189" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1743" />
                    <RANKING order="2" place="2" resultid="1771" />
                    <RANKING order="3" place="3" resultid="1726" />
                    <RANKING order="4" place="4" resultid="1279" />
                    <RANKING order="5" place="5" resultid="1827" />
                    <RANKING order="6" place="6" resultid="1983" />
                    <RANKING order="7" place="-1" resultid="1427" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1190" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1611" />
                    <RANKING order="2" place="2" resultid="1606" />
                    <RANKING order="3" place="3" resultid="1306" />
                    <RANKING order="4" place="4" resultid="1622" />
                    <RANKING order="5" place="5" resultid="1866" />
                    <RANKING order="6" place="6" resultid="1642" />
                    <RANKING order="7" place="7" resultid="2198" />
                    <RANKING order="8" place="8" resultid="2238" />
                    <RANKING order="9" place="9" resultid="2242" />
                    <RANKING order="10" place="10" resultid="2044" />
                    <RANKING order="11" place="-1" resultid="1616" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1191" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1335" />
                    <RANKING order="2" place="2" resultid="1246" />
                    <RANKING order="3" place="3" resultid="1578" />
                    <RANKING order="4" place="4" resultid="2067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1192" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1951" />
                    <RANKING order="2" place="2" resultid="2053" />
                    <RANKING order="3" place="-1" resultid="1838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1193" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1250" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1194" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1195" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2332" daytime="19:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2333" daytime="19:50" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2334" daytime="19:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2335" daytime="20:00" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1196" daytime="20:04" gender="M" number="18" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1197" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1761" />
                    <RANKING order="2" place="2" resultid="1694" />
                    <RANKING order="3" place="3" resultid="1936" />
                    <RANKING order="4" place="-1" resultid="2149" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1814" />
                    <RANKING order="2" place="2" resultid="1632" />
                    <RANKING order="3" place="3" resultid="1601" />
                    <RANKING order="4" place="4" resultid="2210" />
                    <RANKING order="5" place="5" resultid="1931" />
                    <RANKING order="6" place="6" resultid="1463" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1199" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1340" />
                    <RANKING order="2" place="2" resultid="1854" />
                    <RANKING order="3" place="3" resultid="1225" />
                    <RANKING order="4" place="4" resultid="1977" />
                    <RANKING order="5" place="5" resultid="2206" />
                    <RANKING order="6" place="6" resultid="2122" />
                    <RANKING order="7" place="7" resultid="1584" />
                    <RANKING order="8" place="8" resultid="1961" />
                    <RANKING order="9" place="9" resultid="1407" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1200" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1502" />
                    <RANKING order="2" place="2" resultid="1588" />
                    <RANKING order="3" place="3" resultid="1551" />
                    <RANKING order="4" place="4" resultid="1560" />
                    <RANKING order="5" place="5" resultid="1548" />
                    <RANKING order="6" place="6" resultid="1887" />
                    <RANKING order="7" place="7" resultid="1303" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1201" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1851" />
                    <RANKING order="2" place="2" resultid="1908" />
                    <RANKING order="3" place="-1" resultid="1913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1202" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1203" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2336" daytime="20:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2337" daytime="20:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2338" daytime="20:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2339" daytime="20:18" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1204" daytime="20:22" gender="F" number="19" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1205" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1779" />
                    <RANKING order="2" place="2" resultid="1831" />
                    <RANKING order="3" place="3" resultid="1918" />
                    <RANKING order="4" place="4" resultid="1826" />
                    <RANKING order="5" place="5" resultid="1894" />
                    <RANKING order="6" place="6" resultid="1710" />
                    <RANKING order="7" place="7" resultid="1315" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1206" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1654" />
                    <RANKING order="2" place="2" resultid="2169" />
                    <RANKING order="3" place="3" resultid="2227" />
                    <RANKING order="4" place="4" resultid="1526" />
                    <RANKING order="5" place="5" resultid="1664" />
                    <RANKING order="6" place="6" resultid="2048" />
                    <RANKING order="7" place="7" resultid="2043" />
                    <RANKING order="8" place="-1" resultid="1610" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2099" />
                    <RANKING order="2" place="2" resultid="1903" />
                    <RANKING order="3" place="3" resultid="2066" />
                    <RANKING order="4" place="4" resultid="1890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1208" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1491" />
                    <RANKING order="2" place="2" resultid="1294" />
                    <RANKING order="3" place="3" resultid="1417" />
                    <RANKING order="4" place="4" resultid="1313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1209" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1210" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2109" />
                    <RANKING order="2" place="2" resultid="1241" />
                    <RANKING order="3" place="3" resultid="1989" />
                    <RANKING order="4" place="4" resultid="2028" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2038" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2340" daytime="20:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2341" daytime="20:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2342" daytime="20:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2343" daytime="20:30" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1212" daytime="20:34" gender="M" number="20" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1213" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2179" />
                    <RANKING order="2" place="2" resultid="1715" />
                    <RANKING order="3" place="3" resultid="1684" />
                    <RANKING order="4" place="4" resultid="1760" />
                    <RANKING order="5" place="5" resultid="1678" />
                    <RANKING order="6" place="6" resultid="2157" />
                    <RANKING order="7" place="7" resultid="1788" />
                    <RANKING order="8" place="8" resultid="1738" />
                    <RANKING order="9" place="-1" resultid="2213" />
                    <RANKING order="10" place="-1" resultid="2055" />
                    <RANKING order="11" place="-1" resultid="1370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1375" />
                    <RANKING order="2" place="2" resultid="2153" />
                    <RANKING order="3" place="3" resultid="1647" />
                    <RANKING order="4" place="4" resultid="2202" />
                    <RANKING order="5" place="5" resultid="1659" />
                    <RANKING order="6" place="6" resultid="2083" />
                    <RANKING order="7" place="-1" resultid="2165" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1841" />
                    <RANKING order="2" place="2" resultid="1231" />
                    <RANKING order="3" place="3" resultid="2119" />
                    <RANKING order="4" place="4" resultid="1256" />
                    <RANKING order="5" place="5" resultid="1366" />
                    <RANKING order="6" place="6" resultid="1378" />
                    <RANKING order="7" place="7" resultid="1580" />
                    <RANKING order="8" place="8" resultid="2070" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1216" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1554" />
                    <RANKING order="2" place="2" resultid="1818" />
                    <RANKING order="3" place="3" resultid="1422" />
                    <RANKING order="4" place="4" resultid="2094" />
                    <RANKING order="5" place="-1" resultid="1509" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1217" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1540" />
                    <RANKING order="2" place="2" resultid="1955" />
                    <RANKING order="3" place="3" resultid="2105" />
                    <RANKING order="4" place="4" resultid="2088" />
                    <RANKING order="5" place="-1" resultid="1519" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1673" />
                    <RANKING order="2" place="2" resultid="1847" />
                    <RANKING order="3" place="3" resultid="2176" />
                    <RANKING order="4" place="4" resultid="1857" />
                    <RANKING order="5" place="5" resultid="2001" />
                    <RANKING order="6" place="6" resultid="1264" />
                    <RANKING order="7" place="7" resultid="1352" />
                    <RANKING order="8" place="8" resultid="1470" />
                    <RANKING order="9" place="9" resultid="1452" />
                    <RANKING order="10" place="-1" resultid="1883" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1591" />
                    <RANKING order="2" place="2" resultid="1363" />
                    <RANKING order="3" place="3" resultid="1809" />
                    <RANKING order="4" place="4" resultid="1344" />
                    <RANKING order="5" place="5" resultid="1348" />
                    <RANKING order="6" place="6" resultid="2006" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2344" daytime="20:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2345" daytime="20:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2346" daytime="20:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2347" daytime="20:42" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2348" daytime="20:44" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2349" daytime="20:46" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2350" daytime="20:48" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="1899" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Vinicius" lastname="Henrique Ramos" birthdate="2010-02-25" gender="M" nation="BRA" license="406916" athleteid="1928" externalid="406916">
              <RESULTS>
                <RESULT eventid="1116" points="189" reactiontime="+68" swimtime="00:01:29.88" resultid="1929" heatid="2277" lane="5" />
                <RESULT eventid="1084" points="241" swimtime="00:02:43.78" resultid="1930" heatid="2257" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="192" reactiontime="+64" swimtime="00:03:13.79" resultid="1931" heatid="2336" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="256" swimtime="00:01:13.74" resultid="1932" heatid="2305" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Clara Cominato" birthdate="2010-04-09" gender="F" nation="BRA" license="406915" athleteid="1925" externalid="406915">
              <RESULTS>
                <RESULT eventid="1108" points="176" reactiontime="+75" swimtime="00:01:42.18" resultid="1926" heatid="2272" lane="7" />
                <RESULT eventid="1140" status="DSQ" swimtime="00:01:36.13" resultid="1927" heatid="2296" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Ferreira Rais" birthdate="2007-07-04" gender="M" nation="BRA" license="398656" swrid="5697227" athleteid="1910" externalid="398656">
              <RESULTS>
                <RESULT eventid="1116" points="220" reactiontime="+66" swimtime="00:01:25.43" resultid="1911" heatid="2278" lane="5" />
                <RESULT eventid="1084" points="253" swimtime="00:02:41.22" resultid="1912" heatid="2260" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" reactiontime="+82" status="DSQ" swimtime="00:03:12.18" resultid="1913" heatid="2336" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="343" swimtime="00:01:06.94" resultid="1914" heatid="2307" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jennifer" lastname="De Abreu" birthdate="2009-11-07" gender="F" nation="BRA" license="356212" swrid="5600144" athleteid="1900" externalid="356212">
              <RESULTS>
                <RESULT eventid="1124" points="384" swimtime="00:01:28.23" resultid="1901" heatid="2283" lane="4" />
                <RESULT eventid="1076" points="471" swimtime="00:02:24.99" resultid="1902" heatid="2255" lane="3" entrytime="00:02:23.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="373" swimtime="00:01:17.06" resultid="1903" heatid="2341" lane="2" />
                <RESULT eventid="1140" points="498" swimtime="00:01:05.23" resultid="1904" heatid="2301" lane="4" entrytime="00:01:05.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rodrigo" lastname="Zanatta Duda" birthdate="2011-09-12" gender="M" nation="BRA" license="406917" swrid="5717307" athleteid="1933" externalid="406917">
              <RESULTS>
                <RESULT eventid="1132" status="DSQ" swimtime="00:00:00.00" resultid="1934" heatid="2288" lane="3" />
                <RESULT eventid="1116" points="191" reactiontime="+80" swimtime="00:01:29.57" resultid="1935" heatid="2278" lane="6" />
                <RESULT eventid="1196" points="202" reactiontime="+73" swimtime="00:03:10.66" resultid="1936" heatid="2337" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="143" swimtime="00:01:29.58" resultid="1937" heatid="2305" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Ribeiro Melo" birthdate="2011-07-01" gender="F" nation="BRA" license="390923" swrid="5602577" athleteid="1915" externalid="390923">
              <RESULTS>
                <RESULT eventid="1108" points="292" reactiontime="+72" swimtime="00:01:26.41" resultid="1916" heatid="2271" lane="2" />
                <RESULT eventid="1076" points="393" swimtime="00:02:34.05" resultid="1917" heatid="2252" lane="7" entrytime="00:02:50.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="186" swimtime="00:01:37.04" resultid="1918" heatid="2341" lane="4" />
                <RESULT eventid="1156" points="267" swimtime="00:03:33.54" resultid="1919" heatid="2316" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aline" lastname="Hirano" birthdate="2007-11-13" gender="F" nation="BRA" license="358898" swrid="5622283" athleteid="1920" externalid="358898">
              <RESULTS>
                <RESULT eventid="1108" points="329" reactiontime="+70" swimtime="00:01:22.99" resultid="1921" heatid="2274" lane="6" entrytime="00:01:22.87" entrycourse="LCM" />
                <RESULT eventid="1076" points="399" swimtime="00:02:33.20" resultid="1922" heatid="2253" lane="6" entrytime="00:02:34.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="389" swimtime="00:11:03.62" resultid="1923" heatid="2326" lane="4" entrytime="00:11:26.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.85" />
                    <SPLIT distance="200" swimtime="00:02:42.42" />
                    <SPLIT distance="300" swimtime="00:04:05.50" />
                    <SPLIT distance="400" swimtime="00:05:28.77" />
                    <SPLIT distance="500" swimtime="00:06:53.07" />
                    <SPLIT distance="600" swimtime="00:08:18.41" />
                    <SPLIT distance="700" swimtime="00:09:44.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="413" swimtime="00:01:09.39" resultid="1924" heatid="2300" lane="1" entrytime="00:01:10.26" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Guilherme Ballatka" birthdate="2007-06-24" gender="M" nation="BRA" license="398616" swrid="5697228" athleteid="1905" externalid="398616">
              <RESULTS>
                <RESULT eventid="1116" points="342" reactiontime="+84" swimtime="00:01:13.76" resultid="1906" heatid="2277" lane="2" />
                <RESULT eventid="1084" points="297" swimtime="00:02:32.85" resultid="1907" heatid="2258" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="311" reactiontime="+83" swimtime="00:02:45.06" resultid="1908" heatid="2336" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="368" swimtime="00:01:05.35" resultid="1909" heatid="2305" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Camillo Sabim" birthdate="2010-08-02" gender="F" nation="BRA" license="406931" athleteid="1938" externalid="406931">
              <RESULTS>
                <RESULT eventid="1108" points="199" reactiontime="+74" swimtime="00:01:38.08" resultid="1939" heatid="2272" lane="2" />
                <RESULT eventid="1140" points="224" swimtime="00:01:25.08" resultid="1940" heatid="2297" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11303" nation="BRA" region="PR" clubid="1332" swrid="93760" name="Associação De Talentos Da Natação" shortname="Atn/Curitiba">
          <ATHLETES>
            <ATHLETE firstname="Jhon" lastname="Caleb Dos Santos" birthdate="2010-03-02" gender="M" nation="BRA" license="359020" swrid="5588574" athleteid="1372" externalid="359020">
              <RESULTS>
                <RESULT eventid="1132" points="376" swimtime="00:01:18.75" resultid="1373" heatid="2294" lane="6" entrytime="00:01:18.40" entrycourse="LCM" />
                <RESULT eventid="1068" points="378" swimtime="00:05:35.27" resultid="1374" heatid="2248" lane="6" entrytime="00:05:24.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.70" />
                    <SPLIT distance="200" swimtime="00:02:33.14" />
                    <SPLIT distance="300" swimtime="00:04:15.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="426" swimtime="00:01:05.68" resultid="1375" heatid="2348" lane="5" entrytime="00:01:06.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelo" lastname="Correia Bonfim" birthdate="2009-06-21" gender="M" nation="BRA" license="391663" swrid="5622271" athleteid="1404" externalid="391663">
              <RESULTS>
                <RESULT eventid="1132" points="264" swimtime="00:01:28.62" resultid="1405" heatid="2292" lane="4" entrytime="00:01:32.05" entrycourse="LCM" />
                <RESULT eventid="1084" points="352" swimtime="00:02:24.46" resultid="1406" heatid="2259" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="312" reactiontime="+69" swimtime="00:02:44.91" resultid="1407" heatid="2337" lane="6" entrytime="00:02:48.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="403" swimtime="00:01:03.44" resultid="1408" heatid="2309" lane="8" entrytime="00:01:11.10" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Iglesias Prado" birthdate="2010-06-15" gender="M" nation="BRA" license="408052" athleteid="1440" externalid="408052">
              <RESULTS>
                <RESULT eventid="1132" points="166" swimtime="00:01:43.32" resultid="1441" heatid="2289" lane="1" />
                <RESULT eventid="1116" points="161" reactiontime="+68" swimtime="00:01:34.71" resultid="1442" heatid="2279" lane="7" />
                <RESULT eventid="1084" points="230" swimtime="00:02:46.41" resultid="1443" heatid="2260" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="271" swimtime="00:01:12.35" resultid="1444" heatid="2303" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Faria Del Valle" birthdate="2009-08-28" gender="M" nation="BRA" license="376328" swrid="5600155" athleteid="1376" externalid="376328">
              <RESULTS>
                <RESULT eventid="1132" points="348" swimtime="00:01:20.86" resultid="1377" heatid="2290" lane="2" />
                <RESULT eventid="1212" points="304" swimtime="00:01:13.51" resultid="1378" heatid="2345" lane="1" />
                <RESULT eventid="1148" points="489" swimtime="00:00:59.47" resultid="1379" heatid="2313" lane="8" entrytime="00:01:00.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Angelo" lastname="De Queiroz Neto" birthdate="2003-10-31" gender="M" nation="BRA" license="342814" swrid="5600149" athleteid="1346" externalid="342814" level="AERC">
              <RESULTS>
                <RESULT eventid="1084" points="394" swimtime="00:02:19.06" resultid="1347" heatid="2265" lane="2" entrytime="00:02:15.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="379" swimtime="00:01:08.28" resultid="1348" heatid="2348" lane="6" entrytime="00:01:07.67" entrycourse="LCM" />
                <RESULT eventid="1148" points="444" swimtime="00:01:01.40" resultid="1349" heatid="2312" lane="4" entrytime="00:01:00.52" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Muller" birthdate="2009-10-10" gender="F" nation="BRA" license="376952" swrid="5600221" athleteid="1380" externalid="376952">
              <RESULTS>
                <RESULT eventid="1124" points="425" swimtime="00:01:25.26" resultid="1381" heatid="2287" lane="7" entrytime="00:01:21.69" entrycourse="LCM" />
                <RESULT eventid="1156" points="418" swimtime="00:03:03.89" resultid="1382" heatid="2320" lane="1" entrytime="00:02:59.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Kerppers Kreia" birthdate="2006-12-01" gender="M" nation="BRA" license="366815" swrid="5600195" athleteid="1350" externalid="366815">
              <RESULTS>
                <RESULT eventid="1084" points="462" swimtime="00:02:11.88" resultid="1351" heatid="2265" lane="4" entrytime="00:02:13.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="314" swimtime="00:01:12.73" resultid="1352" heatid="2345" lane="6" />
                <RESULT eventid="1148" points="493" swimtime="00:00:59.28" resultid="1353" heatid="2313" lane="3" entrytime="00:00:59.59" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Bortoleto" birthdate="2008-09-05" gender="M" nation="BRA" license="406709" swrid="5717249" athleteid="1419" externalid="406709">
              <RESULTS>
                <RESULT eventid="1116" reactiontime="+47" status="DSQ" swimtime="00:01:19.99" resultid="1420" heatid="2279" lane="6" />
                <RESULT eventid="1100" points="180" swimtime="00:03:15.16" resultid="1421" heatid="2269" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="310" swimtime="00:01:13.02" resultid="1422" heatid="2344" lane="5" />
                <RESULT eventid="1148" points="383" swimtime="00:01:04.50" resultid="1423" heatid="2304" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Fonseca Vendramin" birthdate="2008-09-28" gender="F" nation="BRA" license="393918" swrid="5622282" athleteid="1416" externalid="393918">
              <RESULTS>
                <RESULT eventid="1204" points="275" swimtime="00:01:25.31" resultid="1417" heatid="2341" lane="6" />
                <RESULT eventid="1140" points="369" swimtime="00:01:12.04" resultid="1418" heatid="2299" lane="8" entrytime="00:01:15.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Inacio Carneiro" birthdate="2009-09-09" gender="M" nation="BRA" license="408023" athleteid="1429" externalid="408023">
              <RESULTS>
                <RESULT eventid="1084" points="189" swimtime="00:02:57.66" resultid="1430" heatid="2261" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="252" swimtime="00:01:14.15" resultid="1431" heatid="2306" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mauricio" lastname="Furtado Niwa" birthdate="1978-05-30" gender="M" nation="BRA" license="398757" swrid="5653291" athleteid="1361" externalid="398757">
              <RESULTS>
                <RESULT eventid="1100" points="356" swimtime="00:02:35.57" resultid="1362" heatid="2270" lane="6" entrytime="00:02:31.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="486" swimtime="00:01:02.87" resultid="1363" heatid="2349" lane="5" entrytime="00:01:01.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Riccieri" lastname="Rodrigues Muzolon" birthdate="2010-11-08" gender="M" nation="BRA" license="385439" swrid="5588887" athleteid="1387" externalid="385439">
              <RESULTS>
                <RESULT eventid="1132" points="250" swimtime="00:01:30.27" resultid="1388" heatid="2292" lane="3" entrytime="00:01:33.11" entrycourse="LCM" />
                <RESULT eventid="1116" points="248" reactiontime="+78" swimtime="00:01:22.03" resultid="1389" heatid="2280" lane="2" entrytime="00:01:22.21" entrycourse="LCM" />
                <RESULT eventid="1084" points="254" swimtime="00:02:41.05" resultid="1390" heatid="2262" lane="7" entrytime="00:02:40.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="312" swimtime="00:01:09.08" resultid="1391" heatid="2308" lane="6" entrytime="00:01:11.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Kerniski Demantova" birthdate="1982-05-25" gender="M" nation="BRA" license="398222" swrid="5653293" athleteid="1354" externalid="398222">
              <RESULTS>
                <RESULT eventid="1132" points="326" swimtime="00:01:22.61" resultid="1355" heatid="2289" lane="3" />
                <RESULT eventid="1084" points="373" swimtime="00:02:21.69" resultid="1356" heatid="2264" lane="2" entrytime="00:02:20.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="365" swimtime="00:10:32.52" resultid="1357" heatid="2330" lane="6" entrytime="00:10:29.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.64" />
                    <SPLIT distance="200" swimtime="00:02:33.47" />
                    <SPLIT distance="300" swimtime="00:03:54.03" />
                    <SPLIT distance="400" swimtime="00:05:14.06" />
                    <SPLIT distance="500" swimtime="00:06:34.20" />
                    <SPLIT distance="600" swimtime="00:07:54.75" />
                    <SPLIT distance="700" swimtime="00:09:15.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="James" lastname="Roberto Zoschke" birthdate="1976-02-08" gender="M" nation="BRA" license="312251" swrid="5688617" athleteid="1358" externalid="312251">
              <RESULTS>
                <RESULT eventid="1132" points="450" swimtime="00:01:14.18" resultid="1359" heatid="2291" lane="5" />
                <RESULT eventid="1164" points="401" swimtime="00:02:50.10" resultid="1360" heatid="2322" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Navarro Silva" birthdate="2011-01-10" gender="F" nation="BRA" license="406711" swrid="5717284" athleteid="1424" externalid="406711">
              <RESULTS>
                <RESULT eventid="1108" points="261" reactiontime="+83" swimtime="00:01:29.62" resultid="1425" heatid="2271" lane="3" />
                <RESULT eventid="1076" points="272" swimtime="00:02:53.97" resultid="1426" heatid="2250" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" status="DNS" swimtime="00:00:00.00" resultid="1427" heatid="2333" lane="7" />
                <RESULT eventid="1140" status="DNS" swimtime="00:00:00.00" resultid="1428" heatid="2296" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Arthur Ribeiro" birthdate="2010-02-05" gender="M" nation="BRA" license="408025" athleteid="1437" externalid="408025">
              <RESULTS>
                <RESULT eventid="1132" points="208" swimtime="00:01:35.86" resultid="1438" heatid="2289" lane="2" />
                <RESULT eventid="1148" points="204" swimtime="00:01:19.52" resultid="1439" heatid="2304" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabiana" lastname="Zaleski Dallazem" birthdate="2009-05-16" gender="F" nation="BRA" license="344287" swrid="5600279" athleteid="1333" externalid="344287" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1108" points="479" reactiontime="+59" swimtime="00:01:13.23" resultid="1334" heatid="2276" lane="6" entrytime="00:01:10.23" entrycourse="LCM" />
                <RESULT eventid="1188" points="470" reactiontime="+64" swimtime="00:02:38.35" resultid="1335" heatid="2335" lane="5" entrytime="00:02:38.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="489" swimtime="00:01:05.60" resultid="1336" heatid="2301" lane="3" entrytime="00:01:06.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Zaleski Dallazem" birthdate="2009-05-16" gender="M" nation="BRA" license="344286" swrid="5600280" athleteid="1364" externalid="344286" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1132" points="396" swimtime="00:01:17.44" resultid="1365" heatid="2293" lane="4" entrytime="00:01:22.82" entrycourse="LCM" />
                <RESULT eventid="1212" points="320" swimtime="00:01:12.24" resultid="1366" heatid="2346" lane="3" />
                <RESULT eventid="1164" points="381" swimtime="00:02:53.04" resultid="1367" heatid="2323" lane="2" entrytime="00:03:01.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcos" lastname="Demchuk" birthdate="2011-06-15" gender="M" nation="BRA" license="388540" swrid="5602530" athleteid="1392" externalid="388540">
              <RESULTS>
                <RESULT eventid="1132" points="194" swimtime="00:01:38.13" resultid="1393" heatid="2291" lane="4" entrytime="00:01:54.58" entrycourse="LCM" />
                <RESULT eventid="1164" points="170" swimtime="00:03:46.24" resultid="1394" heatid="2321" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="218" swimtime="00:01:17.76" resultid="1395" heatid="2307" lane="2" entrytime="00:01:21.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Neves Vianna" birthdate="2007-12-30" gender="F" nation="BRA" license="391106" swrid="5600223" athleteid="1401" externalid="391106">
              <RESULTS>
                <RESULT eventid="1108" points="206" reactiontime="+61" swimtime="00:01:37.06" resultid="1402" heatid="2273" lane="8" entrytime="00:01:36.54" entrycourse="LCM" />
                <RESULT eventid="1076" points="224" swimtime="00:03:05.59" resultid="1403" heatid="2251" lane="3" entrytime="00:03:00.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Sofia Silva" birthdate="2007-05-28" gender="F" nation="BRA" license="390921" swrid="5600260" athleteid="1396" externalid="390921">
              <RESULTS>
                <RESULT eventid="1124" points="189" swimtime="00:01:51.65" resultid="1397" heatid="2284" lane="7" entrytime="00:01:57.68" entrycourse="LCM" />
                <RESULT eventid="1076" points="213" swimtime="00:03:08.82" resultid="1398" heatid="2250" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="1399" heatid="2317" lane="5" entrytime="00:04:15.91" entrycourse="LCM" />
                <RESULT eventid="1140" status="DNS" swimtime="00:00:00.00" resultid="1400" heatid="2297" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Castellano Purkot" birthdate="2010-01-25" gender="M" nation="BRA" license="392484" swrid="5622268" athleteid="1409" externalid="392484">
              <RESULTS>
                <RESULT eventid="1116" points="186" reactiontime="+82" swimtime="00:01:30.27" resultid="1410" heatid="2277" lane="4" />
                <RESULT eventid="1084" points="184" swimtime="00:02:59.24" resultid="1411" heatid="2258" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="226" swimtime="00:01:16.90" resultid="1412" heatid="2310" lane="8" entrytime="00:01:08.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Dallastra" birthdate="2010-08-21" gender="M" nation="BRA" license="408024" athleteid="1432" externalid="408024">
              <RESULTS>
                <RESULT eventid="1132" status="DSQ" swimtime="00:01:46.41" resultid="1433" heatid="2291" lane="3" />
                <RESULT eventid="1116" points="145" reactiontime="+75" swimtime="00:01:38.16" resultid="1434" heatid="2278" lane="3" />
                <RESULT eventid="1084" points="291" swimtime="00:02:33.88" resultid="1435" heatid="2260" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="281" swimtime="00:01:11.52" resultid="1436" heatid="2306" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Yuji Yamazato" birthdate="2008-10-01" gender="M" nation="BRA" license="392664" swrid="5622313" athleteid="1413" externalid="392664">
              <RESULTS>
                <RESULT eventid="1084" points="289" swimtime="00:02:34.20" resultid="1414" heatid="2262" lane="3" entrytime="00:02:36.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="346" swimtime="00:01:06.72" resultid="1415" heatid="2310" lane="6" entrytime="00:01:06.10" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Garcia Fraga" birthdate="2003-10-07" gender="M" nation="BRA" license="283467" swrid="5717265" athleteid="1343" externalid="283467" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1212" points="441" swimtime="00:01:04.95" resultid="1344" heatid="2345" lane="7" />
                <RESULT eventid="1164" points="440" swimtime="00:02:44.88" resultid="1345" heatid="2321" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Garcia De Fraga" birthdate="2009-03-24" gender="M" nation="BRA" license="342147" swrid="5600172" athleteid="1337" externalid="342147" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1116" points="577" reactiontime="+60" swimtime="00:01:01.95" resultid="1338" heatid="2282" lane="6" entrytime="00:01:02.29" entrycourse="LCM" />
                <RESULT eventid="1068" points="517" swimtime="00:05:02.02" resultid="1339" heatid="2248" lane="3" entrytime="00:05:08.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.90" />
                    <SPLIT distance="200" swimtime="00:02:21.91" />
                    <SPLIT distance="300" swimtime="00:03:51.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="511" reactiontime="+61" swimtime="00:02:19.92" resultid="1340" heatid="2339" lane="5" entrytime="00:02:17.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Camila" lastname="Duarte De Almeida" birthdate="2009-11-26" gender="F" nation="BRA" license="378819" swrid="5600152" athleteid="1383" externalid="378819">
              <RESULTS>
                <RESULT eventid="1108" points="334" reactiontime="+105" swimtime="00:01:22.57" resultid="1384" heatid="2273" lane="4" entrytime="00:01:27.48" entrycourse="LCM" />
                <RESULT eventid="1076" points="390" swimtime="00:02:34.36" resultid="1385" heatid="2253" lane="2" entrytime="00:02:35.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="442" swimtime="00:01:07.85" resultid="1386" heatid="2300" lane="5" entrytime="00:01:08.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Ocanha" birthdate="2005-06-21" gender="M" nation="BRA" license="313769" swrid="5600231" athleteid="1341" externalid="313769" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1148" points="613" swimtime="00:00:55.15" resultid="1342" heatid="2314" lane="4" entrytime="00:00:54.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Freitas Szucs" birthdate="2011-10-02" gender="M" nation="BRA" license="377272" swrid="5588708" athleteid="1368" externalid="377272">
              <RESULTS>
                <RESULT eventid="1084" points="188" swimtime="00:02:58.01" resultid="1369" heatid="2261" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" status="DSQ" swimtime="00:02:04.39" resultid="1370" heatid="2344" lane="3" />
                <RESULT eventid="1148" points="201" swimtime="00:01:19.98" resultid="1371" heatid="2307" lane="5" entrytime="00:01:18.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13038" nation="BRA" region="PR" clubid="1284" swrid="93759" name="Associação De Pais E Atletas De Natação Ws/Crb" shortname="Apan/Ws">
          <ATHLETES>
            <ATHLETE firstname="Heloisa" lastname="Daniele Silva" birthdate="2010-07-06" gender="F" nation="BRA" license="359593" swrid="5588628" athleteid="1304" externalid="359593" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1108" points="403" swimtime="00:01:17.58" resultid="1305" heatid="2275" lane="1" entrytime="00:01:21.30" entrycourse="LCM" />
                <RESULT eventid="1188" points="352" reactiontime="+72" swimtime="00:02:54.36" resultid="1306" heatid="2334" lane="6" entrytime="00:02:59.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="394" swimtime="00:01:10.50" resultid="1307" heatid="2300" lane="7" entrytime="00:01:09.94" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Zeclhynski Silva" birthdate="2006-09-14" gender="F" nation="BRA" license="330727" swrid="5600283" athleteid="1285" externalid="330727" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1108" points="617" reactiontime="+69" swimtime="00:01:07.34" resultid="1286" heatid="2276" lane="4" entrytime="00:01:06.10" entrycourse="LCM" />
                <RESULT eventid="1140" points="585" swimtime="00:01:01.82" resultid="1287" heatid="2302" lane="5" entrytime="00:01:01.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Alexandre Azevedo" birthdate="2008-05-20" gender="M" nation="BRA" license="398694" swrid="5717240" athleteid="1308" externalid="398694">
              <RESULTS>
                <RESULT eventid="1132" points="181" swimtime="00:01:40.53" resultid="1309" heatid="2290" lane="3" />
                <RESULT eventid="1148" points="283" swimtime="00:01:11.37" resultid="1310" heatid="2304" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Rosa Silva" birthdate="2011-03-25" gender="F" nation="BRA" license="392120" swrid="5602579" athleteid="1317" externalid="392120">
              <RESULTS>
                <RESULT eventid="1124" points="184" swimtime="00:01:52.74" resultid="1318" heatid="2284" lane="1" />
                <RESULT eventid="1156" points="179" swimtime="00:04:03.77" resultid="1319" heatid="2316" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabelly" lastname="Mendonca Bello" birthdate="2008-04-15" gender="F" nation="BRA" license="376996" swrid="5600217" athleteid="1295" externalid="376996" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1124" points="370" swimtime="00:01:29.32" resultid="1296" heatid="2286" lane="8" entrytime="00:01:30.08" entrycourse="LCM" />
                <RESULT eventid="1156" points="360" swimtime="00:03:13.19" resultid="1297" heatid="2319" lane="1" entrytime="00:03:11.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Sieck" birthdate="2011-01-20" gender="F" nation="BRA" license="382234" swrid="5602584" athleteid="1314" externalid="382234">
              <RESULTS>
                <RESULT eventid="1204" points="128" swimtime="00:01:49.97" resultid="1315" heatid="2342" lane="2" entrytime="00:01:45.07" entrycourse="LCM" />
                <RESULT eventid="1140" points="199" swimtime="00:01:28.51" resultid="1316" heatid="2298" lane="1" entrytime="00:01:35.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Da Costa Riekes" birthdate="2008-06-19" gender="F" nation="BRA" license="331686" swrid="5600143" athleteid="1291" externalid="331686" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1108" points="403" reactiontime="+91" swimtime="00:01:17.56" resultid="1292" heatid="2275" lane="4" entrytime="00:01:16.33" entrycourse="LCM" />
                <RESULT eventid="1076" points="453" swimtime="00:02:26.89" resultid="1293" heatid="2255" lane="6" entrytime="00:02:24.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="368" swimtime="00:01:17.41" resultid="1294" heatid="2343" lane="2" entrytime="00:01:13.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonia" lastname="Adam  Fracaro" birthdate="2010-04-27" gender="F" nation="BRA" license="382212" swrid="5588512" athleteid="1288" externalid="382212">
              <RESULTS>
                <RESULT eventid="1076" points="304" swimtime="00:02:47.79" resultid="1289" heatid="2252" lane="2" entrytime="00:02:48.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="263" swimtime="00:12:35.94" resultid="1290" heatid="2326" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.21" />
                    <SPLIT distance="200" swimtime="00:02:54.63" />
                    <SPLIT distance="300" swimtime="00:04:32.27" />
                    <SPLIT distance="400" swimtime="00:06:09.49" />
                    <SPLIT distance="500" swimtime="00:07:47.16" />
                    <SPLIT distance="600" swimtime="00:09:26.63" />
                    <SPLIT distance="700" swimtime="00:11:04.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Zanchetta Silva" birthdate="2010-08-05" gender="F" nation="BRA" license="406865" swrid="5717308" athleteid="1323" externalid="406865">
              <RESULTS>
                <RESULT eventid="1108" points="112" reactiontime="+70" swimtime="00:01:58.73" resultid="1324" heatid="2272" lane="8" />
                <RESULT eventid="1140" points="153" swimtime="00:01:36.50" resultid="1325" heatid="2297" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="De Reginalda" birthdate="2011-07-22" gender="M" nation="BRA" license="400323" swrid="5717257" athleteid="1320" externalid="400323">
              <RESULTS>
                <RESULT eventid="1116" points="291" reactiontime="+58" swimtime="00:01:17.81" resultid="1321" heatid="2279" lane="2" />
                <RESULT eventid="1148" points="337" swimtime="00:01:07.31" resultid="1322" heatid="2305" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Arceli Silva" birthdate="2008-03-04" gender="M" nation="BRA" license="331565" swrid="5385686" athleteid="1301" externalid="331565" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1116" points="411" swimtime="00:01:09.40" resultid="1302" heatid="2281" lane="1" entrytime="00:01:12.35" entrycourse="LCM" />
                <RESULT eventid="1196" points="297" reactiontime="+72" swimtime="00:02:47.57" resultid="1303" heatid="2337" lane="2" entrytime="00:02:49.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marjori" lastname="Leticia Oliveira" birthdate="2011-05-23" gender="F" nation="BRA" license="406869" swrid="5717279" athleteid="1329" externalid="406869">
              <RESULTS>
                <RESULT eventid="1108" points="173" reactiontime="+82" swimtime="00:01:42.78" resultid="1330" heatid="2271" lane="6" />
                <RESULT eventid="1140" points="210" swimtime="00:01:26.97" resultid="1331" heatid="2297" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Cravcenco Marcondes" birthdate="2011-05-06" gender="M" nation="BRA" license="406867" athleteid="1326" externalid="406867">
              <RESULTS>
                <RESULT eventid="1116" points="149" swimtime="00:01:37.33" resultid="1327" heatid="2277" lane="1" />
                <RESULT eventid="1148" points="177" swimtime="00:01:23.37" resultid="1328" heatid="2306" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Reis" birthdate="2008-04-07" gender="F" nation="BRA" license="378820" swrid="5600243" athleteid="1311" externalid="378820" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1108" points="238" reactiontime="+80" swimtime="00:01:32.39" resultid="1312" heatid="2273" lane="7" entrytime="00:01:35.30" entrycourse="LCM" />
                <RESULT eventid="1204" points="138" swimtime="00:01:47.18" resultid="1313" heatid="2340" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Zanatta Flizikowski" birthdate="2007-09-14" gender="F" nation="BRA" license="366835" swrid="5600281" athleteid="1298" externalid="366835" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1124" points="275" swimtime="00:01:38.53" resultid="1299" heatid="2284" lane="4" entrytime="00:01:39.59" entrycourse="LCM" />
                <RESULT eventid="1156" points="223" swimtime="00:03:46.51" resultid="1300" heatid="2318" lane="8" entrytime="00:03:39.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:47.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="12782" nation="BRA" region="PR" clubid="1868" swrid="93773" name="Clube Duque De Caxias" shortname="Duque De Caxias">
          <ATHLETES>
            <ATHLETE firstname="Joao" lastname="Vitor Girelli" birthdate="2009-08-01" gender="M" nation="BRA" license="387965" swrid="5622312" athleteid="1869" externalid="387965">
              <RESULTS>
                <RESULT eventid="1116" points="314" reactiontime="+72" swimtime="00:01:15.90" resultid="1870" heatid="2277" lane="3" />
                <RESULT eventid="1084" points="370" swimtime="00:02:21.99" resultid="1871" heatid="2264" lane="6" entrytime="00:02:20.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="418" swimtime="00:01:02.65" resultid="1872" heatid="2312" lane="8" entrytime="00:01:02.36" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2539" nation="BRA" region="PR" clubid="1445" swrid="93771" name="Círculo Militar Do Paraná" shortname="Círculo Militar">
          <ATHLETES>
            <ATHLETE firstname="Fernando" lastname="Jun Melo Ogima" birthdate="2006-07-05" gender="M" nation="BRA" license="378332" swrid="5622284" athleteid="1449" externalid="378332">
              <RESULTS>
                <RESULT eventid="1132" points="274" swimtime="00:01:27.49" resultid="1450" heatid="2290" lane="5" />
                <RESULT eventid="1084" points="333" swimtime="00:02:27.05" resultid="1451" heatid="2263" lane="2" entrytime="00:02:27.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="226" swimtime="00:01:21.13" resultid="1452" heatid="2346" lane="2" />
                <RESULT eventid="1148" points="429" swimtime="00:01:02.12" resultid="1453" heatid="2311" lane="5" entrytime="00:01:02.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Vieira De Macedo Brasil" birthdate="2009-12-19" gender="F" nation="BRA" license="344143" swrid="5622311" athleteid="1446" externalid="344143">
              <RESULTS>
                <RESULT eventid="1076" points="375" swimtime="00:02:36.37" resultid="1447" heatid="2252" lane="3" entrytime="00:02:42.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="256" swimtime="00:03:36.48" resultid="1448" heatid="2318" lane="1" entrytime="00:03:34.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Manocchio" birthdate="2011-07-28" gender="M" nation="BRA" license="384916" swrid="5588573" athleteid="1457" externalid="384916">
              <RESULTS>
                <RESULT eventid="1132" points="214" swimtime="00:01:34.96" resultid="1458" heatid="2291" lane="2" />
                <RESULT eventid="1084" points="332" swimtime="00:02:27.18" resultid="1459" heatid="2262" lane="5" entrytime="00:02:34.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="344" swimtime="00:01:06.82" resultid="1460" heatid="2309" lane="1" entrytime="00:01:10.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Cavalcante Pierin" birthdate="2010-12-28" gender="M" nation="BRA" license="391227" swrid="5622269" athleteid="1461" externalid="391227">
              <RESULTS>
                <RESULT eventid="1116" points="185" reactiontime="+66" swimtime="00:01:30.47" resultid="1462" heatid="2279" lane="4" entrytime="00:01:35.85" entrycourse="LCM" />
                <RESULT eventid="1196" points="182" reactiontime="+86" swimtime="00:03:17.16" resultid="1463" heatid="2336" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="232" swimtime="00:01:16.19" resultid="1464" heatid="2307" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Maria Romanelli" birthdate="2011-04-18" gender="F" nation="BRA" license="378335" swrid="5588803" athleteid="1454" externalid="378335">
              <RESULTS>
                <RESULT eventid="1108" points="255" reactiontime="+86" swimtime="00:01:30.32" resultid="1455" heatid="2272" lane="4" entrytime="00:01:38.45" entrycourse="LCM" />
                <RESULT eventid="1140" points="379" swimtime="00:01:11.42" resultid="1456" heatid="2299" lane="5" entrytime="00:01:11.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Oliveira Martini" birthdate="2008-10-31" gender="M" nation="BRA" license="406953" swrid="5717285" athleteid="1479" externalid="406953">
              <RESULTS>
                <RESULT eventid="1084" points="261" swimtime="00:02:39.59" resultid="1480" heatid="2259" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="353" swimtime="00:01:06.27" resultid="1481" heatid="2304" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Torres Oliveira" birthdate="2008-04-10" gender="M" nation="BRA" license="400274" swrid="5653303" athleteid="1465" externalid="400274">
              <RESULTS>
                <RESULT eventid="1132" points="203" swimtime="00:01:36.78" resultid="1466" heatid="2293" lane="8" entrytime="00:01:30.32" entrycourse="LCM" />
                <RESULT eventid="1164" points="226" swimtime="00:03:25.96" resultid="1467" heatid="2321" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:37.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="320" swimtime="00:01:08.46" resultid="1468" heatid="2309" lane="2" entrytime="00:01:10.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Yamamoto" birthdate="2006-04-22" gender="M" nation="BRA" license="336569" swrid="5717304" athleteid="1469" externalid="336569">
              <RESULTS>
                <RESULT eventid="1212" points="253" swimtime="00:01:18.12" resultid="1470" heatid="2345" lane="3" />
                <RESULT eventid="1148" points="409" swimtime="00:01:03.12" resultid="1471" heatid="2305" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vicente" lastname="Bileski" birthdate="2011-06-29" gender="M" nation="BRA" license="406950" swrid="5717248" athleteid="1475" externalid="406950">
              <RESULTS>
                <RESULT eventid="1132" points="138" swimtime="00:01:49.98" resultid="1476" heatid="2288" lane="5" />
                <RESULT eventid="1116" points="136" reactiontime="+74" swimtime="00:01:40.27" resultid="1477" heatid="2278" lane="2" />
                <RESULT eventid="1148" points="168" swimtime="00:01:24.86" resultid="1478" heatid="2304" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thomas" lastname="Gomes" birthdate="2009-06-15" gender="M" nation="BRA" license="406948" swrid="5717268" athleteid="1472" externalid="406948">
              <RESULTS>
                <RESULT eventid="1084" points="177" swimtime="00:03:01.43" resultid="1473" heatid="2258" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="198" swimtime="00:01:20.37" resultid="1474" heatid="2306" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="263" nation="BRA" region="PR" clubid="1482" swrid="75436" name="Clube Curitibano" shortname="Curitibano">
          <ATHLETES>
            <ATHLETE firstname="Caua" lastname="Coelho" birthdate="2011-11-11" gender="M" nation="BRA" license="366889" swrid="5602527" athleteid="1681" externalid="366889">
              <RESULTS>
                <RESULT eventid="1100" points="251" swimtime="00:02:54.92" resultid="1682" heatid="2269" lane="5" entrytime="00:02:56.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1084" points="355" swimtime="00:02:23.93" resultid="1683" heatid="2263" lane="5" entrytime="00:02:26.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="275" swimtime="00:01:16.04" resultid="1684" heatid="2348" lane="8" entrytime="00:01:16.56" entrycourse="LCM" />
                <RESULT eventid="1180" points="396" swimtime="00:10:15.27" resultid="1685" heatid="2329" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.32" />
                    <SPLIT distance="200" swimtime="00:02:31.68" />
                    <SPLIT distance="300" swimtime="00:03:49.87" />
                    <SPLIT distance="400" swimtime="00:05:08.53" />
                    <SPLIT distance="500" swimtime="00:06:26.65" />
                    <SPLIT distance="600" swimtime="00:07:45.06" />
                    <SPLIT distance="700" swimtime="00:09:01.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Godino" birthdate="2010-04-27" gender="F" nation="BRA" license="356355" swrid="5600176" athleteid="1639" externalid="356355">
              <RESULTS>
                <RESULT eventid="1108" points="305" reactiontime="+79" swimtime="00:01:25.12" resultid="1640" heatid="2271" lane="7" />
                <RESULT eventid="1076" points="421" swimtime="00:02:30.46" resultid="1641" heatid="2254" lane="1" entrytime="00:02:32.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="306" swimtime="00:03:02.54" resultid="1642" heatid="2334" lane="1" entrytime="00:03:05.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="433" swimtime="00:10:40.44" resultid="1643" heatid="2327" lane="7" entrytime="00:10:50.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.23" />
                    <SPLIT distance="200" swimtime="00:02:35.91" />
                    <SPLIT distance="300" swimtime="00:03:56.69" />
                    <SPLIT distance="400" swimtime="00:05:17.77" />
                    <SPLIT distance="500" swimtime="00:06:39.28" />
                    <SPLIT distance="600" swimtime="00:08:00.49" />
                    <SPLIT distance="700" swimtime="00:09:21.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Gustavo Souza" birthdate="2011-08-24" gender="M" nation="BRA" license="366901" swrid="5588733" athleteid="1712" externalid="366901">
              <RESULTS>
                <RESULT eventid="1100" points="275" swimtime="00:02:49.53" resultid="1713" heatid="2269" lane="3" entrytime="00:03:06.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="294" swimtime="00:06:04.60" resultid="1714" heatid="2248" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.35" />
                    <SPLIT distance="200" swimtime="00:02:57.62" />
                    <SPLIT distance="300" swimtime="00:04:48.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="277" swimtime="00:01:15.78" resultid="1715" heatid="2347" lane="5" entrytime="00:01:17.57" entrycourse="LCM" />
                <RESULT eventid="1180" points="341" swimtime="00:10:46.59" resultid="1716" heatid="2328" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.69" />
                    <SPLIT distance="200" swimtime="00:02:42.00" />
                    <SPLIT distance="300" swimtime="00:04:04.09" />
                    <SPLIT distance="400" swimtime="00:05:27.96" />
                    <SPLIT distance="500" swimtime="00:06:48.67" />
                    <SPLIT distance="600" swimtime="00:08:09.51" />
                    <SPLIT distance="700" swimtime="00:09:30.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Bussmann" birthdate="2007-01-16" gender="F" nation="BRA" license="313781" swrid="5579983" athleteid="1513" externalid="313781">
              <RESULTS>
                <RESULT eventid="1124" points="593" swimtime="00:01:16.30" resultid="1514" heatid="2287" lane="5" entrytime="00:01:15.11" entrycourse="LCM" />
                <RESULT eventid="1076" points="537" swimtime="00:02:18.77" resultid="1515" heatid="2256" lane="2" entrytime="00:02:17.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="571" swimtime="00:02:45.77" resultid="1516" heatid="2320" lane="4" entrytime="00:02:39.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Felipe Paes Feres" birthdate="2008-07-28" gender="M" nation="BRA" license="307676" swrid="5600156" athleteid="1549" externalid="307676">
              <RESULTS>
                <RESULT eventid="1116" points="433" swimtime="00:01:08.19" resultid="1550" heatid="2282" lane="1" entrytime="00:01:06.99" entrycourse="LCM" />
                <RESULT eventid="1196" points="425" reactiontime="+64" swimtime="00:02:28.75" resultid="1551" heatid="2338" lane="4" entrytime="00:02:28.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo" lastname="De Lima Cavalcanti" birthdate="2009-12-17" gender="M" nation="BRA" license="380965" swrid="5634589" athleteid="1839" externalid="380965">
              <RESULTS>
                <RESULT eventid="1100" points="434" swimtime="00:02:25.66" resultid="1840" heatid="2270" lane="7" entrytime="00:02:37.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="513" swimtime="00:01:01.75" resultid="1841" heatid="2348" lane="3" entrytime="00:01:07.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Fantin Dias De Andrade" birthdate="2010-11-06" gender="F" nation="BRA" license="339262" swrid="5588684" athleteid="1763" externalid="339262">
              <RESULTS>
                <RESULT eventid="1124" points="274" swimtime="00:01:38.67" resultid="1764" heatid="2285" lane="5" entrytime="00:01:33.13" entrycourse="LCM" />
                <RESULT eventid="1108" points="263" reactiontime="+78" swimtime="00:01:29.38" resultid="1765" heatid="2273" lane="5" entrytime="00:01:28.94" entrycourse="LCM" />
                <RESULT eventid="1156" points="282" swimtime="00:03:29.67" resultid="1766" heatid="2318" lane="5" entrytime="00:03:20.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="342" swimtime="00:01:13.89" resultid="1767" heatid="2299" lane="1" entrytime="00:01:14.87" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Francisco Saldo" birthdate="2007-01-23" gender="M" nation="BRA" license="313537" swrid="5600169" athleteid="1517" externalid="313537">
              <RESULTS>
                <RESULT eventid="1100" status="DNS" swimtime="00:00:00.00" resultid="1518" heatid="2270" lane="4" entrytime="00:02:02.95" entrycourse="LCM" />
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="1519" heatid="2350" lane="5" entrytime="00:00:56.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Brandt De Macedo" birthdate="2010-01-13" gender="M" nation="BRA" license="338925" swrid="5588565" athleteid="1666" externalid="338925">
              <RESULTS>
                <RESULT eventid="1132" points="287" swimtime="00:01:26.16" resultid="1667" heatid="2290" lane="1" />
                <RESULT eventid="1084" points="433" swimtime="00:02:14.79" resultid="1668" heatid="2265" lane="6" entrytime="00:02:14.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="464" swimtime="00:09:43.59" resultid="1669" heatid="2331" lane="3" entrytime="00:09:34.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.93" />
                    <SPLIT distance="200" swimtime="00:02:18.33" />
                    <SPLIT distance="300" swimtime="00:03:31.61" />
                    <SPLIT distance="400" swimtime="00:04:46.23" />
                    <SPLIT distance="500" swimtime="00:06:01.35" />
                    <SPLIT distance="600" swimtime="00:07:15.97" />
                    <SPLIT distance="700" swimtime="00:08:30.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="433" swimtime="00:01:01.92" resultid="1670" heatid="2311" lane="3" entrytime="00:01:02.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Clivatti" birthdate="2010-05-24" gender="M" nation="BRA" license="368007" swrid="5600139" athleteid="1752" externalid="368007">
              <RESULTS>
                <RESULT eventid="1116" points="335" swimtime="00:01:14.24" resultid="1753" heatid="2279" lane="1" />
                <RESULT eventid="1084" points="492" swimtime="00:02:09.17" resultid="1754" heatid="2266" lane="7" entrytime="00:02:09.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="456" swimtime="00:09:47.14" resultid="1755" heatid="2331" lane="7" entrytime="00:09:46.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.62" />
                    <SPLIT distance="200" swimtime="00:02:17.08" />
                    <SPLIT distance="300" swimtime="00:03:30.31" />
                    <SPLIT distance="400" swimtime="00:04:44.78" />
                    <SPLIT distance="500" swimtime="00:06:00.75" />
                    <SPLIT distance="600" swimtime="00:07:17.25" />
                    <SPLIT distance="700" swimtime="00:08:33.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="480" swimtime="00:00:59.82" resultid="1756" heatid="2313" lane="1" entrytime="00:01:00.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Muxfeldt" birthdate="2011-05-13" gender="F" nation="BRA" license="366903" swrid="5602563" athleteid="1717" externalid="366903">
              <RESULTS>
                <RESULT eventid="1124" points="342" swimtime="00:01:31.66" resultid="1718" heatid="2286" lane="1" entrytime="00:01:28.54" entrycourse="LCM" />
                <RESULT eventid="1108" points="270" reactiontime="+82" swimtime="00:01:28.67" resultid="1719" heatid="2271" lane="4" />
                <RESULT eventid="1076" points="413" swimtime="00:02:31.44" resultid="1720" heatid="2253" lane="7" entrytime="00:02:37.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="359" swimtime="00:03:13.47" resultid="1721" heatid="2319" lane="2" entrytime="00:03:08.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="401" swimtime="00:01:10.07" resultid="1722" heatid="2296" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Moreira Segadaes" birthdate="2008-05-15" gender="M" nation="BRA" license="331574" swrid="5600220" athleteid="1510" externalid="331574">
              <RESULTS>
                <RESULT eventid="1132" points="547" swimtime="00:01:09.52" resultid="1511" heatid="2295" lane="2" entrytime="00:01:10.01" entrycourse="LCM" />
                <RESULT eventid="1164" points="545" swimtime="00:02:33.55" resultid="1512" heatid="2324" lane="2" entrytime="00:02:38.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Pereira Galle" birthdate="2011-08-02" gender="F" nation="BRA" license="369465" swrid="5627330" athleteid="1828" externalid="369465">
              <RESULTS>
                <RESULT eventid="1124" points="333" swimtime="00:01:32.46" resultid="1829" heatid="2286" lane="7" entrytime="00:01:28.00" entrycourse="LCM" />
                <RESULT eventid="1076" points="367" swimtime="00:02:37.59" resultid="1830" heatid="2254" lane="8" entrytime="00:02:33.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="230" swimtime="00:01:30.54" resultid="1831" heatid="2341" lane="1" />
                <RESULT eventid="1156" points="316" swimtime="00:03:21.89" resultid="1832" heatid="2317" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Artigas Pinheiro" birthdate="2011-08-25" gender="M" nation="BRA" license="377040" swrid="5588535" athleteid="1784" externalid="377040">
              <RESULTS>
                <RESULT eventid="1132" status="DSQ" swimtime="00:01:33.71" resultid="1785" heatid="2292" lane="5" entrytime="00:01:32.95" entrycourse="LCM" />
                <RESULT eventid="1100" points="208" swimtime="00:03:06.04" resultid="1786" heatid="2269" lane="6" entrytime="00:03:26.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1084" points="280" swimtime="00:02:35.91" resultid="1787" heatid="2257" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="186" swimtime="00:01:26.60" resultid="1788" heatid="2346" lane="5" entrytime="00:01:37.54" entrycourse="LCM" />
                <RESULT eventid="1164" points="285" swimtime="00:03:10.46" resultid="1789" heatid="2322" lane="6" entrytime="00:03:26.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Laurindo Netto" birthdate="2005-07-15" gender="M" nation="BRA" license="289995" swrid="5600198" athleteid="1495" externalid="289995">
              <RESULTS>
                <RESULT eventid="1068" points="544" swimtime="00:04:56.93" resultid="1496" heatid="2248" lane="4" entrytime="00:04:44.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.17" />
                    <SPLIT distance="200" swimtime="00:02:21.20" />
                    <SPLIT distance="300" swimtime="00:03:47.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="511" reactiontime="+71" swimtime="00:02:19.93" resultid="1497" heatid="2339" lane="3" entrytime="00:02:18.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="485" swimtime="00:02:39.69" resultid="1498" heatid="2324" lane="3" entrytime="00:02:32.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Cabrera Cirino" birthdate="2011-01-28" gender="M" nation="BRA" license="369531" swrid="5588569" athleteid="1757" externalid="369531">
              <RESULTS>
                <RESULT eventid="1116" points="393" reactiontime="+59" swimtime="00:01:10.40" resultid="1758" heatid="2281" lane="2" entrytime="00:01:11.59" entrycourse="LCM" />
                <RESULT eventid="1084" points="407" swimtime="00:02:17.63" resultid="1759" heatid="2258" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="262" swimtime="00:01:17.19" resultid="1760" heatid="2345" lane="2" />
                <RESULT eventid="1196" points="399" reactiontime="+64" swimtime="00:02:31.93" resultid="1761" heatid="2337" lane="5" entrytime="00:02:40.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="429" swimtime="00:01:02.09" resultid="1762" heatid="2311" lane="2" entrytime="00:01:03.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Sachser Rocha" birthdate="2008-07-09" gender="M" nation="BRA" license="330072" swrid="5600254" athleteid="1552" externalid="330072">
              <RESULTS>
                <RESULT eventid="1100" points="342" swimtime="00:02:37.64" resultid="1553" heatid="2269" lane="4" entrytime="00:02:56.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="500" swimtime="00:01:02.28" resultid="1554" heatid="2349" lane="3" entrytime="00:01:02.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Albuquerque" birthdate="2008-03-14" gender="F" nation="BRA" license="324787" swrid="5315259" athleteid="1483" externalid="324787">
              <RESULTS>
                <RESULT eventid="1124" points="546" swimtime="00:01:18.44" resultid="1484" heatid="2287" lane="3" entrytime="00:01:16.67" entrycourse="LCM" />
                <RESULT eventid="1156" points="509" swimtime="00:02:52.19" resultid="1485" heatid="2320" lane="3" entrytime="00:02:48.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Fontolan Gomes" birthdate="2010-07-02" gender="M" nation="BRA" license="356245" swrid="5588705" athleteid="1598" externalid="356245">
              <RESULTS>
                <RESULT eventid="1132" points="187" swimtime="00:01:39.34" resultid="1599" heatid="2290" lane="6" />
                <RESULT eventid="1116" points="356" reactiontime="+51" swimtime="00:01:12.75" resultid="1600" heatid="2281" lane="8" entrytime="00:01:14.51" entrycourse="LCM" />
                <RESULT eventid="1196" points="366" reactiontime="+77" swimtime="00:02:36.38" resultid="1601" heatid="2337" lane="4" entrytime="00:02:38.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="345" swimtime="00:01:06.79" resultid="1602" heatid="2308" lane="5" entrytime="00:01:11.51" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="De Krinski" birthdate="2007-07-20" gender="M" nation="BRA" license="334494" swrid="5600148" athleteid="1849" externalid="334494">
              <RESULTS>
                <RESULT eventid="1116" points="547" reactiontime="+71" swimtime="00:01:03.08" resultid="1850" heatid="2282" lane="5" entrytime="00:01:01.65" entrycourse="LCM" />
                <RESULT eventid="1196" points="488" swimtime="00:02:22.07" resultid="1851" heatid="2339" lane="1" entrytime="00:02:19.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicole" lastname="Rosario Osternack" birthdate="2008-04-11" gender="F" nation="BRA" license="331584" swrid="5600248" athleteid="1489" externalid="331584">
              <RESULTS>
                <RESULT eventid="1108" points="485" reactiontime="+67" swimtime="00:01:12.93" resultid="1490" heatid="2276" lane="2" entrytime="00:01:10.78" entrycourse="LCM" />
                <RESULT eventid="1204" points="531" swimtime="00:01:08.51" resultid="1491" heatid="2343" lane="3" entrytime="00:01:07.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="De Albuquerque" birthdate="2010-06-08" gender="F" nation="BRA" license="356249" swrid="5600145" athleteid="1603" externalid="356249">
              <RESULTS>
                <RESULT eventid="1124" points="267" swimtime="00:01:39.53" resultid="1604" heatid="2283" lane="6" />
                <RESULT eventid="1108" points="404" reactiontime="+61" swimtime="00:01:17.53" resultid="1605" heatid="2276" lane="8" entrytime="00:01:16.20" entrycourse="LCM" />
                <RESULT eventid="1188" points="387" reactiontime="+78" swimtime="00:02:48.93" resultid="1606" heatid="2335" lane="2" entrytime="00:02:45.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="390" swimtime="00:01:10.76" resultid="1607" heatid="2300" lane="8" entrytime="00:01:10.55" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Schiavon" birthdate="2010-05-03" gender="M" nation="BRA" license="356354" swrid="5600256" athleteid="1634" externalid="356354">
              <RESULTS>
                <RESULT eventid="1116" points="283" reactiontime="+60" swimtime="00:01:18.59" resultid="1635" heatid="2279" lane="3" />
                <RESULT eventid="1084" points="432" swimtime="00:02:14.92" resultid="1636" heatid="2265" lane="8" entrytime="00:02:17.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="479" swimtime="00:09:37.49" resultid="1637" heatid="2331" lane="1" entrytime="00:09:50.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.09" />
                    <SPLIT distance="200" swimtime="00:02:18.11" />
                    <SPLIT distance="300" swimtime="00:03:31.23" />
                    <SPLIT distance="400" swimtime="00:04:45.21" />
                    <SPLIT distance="500" swimtime="00:05:59.11" />
                    <SPLIT distance="600" swimtime="00:07:12.68" />
                    <SPLIT distance="700" swimtime="00:08:26.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="414" swimtime="00:01:02.83" resultid="1638" heatid="2310" lane="5" entrytime="00:01:05.05" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helen" lastname="Barato Bernardi" birthdate="2006-07-27" gender="F" nation="BRA" license="317031" swrid="5717244" athleteid="1842" externalid="317031">
              <RESULTS>
                <RESULT eventid="1124" points="606" swimtime="00:01:15.75" resultid="1843" heatid="2287" lane="4" entrytime="00:01:14.91" entrycourse="LCM" />
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="1844" heatid="2320" lane="5" entrytime="00:02:45.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Clara Fernandes Pereira" birthdate="2009-11-19" gender="F" nation="BRA" license="344340" swrid="5600137" athleteid="1486" externalid="344340">
              <RESULTS>
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="1487" heatid="2256" lane="7" entrytime="00:02:17.87" entrycourse="LCM" />
                <RESULT eventid="1172" status="WDR" swimtime="00:00:00.00" resultid="1488" heatid="2327" lane="5" entrytime="00:10:05.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Kirchgassner" birthdate="2007-02-10" gender="M" nation="BRA" license="313535" swrid="5600230" athleteid="1538" externalid="313535">
              <RESULTS>
                <RESULT eventid="1132" points="597" swimtime="00:01:07.55" resultid="1539" heatid="2295" lane="5" entrytime="00:01:05.67" entrycourse="LCM" />
                <RESULT eventid="1212" points="501" swimtime="00:01:02.25" resultid="1540" heatid="2349" lane="4" entrytime="00:01:01.35" entrycourse="LCM" />
                <RESULT eventid="1164" points="606" swimtime="00:02:28.27" resultid="1541" heatid="2324" lane="4" entrytime="00:02:21.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Pellanda" birthdate="2010-11-12" gender="M" nation="BRA" license="356352" swrid="5600233" athleteid="1624" externalid="356352">
              <RESULTS>
                <RESULT eventid="1116" points="340" reactiontime="+81" swimtime="00:01:13.88" resultid="1625" heatid="2280" lane="3" entrytime="00:01:17.90" entrycourse="LCM" />
                <RESULT eventid="1084" points="513" swimtime="00:02:07.35" resultid="1626" heatid="2266" lane="8" entrytime="00:02:11.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="539" swimtime="00:09:15.51" resultid="1627" heatid="2331" lane="4" entrytime="00:09:22.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.93" />
                    <SPLIT distance="200" swimtime="00:02:16.93" />
                    <SPLIT distance="300" swimtime="00:03:27.77" />
                    <SPLIT distance="400" swimtime="00:04:38.89" />
                    <SPLIT distance="500" swimtime="00:05:48.36" />
                    <SPLIT distance="600" swimtime="00:06:58.39" />
                    <SPLIT distance="700" swimtime="00:08:08.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="479" swimtime="00:00:59.88" resultid="1628" heatid="2312" lane="6" entrytime="00:01:00.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolau" lastname="Neto" birthdate="2011-03-22" gender="M" nation="BRA" license="366906" swrid="5602565" athleteid="1729" externalid="366906">
              <RESULTS>
                <RESULT eventid="1132" points="305" swimtime="00:01:24.42" resultid="1730" heatid="2293" lane="7" entrytime="00:01:28.66" entrycourse="LCM" />
                <RESULT eventid="1068" points="312" swimtime="00:05:57.46" resultid="1731" heatid="2247" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.70" />
                    <SPLIT distance="200" swimtime="00:03:07.44" />
                    <SPLIT distance="300" swimtime="00:04:40.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="357" swimtime="00:10:36.88" resultid="1732" heatid="2329" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.81" />
                    <SPLIT distance="200" swimtime="00:02:34.24" />
                    <SPLIT distance="300" swimtime="00:03:56.18" />
                    <SPLIT distance="400" swimtime="00:05:17.14" />
                    <SPLIT distance="500" swimtime="00:06:39.34" />
                    <SPLIT distance="600" swimtime="00:08:01.31" />
                    <SPLIT distance="700" swimtime="00:09:20.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="302" swimtime="00:03:07.01" resultid="1733" heatid="2323" lane="8" entrytime="00:03:08.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="380" swimtime="00:01:04.66" resultid="1734" heatid="2304" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Sabedotti" birthdate="2002-07-07" gender="M" nation="BRA" license="134704" swrid="5600252" athleteid="1589" externalid="134704" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1132" points="658" swimtime="00:01:05.38" resultid="1590" heatid="2295" lane="4" entrytime="00:01:04.14" entrycourse="LCM" />
                <RESULT eventid="1212" points="657" swimtime="00:00:56.88" resultid="1591" heatid="2350" lane="4" entrytime="00:00:55.31" entrycourse="LCM" />
                <RESULT eventid="1148" points="698" swimtime="00:00:52.82" resultid="1592" heatid="2315" lane="3" entrytime="00:00:52.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Fontana Moraes" birthdate="2006-08-17" gender="M" nation="BRA" license="296593" swrid="5600163" athleteid="1542" externalid="296593">
              <RESULTS>
                <RESULT eventid="1084" points="274" swimtime="00:02:36.86" resultid="1543" heatid="2263" lane="8" entrytime="00:02:31.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="293" swimtime="00:11:20.15" resultid="1544" heatid="2329" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.16" />
                    <SPLIT distance="200" swimtime="00:02:46.55" />
                    <SPLIT distance="300" swimtime="00:04:14.18" />
                    <SPLIT distance="400" swimtime="00:05:41.20" />
                    <SPLIT distance="500" swimtime="00:07:07.57" />
                    <SPLIT distance="600" swimtime="00:08:33.89" />
                    <SPLIT distance="700" swimtime="00:09:59.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="301" swimtime="00:01:09.90" resultid="1545" heatid="2310" lane="2" entrytime="00:01:06.57" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Galvao" birthdate="2011-03-11" gender="M" nation="BRA" license="381989" swrid="5602541" athleteid="1793" externalid="381989">
              <RESULTS>
                <RESULT eventid="1132" points="184" swimtime="00:01:39.98" resultid="1794" heatid="2291" lane="8" />
                <RESULT eventid="1116" points="154" reactiontime="+62" swimtime="00:01:36.12" resultid="1795" heatid="2278" lane="8" />
                <RESULT eventid="1084" points="290" swimtime="00:02:33.96" resultid="1796" heatid="2262" lane="2" entrytime="00:02:38.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="317" swimtime="00:11:03.00" resultid="1797" heatid="2329" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.09" />
                    <SPLIT distance="200" swimtime="00:02:43.05" />
                    <SPLIT distance="300" swimtime="00:04:06.85" />
                    <SPLIT distance="400" swimtime="00:05:31.24" />
                    <SPLIT distance="500" swimtime="00:06:56.15" />
                    <SPLIT distance="600" swimtime="00:08:20.90" />
                    <SPLIT distance="700" swimtime="00:09:44.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="321" swimtime="00:01:08.37" resultid="1798" heatid="2308" lane="3" entrytime="00:01:11.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Kremer De Aguiar" birthdate="2009-12-22" gender="F" nation="BRA" license="338987" swrid="5600196" athleteid="1570" externalid="338987">
              <RESULTS>
                <RESULT eventid="1124" points="427" swimtime="00:01:25.14" resultid="1571" heatid="2286" lane="5" entrytime="00:01:25.51" entrycourse="LCM" />
                <RESULT eventid="1156" points="411" swimtime="00:03:04.87" resultid="1572" heatid="2319" lane="5" entrytime="00:03:03.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Leao" birthdate="2011-09-18" gender="M" nation="BRA" license="366880" swrid="5602553" athleteid="1675" externalid="366880">
              <RESULTS>
                <RESULT eventid="1116" points="240" reactiontime="+76" swimtime="00:01:23.02" resultid="1676" heatid="2278" lane="4" />
                <RESULT eventid="1084" points="346" swimtime="00:02:25.17" resultid="1677" heatid="2261" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="226" swimtime="00:01:21.13" resultid="1678" heatid="2346" lane="4" entrytime="00:01:31.40" entrycourse="LCM" />
                <RESULT eventid="1180" points="379" swimtime="00:10:24.25" resultid="1679" heatid="2329" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.86" />
                    <SPLIT distance="200" swimtime="00:02:34.81" />
                    <SPLIT distance="300" swimtime="00:03:54.30" />
                    <SPLIT distance="400" swimtime="00:05:13.17" />
                    <SPLIT distance="500" swimtime="00:06:32.69" />
                    <SPLIT distance="600" swimtime="00:07:51.66" />
                    <SPLIT distance="700" swimtime="00:09:10.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="357" swimtime="00:01:06.02" resultid="1680" heatid="2309" lane="3" entrytime="00:01:09.41" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Krupacz" birthdate="2008-04-18" gender="F" nation="BRA" license="329187" swrid="5634611" athleteid="1836" externalid="329187">
              <RESULTS>
                <RESULT eventid="1108" points="550" reactiontime="+66" swimtime="00:01:09.97" resultid="1837" heatid="2276" lane="3" entrytime="00:01:08.91" entrycourse="LCM" />
                <RESULT eventid="1188" status="DNS" swimtime="00:00:00.00" resultid="1838" heatid="2335" lane="4" entrytime="00:02:32.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Fontoura" birthdate="2010-08-26" gender="M" nation="BRA" license="338922" swrid="5600167" athleteid="1656" externalid="338922">
              <RESULTS>
                <RESULT eventid="1132" points="249" swimtime="00:01:30.37" resultid="1657" heatid="2291" lane="6" />
                <RESULT eventid="1068" points="308" swimtime="00:05:59.03" resultid="1658" heatid="2247" lane="5" />
                <RESULT eventid="1212" points="258" swimtime="00:01:17.61" resultid="1659" heatid="2347" lane="2" entrytime="00:01:24.76" entrycourse="LCM" />
                <RESULT eventid="1148" points="368" swimtime="00:01:05.38" resultid="1660" heatid="2309" lane="4" entrytime="00:01:08.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joshua" lastname="Gomide Capraro" birthdate="2009-01-18" gender="M" nation="BRA" license="339030" swrid="5600177" athleteid="1503" externalid="339030">
              <RESULTS>
                <RESULT eventid="1084" points="535" swimtime="00:02:05.62" resultid="1504" heatid="2267" lane="7" entrytime="00:02:03.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="404" swimtime="00:10:11.49" resultid="1505" heatid="2331" lane="6" entrytime="00:09:42.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.53" />
                    <SPLIT distance="200" swimtime="00:02:17.24" />
                    <SPLIT distance="300" swimtime="00:03:32.57" />
                    <SPLIT distance="400" swimtime="00:04:51.03" />
                    <SPLIT distance="500" swimtime="00:06:11.44" />
                    <SPLIT distance="600" swimtime="00:07:32.41" />
                    <SPLIT distance="700" swimtime="00:08:52.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="601" swimtime="00:00:55.50" resultid="1506" heatid="2314" lane="5" entrytime="00:00:55.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Presiazniuk" birthdate="2010-10-14" gender="M" nation="BRA" license="356353" swrid="5600237" athleteid="1629" externalid="356353">
              <RESULTS>
                <RESULT eventid="1116" points="376" reactiontime="+67" swimtime="00:01:11.43" resultid="1630" heatid="2281" lane="6" entrytime="00:01:11.48" entrycourse="LCM" />
                <RESULT eventid="1084" points="431" swimtime="00:02:14.95" resultid="1631" heatid="2265" lane="3" entrytime="00:02:14.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="390" reactiontime="+70" swimtime="00:02:33.13" resultid="1632" heatid="2338" lane="2" entrytime="00:02:33.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="457" swimtime="00:01:00.81" resultid="1633" heatid="2312" lane="5" entrytime="00:01:00.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="LIV" lastname="Carvalho" birthdate="2011-09-13" gender="F" nation="BRA" license="366899" swrid="5602524" athleteid="1707" externalid="366899">
              <RESULTS>
                <RESULT eventid="1124" points="284" swimtime="00:01:37.48" resultid="1708" heatid="2284" lane="6" entrytime="00:01:47.56" entrycourse="LCM" />
                <RESULT eventid="1076" points="279" swimtime="00:02:52.54" resultid="1709" heatid="2252" lane="8" entrytime="00:02:53.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="136" swimtime="00:01:47.76" resultid="1710" heatid="2342" lane="7" entrytime="00:01:47.78" entrycourse="LCM" />
                <RESULT eventid="1156" points="310" swimtime="00:03:23.22" resultid="1711" heatid="2316" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Lacerda" birthdate="2011-05-09" gender="M" nation="BRA" license="366909" swrid="5602550" athleteid="1746" externalid="366909">
              <RESULTS>
                <RESULT eventid="1132" points="257" swimtime="00:01:29.37" resultid="1747" heatid="2293" lane="1" entrytime="00:01:28.88" entrycourse="LCM" />
                <RESULT eventid="1084" points="334" swimtime="00:02:27.00" resultid="1748" heatid="2259" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="310" swimtime="00:05:57.95" resultid="1749" heatid="2248" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.76" />
                    <SPLIT distance="200" swimtime="00:03:01.64" />
                    <SPLIT distance="300" swimtime="00:04:42.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="289" swimtime="00:03:09.73" resultid="1750" heatid="2322" lane="5" entrytime="00:03:14.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="343" swimtime="00:01:06.89" resultid="1751" heatid="2309" lane="6" entrytime="00:01:09.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Mattioli" birthdate="2011-10-22" gender="F" nation="BRA" license="366896" swrid="5602559" athleteid="1696" externalid="366896">
              <RESULTS>
                <RESULT eventid="1124" points="335" swimtime="00:01:32.25" resultid="1697" heatid="2285" lane="3" entrytime="00:01:33.28" entrycourse="LCM" />
                <RESULT eventid="1076" points="420" swimtime="00:02:30.68" resultid="1698" heatid="2249" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="336" swimtime="00:03:17.75" resultid="1699" heatid="2318" lane="4" entrytime="00:03:18.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="405" swimtime="00:01:09.84" resultid="1700" heatid="2296" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Rocha Silva" birthdate="2007-10-10" gender="M" nation="BRA" license="372280" swrid="5717294" athleteid="1535" externalid="372280">
              <RESULTS>
                <RESULT eventid="1084" points="701" swimtime="00:01:54.78" resultid="1536" heatid="2267" lane="5" entrytime="00:01:54.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="717" swimtime="00:00:52.34" resultid="1537" heatid="2315" lane="4" entrytime="00:00:51.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manoela" lastname="Andrade" birthdate="2010-03-10" gender="F" nation="BRA" license="339042" swrid="5363102" athleteid="1661" externalid="339042">
              <RESULTS>
                <RESULT eventid="1108" points="238" reactiontime="+67" swimtime="00:01:32.40" resultid="1662" heatid="2274" lane="8" entrytime="00:01:26.95" entrycourse="LCM" />
                <RESULT eventid="1076" points="364" swimtime="00:02:37.96" resultid="1663" heatid="2253" lane="5" entrytime="00:02:34.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="225" swimtime="00:01:31.11" resultid="1664" heatid="2342" lane="4" entrytime="00:01:19.51" entrycourse="LCM" />
                <RESULT eventid="1172" points="402" swimtime="00:10:56.37" resultid="1665" heatid="2327" lane="2" entrytime="00:10:49.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.28" />
                    <SPLIT distance="200" swimtime="00:02:38.85" />
                    <SPLIT distance="300" swimtime="00:04:02.79" />
                    <SPLIT distance="400" swimtime="00:05:27.29" />
                    <SPLIT distance="500" swimtime="00:06:52.69" />
                    <SPLIT distance="600" swimtime="00:08:14.59" />
                    <SPLIT distance="700" swimtime="00:09:36.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Correa Nascimento" birthdate="2009-01-19" gender="M" nation="BRA" license="342235" swrid="5600140" athleteid="1564" externalid="342235">
              <RESULTS>
                <RESULT eventid="1132" status="DNS" swimtime="00:00:00.00" resultid="1565" heatid="2290" lane="8" />
                <RESULT eventid="1148" status="DNS" swimtime="00:00:00.00" resultid="1566" heatid="2313" lane="5" entrytime="00:00:58.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietra" lastname="Ruschel Carvalho" birthdate="2009-03-21" gender="F" nation="BRA" license="324999" swrid="5600250" athleteid="1492" externalid="324999">
              <RESULTS>
                <RESULT eventid="1076" points="573" swimtime="00:02:15.84" resultid="1493" heatid="2256" lane="3" entrytime="00:02:13.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="606" swimtime="00:01:01.08" resultid="1494" heatid="2302" lane="3" entrytime="00:01:01.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Carneiro Silva" birthdate="2011-02-21" gender="F" nation="BRA" license="390924" swrid="5602522" athleteid="1823" externalid="390924">
              <RESULTS>
                <RESULT eventid="1108" points="351" reactiontime="+75" swimtime="00:01:21.20" resultid="1824" heatid="2274" lane="3" entrytime="00:01:22.75" entrycourse="LCM" />
                <RESULT eventid="1076" points="336" swimtime="00:02:42.32" resultid="1825" heatid="2252" lane="6" entrytime="00:02:43.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="148" swimtime="00:01:44.66" resultid="1826" heatid="2341" lane="7" />
                <RESULT eventid="1188" points="298" reactiontime="+74" swimtime="00:03:04.26" resultid="1827" heatid="2334" lane="8" entrytime="00:03:05.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Estevao" lastname="Valduga Artigas" birthdate="2009-06-01" gender="M" nation="BRA" license="339556" swrid="5600267" athleteid="1561" externalid="339556">
              <RESULTS>
                <RESULT eventid="1116" points="273" swimtime="00:01:19.46" resultid="1562" heatid="2280" lane="1" entrytime="00:01:23.63" entrycourse="LCM" />
                <RESULT eventid="1180" points="332" swimtime="00:10:52.57" resultid="1563" heatid="2330" lane="2" entrytime="00:10:48.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.26" />
                    <SPLIT distance="200" swimtime="00:02:36.28" />
                    <SPLIT distance="300" swimtime="00:03:58.94" />
                    <SPLIT distance="400" swimtime="00:05:22.90" />
                    <SPLIT distance="500" swimtime="00:06:47.03" />
                    <SPLIT distance="600" swimtime="00:08:10.36" />
                    <SPLIT distance="700" swimtime="00:09:33.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Zaroni" birthdate="2010-03-03" gender="F" nation="BRA" license="356345" swrid="5600282" athleteid="1523" externalid="356345">
              <RESULTS>
                <RESULT eventid="1124" points="423" swimtime="00:01:25.39" resultid="1524" heatid="2287" lane="2" entrytime="00:01:21.40" entrycourse="LCM" />
                <RESULT eventid="1076" points="421" swimtime="00:02:30.49" resultid="1525" heatid="2254" lane="4" entrytime="00:02:30.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="230" swimtime="00:01:30.46" resultid="1526" heatid="2342" lane="8" />
                <RESULT eventid="1156" points="442" swimtime="00:03:00.48" resultid="1527" heatid="2320" lane="2" entrytime="00:02:56.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabelly" lastname="Sinnott" birthdate="2009-03-14" gender="F" nation="BRA" license="367255" swrid="5600258" athleteid="1520" externalid="367255">
              <RESULTS>
                <RESULT eventid="1076" points="595" swimtime="00:02:14.14" resultid="1521" heatid="2256" lane="5" entrytime="00:02:12.13" entrycourse="LCM" />
                <RESULT eventid="1172" points="526" swimtime="00:10:00.22" resultid="1522" heatid="2327" lane="4" entrytime="00:09:47.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.43" />
                    <SPLIT distance="200" swimtime="00:02:22.63" />
                    <SPLIT distance="300" swimtime="00:03:38.48" />
                    <SPLIT distance="400" swimtime="00:04:55.04" />
                    <SPLIT distance="500" swimtime="00:06:11.63" />
                    <SPLIT distance="600" swimtime="00:07:28.28" />
                    <SPLIT distance="700" swimtime="00:08:45.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fernandes" birthdate="2010-03-13" gender="M" nation="BRA" license="339266" swrid="5588695" athleteid="1811" externalid="339266">
              <RESULTS>
                <RESULT eventid="1116" points="425" reactiontime="+68" swimtime="00:01:08.63" resultid="1812" heatid="2281" lane="3" entrytime="00:01:09.53" entrycourse="LCM" />
                <RESULT eventid="1084" points="437" swimtime="00:02:14.39" resultid="1813" heatid="2265" lane="5" entrytime="00:02:14.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="404" reactiontime="+73" swimtime="00:02:31.33" resultid="1814" heatid="2338" lane="5" entrytime="00:02:30.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="491" swimtime="00:00:59.39" resultid="1815" heatid="2313" lane="2" entrytime="00:00:59.82" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Fontana" birthdate="2011-12-29" gender="M" nation="BRA" license="366897" swrid="5602539" athleteid="1701" externalid="366897">
              <RESULTS>
                <RESULT eventid="1132" points="152" swimtime="00:01:46.55" resultid="1702" heatid="2292" lane="8" entrytime="00:01:51.66" entrycourse="LCM" />
                <RESULT eventid="1116" points="172" swimtime="00:01:32.65" resultid="1703" heatid="2279" lane="8" />
                <RESULT eventid="1084" points="190" swimtime="00:02:57.40" resultid="1704" heatid="2260" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="174" swimtime="00:03:44.36" resultid="1705" heatid="2322" lane="7" entrytime="00:04:00.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:49.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="194" swimtime="00:01:20.87" resultid="1706" heatid="2307" lane="6" entrytime="00:01:20.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Henrique Pasqual" birthdate="2005-05-07" gender="M" nation="BRA" license="329284" swrid="5600185" athleteid="1855" externalid="329284">
              <RESULTS>
                <RESULT eventid="1084" points="531" swimtime="00:02:05.95" resultid="1856" heatid="2267" lane="2" entrytime="00:02:01.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="480" swimtime="00:01:03.12" resultid="1857" heatid="2350" lane="2" entrytime="00:00:58.79" entrycourse="LCM" />
                <RESULT eventid="1148" points="613" swimtime="00:00:55.15" resultid="1858" heatid="2315" lane="6" entrytime="00:00:53.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelo" lastname="Vanhazebrouck" birthdate="2010-01-09" gender="M" nation="BRA" license="339043" swrid="5600269" athleteid="1593" externalid="339043">
              <RESULTS>
                <RESULT eventid="1132" points="310" swimtime="00:01:24.04" resultid="1594" heatid="2293" lane="3" entrytime="00:01:23.11" entrycourse="LCM" />
                <RESULT eventid="1084" points="415" swimtime="00:02:16.65" resultid="1595" heatid="2265" lane="1" entrytime="00:02:17.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="295" swimtime="00:03:08.41" resultid="1596" heatid="2323" lane="7" entrytime="00:03:02.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="447" swimtime="00:01:01.27" resultid="1597" heatid="2312" lane="3" entrytime="00:01:00.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Fontolan Gomes" birthdate="2008-05-01" gender="M" nation="BRA" license="307667" swrid="5600166" athleteid="1546" externalid="307667">
              <RESULTS>
                <RESULT eventid="1116" points="379" reactiontime="+75" swimtime="00:01:11.25" resultid="1547" heatid="2281" lane="5" entrytime="00:01:09.02" entrycourse="LCM" />
                <RESULT eventid="1196" points="384" reactiontime="+76" swimtime="00:02:33.88" resultid="1548" heatid="2338" lane="6" entrytime="00:02:32.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Emili Da Silva Gomes Xavier" birthdate="2010-09-08" gender="F" nation="BRA" license="372519" swrid="5717260" athleteid="1862" externalid="372519">
              <RESULTS>
                <RESULT eventid="1124" points="351" swimtime="00:01:30.91" resultid="1863" heatid="2285" lane="6" entrytime="00:01:33.31" entrycourse="LCM" />
                <RESULT eventid="1108" points="320" reactiontime="+74" swimtime="00:01:23.79" resultid="1864" heatid="2274" lane="2" entrytime="00:01:22.97" entrycourse="LCM" />
                <RESULT eventid="1076" points="379" swimtime="00:02:35.87" resultid="1865" heatid="2250" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="333" swimtime="00:02:57.49" resultid="1866" heatid="2334" lane="7" entrytime="00:03:04.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="291" swimtime="00:03:27.36" resultid="1867" heatid="2318" lane="6" entrytime="00:03:30.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:40.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Geremia" birthdate="2011-07-20" gender="F" nation="BRA" license="366908" swrid="5602543" athleteid="1740" externalid="366908">
              <RESULTS>
                <RESULT eventid="1108" points="392" reactiontime="+62" swimtime="00:01:18.33" resultid="1741" heatid="2275" lane="6" entrytime="00:01:19.15" entrycourse="LCM" />
                <RESULT eventid="1076" points="479" swimtime="00:02:24.21" resultid="1742" heatid="2250" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="394" reactiontime="+68" swimtime="00:02:47.87" resultid="1743" heatid="2334" lane="5" entrytime="00:02:53.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="459" swimtime="00:10:28.08" resultid="1744" heatid="2326" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.82" />
                    <SPLIT distance="200" swimtime="00:02:35.57" />
                    <SPLIT distance="300" swimtime="00:03:56.49" />
                    <SPLIT distance="400" swimtime="00:05:16.67" />
                    <SPLIT distance="500" swimtime="00:06:36.12" />
                    <SPLIT distance="600" swimtime="00:07:54.58" />
                    <SPLIT distance="700" swimtime="00:09:12.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="473" swimtime="00:01:06.33" resultid="1745" heatid="2301" lane="8" entrytime="00:01:07.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorena" lastname="Mascarenhas" birthdate="2011-08-31" gender="F" nation="BRA" license="370581" swrid="5602558" athleteid="1768" externalid="370581">
              <RESULTS>
                <RESULT eventid="1108" points="361" reactiontime="+39" swimtime="00:01:20.45" resultid="1769" heatid="2274" lane="5" entrytime="00:01:22.71" entrycourse="LCM" />
                <RESULT eventid="1076" points="391" swimtime="00:02:34.25" resultid="1770" heatid="2252" lane="4" entrytime="00:02:41.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="383" reactiontime="+69" swimtime="00:02:49.49" resultid="1771" heatid="2334" lane="2" entrytime="00:02:59.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="397" swimtime="00:01:10.32" resultid="1772" heatid="2297" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gael" lastname="Gluck" birthdate="2011-01-28" gender="M" nation="BRA" license="366891" swrid="5588726" athleteid="1686" externalid="366891">
              <RESULTS>
                <RESULT eventid="1132" points="305" swimtime="00:01:24.43" resultid="1687" heatid="2293" lane="6" entrytime="00:01:27.02" entrycourse="LCM" />
                <RESULT eventid="1084" points="346" swimtime="00:02:25.19" resultid="1688" heatid="2258" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="319" swimtime="00:03:03.53" resultid="1689" heatid="2323" lane="1" entrytime="00:03:05.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="348" swimtime="00:01:06.61" resultid="1690" heatid="2305" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Vieira Motta" birthdate="2009-09-19" gender="M" nation="BRA" license="339064" swrid="5600271" athleteid="1582" externalid="339064">
              <RESULTS>
                <RESULT eventid="1116" points="418" reactiontime="+72" swimtime="00:01:09.00" resultid="1583" heatid="2281" lane="7" entrytime="00:01:11.84" entrycourse="LCM" />
                <RESULT eventid="1196" points="388" swimtime="00:02:33.35" resultid="1584" heatid="2338" lane="1" entrytime="00:02:36.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="442" swimtime="00:09:53.50" resultid="1585" heatid="2330" lane="5" entrytime="00:10:03.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.57" />
                    <SPLIT distance="200" swimtime="00:02:24.94" />
                    <SPLIT distance="300" swimtime="00:03:39.47" />
                    <SPLIT distance="400" swimtime="00:04:54.75" />
                    <SPLIT distance="500" swimtime="00:06:09.45" />
                    <SPLIT distance="600" swimtime="00:07:24.49" />
                    <SPLIT distance="700" swimtime="00:08:39.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rene" lastname="Osternack Erbe" birthdate="2011-04-03" gender="M" nation="BRA" license="366907" swrid="5588842" athleteid="1735" externalid="366907">
              <RESULTS>
                <RESULT eventid="1116" points="255" reactiontime="+84" swimtime="00:01:21.28" resultid="1736" heatid="2280" lane="6" entrytime="00:01:21.81" entrycourse="LCM" />
                <RESULT eventid="1068" points="246" swimtime="00:06:26.82" resultid="1737" heatid="2247" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.85" />
                    <SPLIT distance="200" swimtime="00:03:03.95" />
                    <SPLIT distance="300" swimtime="00:05:04.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="163" swimtime="00:01:30.41" resultid="1738" heatid="2347" lane="8" entrytime="00:01:26.65" entrycourse="LCM" />
                <RESULT eventid="1180" points="307" swimtime="00:11:09.94" resultid="1739" heatid="2328" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.81" />
                    <SPLIT distance="200" swimtime="00:02:44.42" />
                    <SPLIT distance="300" swimtime="00:04:09.10" />
                    <SPLIT distance="400" swimtime="00:05:34.59" />
                    <SPLIT distance="500" swimtime="00:06:58.97" />
                    <SPLIT distance="600" swimtime="00:08:25.33" />
                    <SPLIT distance="700" swimtime="00:09:49.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="David Cella" birthdate="2008-02-17" gender="M" nation="BRA" license="341107" swrid="5634581" athleteid="1833" externalid="341107">
              <RESULTS>
                <RESULT eventid="1132" points="475" swimtime="00:01:12.89" resultid="1834" heatid="2295" lane="7" entrytime="00:01:11.28" entrycourse="LCM" />
                <RESULT eventid="1148" points="601" swimtime="00:00:55.52" resultid="1835" heatid="2314" lane="3" entrytime="00:00:55.13" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Valduga Artigas" birthdate="2009-06-01" gender="M" nation="BRA" license="339569" swrid="5600268" athleteid="1579" externalid="339569">
              <RESULTS>
                <RESULT eventid="1212" points="282" swimtime="00:01:15.33" resultid="1580" heatid="2347" lane="4" entrytime="00:01:17.32" entrycourse="LCM" />
                <RESULT eventid="1148" points="361" swimtime="00:01:05.80" resultid="1581" heatid="2310" lane="1" entrytime="00:01:07.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Yolanda Ferreira" birthdate="2008-03-17" gender="F" nation="BRA" license="358335" swrid="5600276" athleteid="1773" externalid="358335">
              <RESULTS>
                <RESULT eventid="1124" points="483" swimtime="00:01:21.73" resultid="1774" heatid="2287" lane="6" entrytime="00:01:21.18" entrycourse="LCM" />
                <RESULT eventid="1156" points="463" swimtime="00:02:57.70" resultid="1775" heatid="2320" lane="6" entrytime="00:02:55.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Ramos Marcon" birthdate="2008-01-12" gender="M" nation="BRA" license="372281" swrid="5600240" athleteid="1799" externalid="372281">
              <RESULTS>
                <RESULT eventid="1084" points="466" swimtime="00:02:11.55" resultid="1800" heatid="2266" lane="2" entrytime="00:02:09.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="542" swimtime="00:00:57.45" resultid="1801" heatid="2314" lane="2" entrytime="00:00:56.51" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="De Czarnecki" birthdate="2008-06-24" gender="M" nation="BRA" license="329641" swrid="5600146" athleteid="1499" externalid="329641">
              <RESULTS>
                <RESULT eventid="1116" points="570" reactiontime="+65" swimtime="00:01:02.22" resultid="1500" heatid="2282" lane="4" entrytime="00:01:01.63" entrycourse="LCM" />
                <RESULT eventid="1084" points="504" swimtime="00:02:08.17" resultid="1501" heatid="2266" lane="3" entrytime="00:02:07.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="573" reactiontime="+69" swimtime="00:02:14.73" resultid="1502" heatid="2339" lane="4" entrytime="00:02:13.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Estela" lastname="Albuquerque" birthdate="2010-11-23" gender="F" nation="BRA" license="356344" swrid="5653285" athleteid="1619" externalid="356344">
              <RESULTS>
                <RESULT eventid="1108" points="373" reactiontime="+69" swimtime="00:01:19.61" resultid="1620" heatid="2275" lane="3" entrytime="00:01:19.04" entrycourse="LCM" />
                <RESULT eventid="1076" points="448" swimtime="00:02:27.40" resultid="1621" heatid="2254" lane="2" entrytime="00:02:32.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="346" reactiontime="+70" swimtime="00:02:55.35" resultid="1622" heatid="2334" lane="4" entrytime="00:02:53.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="420" swimtime="00:01:09.04" resultid="1623" heatid="2300" lane="2" entrytime="00:01:09.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Germer Munhoz" birthdate="2010-04-23" gender="F" nation="BRA" license="356632" swrid="5588722" athleteid="1650" externalid="356632">
              <RESULTS>
                <RESULT eventid="1124" points="309" swimtime="00:01:34.76" resultid="1651" heatid="2285" lane="7" entrytime="00:01:37.06" entrycourse="LCM" />
                <RESULT eventid="1092" points="353" swimtime="00:02:52.30" resultid="1652" heatid="2268" lane="3" entrytime="00:02:55.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1076" points="491" swimtime="00:02:22.95" resultid="1653" heatid="2255" lane="1" entrytime="00:02:25.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="360" swimtime="00:01:17.97" resultid="1654" heatid="2343" lane="7" entrytime="00:01:16.66" entrycourse="LCM" />
                <RESULT eventid="1172" points="489" swimtime="00:10:14.94" resultid="1655" heatid="2327" lane="3" entrytime="00:10:16.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.16" />
                    <SPLIT distance="200" swimtime="00:02:30.44" />
                    <SPLIT distance="300" swimtime="00:03:47.91" />
                    <SPLIT distance="400" swimtime="00:05:05.48" />
                    <SPLIT distance="500" swimtime="00:06:23.33" />
                    <SPLIT distance="600" swimtime="00:07:40.65" />
                    <SPLIT distance="700" swimtime="00:08:59.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Heloisa Souza" birthdate="2007-01-15" gender="F" nation="BRA" license="336615" swrid="5600184" athleteid="1531" externalid="336615">
              <RESULTS>
                <RESULT eventid="1076" points="635" swimtime="00:02:11.27" resultid="1532" heatid="2256" lane="4" entrytime="00:02:11.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="577" swimtime="00:09:42.00" resultid="1533" heatid="2326" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.26" />
                    <SPLIT distance="200" swimtime="00:02:22.51" />
                    <SPLIT distance="300" swimtime="00:03:34.59" />
                    <SPLIT distance="400" swimtime="00:04:47.97" />
                    <SPLIT distance="500" swimtime="00:06:01.58" />
                    <SPLIT distance="600" swimtime="00:07:15.93" />
                    <SPLIT distance="700" swimtime="00:08:31.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="609" swimtime="00:01:00.99" resultid="1534" heatid="2302" lane="4" entrytime="00:01:00.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Iglesias Vargas" birthdate="2009-01-11" gender="M" nation="BRA" license="324792" swrid="5600189" athleteid="1528" externalid="324792">
              <RESULTS>
                <RESULT eventid="1084" points="529" swimtime="00:02:06.10" resultid="1529" heatid="2266" lane="6" entrytime="00:02:07.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="494" swimtime="00:09:31.85" resultid="1530" heatid="2331" lane="5" entrytime="00:09:26.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.55" />
                    <SPLIT distance="200" swimtime="00:02:16.34" />
                    <SPLIT distance="300" swimtime="00:03:27.67" />
                    <SPLIT distance="400" swimtime="00:04:39.66" />
                    <SPLIT distance="500" swimtime="00:05:51.47" />
                    <SPLIT distance="600" swimtime="00:07:05.57" />
                    <SPLIT distance="700" swimtime="00:08:19.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariana" lastname="Stoberl" birthdate="2010-07-09" gender="F" nation="BRA" license="356250" swrid="5600265" athleteid="1608" externalid="356250">
              <RESULTS>
                <RESULT eventid="1076" points="513" swimtime="00:02:20.94" resultid="1609" heatid="2255" lane="5" entrytime="00:02:23.42" entrycourse="LCM" />
                <RESULT eventid="1204" status="DSQ" swimtime="00:01:19.34" resultid="1610" heatid="2340" lane="3" />
                <RESULT eventid="1188" points="406" reactiontime="+71" swimtime="00:02:46.19" resultid="1611" heatid="2335" lane="7" entrytime="00:02:47.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="526" swimtime="00:01:04.05" resultid="1612" heatid="2301" lane="5" entrytime="00:01:05.78" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivia" lastname="Jeger" birthdate="2004-12-19" gender="F" nation="BRA" license="325493" swrid="5600193" athleteid="1819" externalid="325493" level="UNIDOMBOSC">
              <RESULTS>
                <RESULT eventid="1092" points="496" swimtime="00:02:33.84" resultid="1820" heatid="2268" lane="5" entrytime="00:02:31.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="532" swimtime="00:05:27.96" resultid="1821" heatid="2246" lane="4" entrytime="00:05:19.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.68" />
                    <SPLIT distance="200" swimtime="00:02:37.92" />
                    <SPLIT distance="300" swimtime="00:04:15.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="549" swimtime="00:01:03.14" resultid="1822" heatid="2302" lane="2" entrytime="00:01:03.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Cury" birthdate="2005-09-28" gender="M" nation="BRA" license="329251" swrid="5600270" athleteid="1671" externalid="329251" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1100" points="614" swimtime="00:02:09.82" resultid="1672" heatid="2270" lane="5" entrytime="00:02:10.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="645" swimtime="00:00:57.21" resultid="1673" heatid="2350" lane="3" entrytime="00:00:57.67" entrycourse="LCM" />
                <RESULT eventid="1148" points="581" swimtime="00:00:56.14" resultid="1674" heatid="2315" lane="7" entrytime="00:00:53.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo" lastname="Gabriel Nascimento" birthdate="2008-11-14" gender="M" nation="BRA" license="348028" swrid="5600171" athleteid="1816" externalid="348028" level="BIG BUM">
              <RESULTS>
                <RESULT eventid="1100" status="DSQ" swimtime="00:02:45.83" resultid="1817" heatid="2270" lane="8" entrytime="00:02:48.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="445" swimtime="00:01:04.76" resultid="1818" heatid="2349" lane="1" entrytime="00:01:04.11" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Saboia" birthdate="2009-01-25" gender="M" nation="BRA" license="342252" swrid="5600253" athleteid="1573" externalid="342252">
              <RESULTS>
                <RESULT eventid="1132" points="424" swimtime="00:01:15.70" resultid="1574" heatid="2294" lane="2" entrytime="00:01:19.33" entrycourse="LCM" />
                <RESULT eventid="1164" points="420" swimtime="00:02:47.53" resultid="1575" heatid="2323" lane="3" entrytime="00:02:53.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ferreira Motta" birthdate="2008-10-24" gender="M" nation="BRA" license="378068" swrid="5600160" athleteid="1790" externalid="378068">
              <RESULTS>
                <RESULT eventid="1132" points="425" swimtime="00:01:15.60" resultid="1791" heatid="2294" lane="3" entrytime="00:01:17.45" entrycourse="LCM" />
                <RESULT eventid="1164" points="427" swimtime="00:02:46.54" resultid="1792" heatid="2323" lane="4" entrytime="00:02:51.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Peret Saboia" birthdate="2009-11-25" gender="F" nation="BRA" license="342238" swrid="5600234" athleteid="1567" externalid="342238">
              <RESULTS>
                <RESULT eventid="1124" points="478" swimtime="00:01:21.98" resultid="1568" heatid="2287" lane="8" entrytime="00:01:22.94" entrycourse="LCM" />
                <RESULT eventid="1156" points="423" swimtime="00:03:03.13" resultid="1569" heatid="2319" lane="4" entrytime="00:03:03.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Cristina Ferreira" birthdate="2011-08-24" gender="F" nation="BRA" license="358334" swrid="5588611" athleteid="1776" externalid="358334">
              <RESULTS>
                <RESULT eventid="1092" points="537" swimtime="00:02:29.80" resultid="1777" heatid="2268" lane="4" entrytime="00:02:27.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="571" swimtime="00:05:20.44" resultid="1778" heatid="2246" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.62" />
                    <SPLIT distance="200" swimtime="00:02:37.15" />
                    <SPLIT distance="300" swimtime="00:04:09.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="604" swimtime="00:01:05.61" resultid="1779" heatid="2343" lane="5" entrytime="00:01:04.99" entrycourse="LCM" />
                <RESULT eventid="1156" points="490" swimtime="00:02:54.46" resultid="1780" heatid="2317" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diego" lastname="Rafael Faria Vellozo" birthdate="2008-02-21" gender="M" nation="BRA" license="342231" swrid="5600239" athleteid="1558" externalid="342231">
              <RESULTS>
                <RESULT eventid="1116" points="438" reactiontime="+64" swimtime="00:01:07.92" resultid="1559" heatid="2282" lane="8" entrytime="00:01:07.94" entrycourse="LCM" />
                <RESULT eventid="1196" points="408" reactiontime="+64" swimtime="00:02:30.85" resultid="1560" heatid="2338" lane="7" entrytime="00:02:34.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Martinez Diniz" birthdate="2008-11-22" gender="M" nation="BRA" license="339400" swrid="5717283" athleteid="1859" externalid="339400">
              <RESULTS>
                <RESULT eventid="1084" points="433" swimtime="00:02:14.73" resultid="1860" heatid="2260" lane="4" />
                <RESULT eventid="1180" points="374" swimtime="00:10:27.37" resultid="1861" heatid="2328" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.71" />
                    <SPLIT distance="200" swimtime="00:02:32.22" />
                    <SPLIT distance="300" swimtime="00:03:53.36" />
                    <SPLIT distance="400" swimtime="00:05:14.00" />
                    <SPLIT distance="500" swimtime="00:06:34.21" />
                    <SPLIT distance="600" swimtime="00:07:53.24" />
                    <SPLIT distance="700" swimtime="00:09:11.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Prosdocimo" birthdate="2010-11-23" gender="F" nation="BRA" license="356251" swrid="5600238" athleteid="1613" externalid="356251">
              <RESULTS>
                <RESULT eventid="1108" points="411" reactiontime="+71" swimtime="00:01:17.08" resultid="1614" heatid="2275" lane="5" entrytime="00:01:16.78" entrycourse="LCM" />
                <RESULT eventid="1076" points="489" swimtime="00:02:23.22" resultid="1615" heatid="2255" lane="2" entrytime="00:02:24.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" status="DSQ" swimtime="00:02:53.37" resultid="1616" heatid="2335" lane="1" entrytime="00:02:48.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="432" swimtime="00:10:41.28" resultid="1617" heatid="2327" lane="6" entrytime="00:10:34.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.81" />
                    <SPLIT distance="200" swimtime="00:02:35.14" />
                    <SPLIT distance="300" swimtime="00:03:56.95" />
                    <SPLIT distance="400" swimtime="00:05:19.07" />
                    <SPLIT distance="500" swimtime="00:06:41.01" />
                    <SPLIT distance="600" swimtime="00:08:03.49" />
                    <SPLIT distance="700" swimtime="00:09:25.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="463" swimtime="00:01:06.84" resultid="1618" heatid="2300" lane="4" entrytime="00:01:07.41" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Severo" lastname="Berger Leal" birthdate="2008-08-05" gender="M" nation="BRA" license="330073" swrid="5449277" athleteid="1555" externalid="330073">
              <RESULTS>
                <RESULT eventid="1132" status="DNS" swimtime="00:00:00.00" resultid="1556" heatid="2294" lane="4" entrytime="00:01:17.01" entrycourse="LCM" />
                <RESULT eventid="1164" status="DNS" swimtime="00:00:00.00" resultid="1557" heatid="2324" lane="8" entrytime="00:02:51.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Magalhaes Dos Reis" birthdate="2010-05-05" gender="M" nation="BRA" license="356361" swrid="5600207" athleteid="1644" externalid="356361">
              <RESULTS>
                <RESULT eventid="1132" points="331" swimtime="00:01:22.21" resultid="1645" heatid="2294" lane="8" entrytime="00:01:21.07" entrycourse="LCM" />
                <RESULT eventid="1084" points="377" swimtime="00:02:21.15" resultid="1646" heatid="2264" lane="7" entrytime="00:02:20.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="269" swimtime="00:01:16.51" resultid="1647" heatid="2347" lane="3" entrytime="00:01:18.89" entrycourse="LCM" />
                <RESULT eventid="1164" points="347" swimtime="00:02:58.52" resultid="1648" heatid="2323" lane="6" entrytime="00:02:56.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="463" swimtime="00:01:00.56" resultid="1649" heatid="2312" lane="2" entrytime="00:01:01.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Braun Prado" birthdate="2008-04-07" gender="M" nation="BRA" license="307663" swrid="5484324" athleteid="1586" externalid="307663">
              <RESULTS>
                <RESULT eventid="1116" points="526" reactiontime="+65" swimtime="00:01:03.92" resultid="1587" heatid="2282" lane="2" entrytime="00:01:03.74" entrycourse="LCM" />
                <RESULT eventid="1196" points="505" reactiontime="+61" swimtime="00:02:20.50" resultid="1588" heatid="2339" lane="7" entrytime="00:02:19.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Martynychen" birthdate="2011-12-19" gender="M" nation="BRA" license="366893" swrid="5602557" athleteid="1691" externalid="366893">
              <RESULTS>
                <RESULT eventid="1116" points="253" reactiontime="+31" swimtime="00:01:21.50" resultid="1692" heatid="2280" lane="7" entrytime="00:01:22.84" entrycourse="LCM" />
                <RESULT eventid="1084" points="330" swimtime="00:02:27.52" resultid="1693" heatid="2263" lane="1" entrytime="00:02:31.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="288" swimtime="00:02:49.35" resultid="1694" heatid="2337" lane="1" entrytime="00:02:56.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="366" swimtime="00:10:31.87" resultid="1695" heatid="2328" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.59" />
                    <SPLIT distance="200" swimtime="00:02:34.45" />
                    <SPLIT distance="300" swimtime="00:03:55.07" />
                    <SPLIT distance="400" swimtime="00:05:16.83" />
                    <SPLIT distance="500" swimtime="00:06:36.81" />
                    <SPLIT distance="600" swimtime="00:07:57.31" />
                    <SPLIT distance="700" swimtime="00:09:17.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Pedro Pasqual" birthdate="2009-06-17" gender="M" nation="BRA" license="386136" swrid="5600232" athleteid="1852" externalid="386136">
              <RESULTS>
                <RESULT eventid="1116" points="509" reactiontime="+63" swimtime="00:01:04.59" resultid="1853" heatid="2282" lane="7" entrytime="00:01:03.74" entrycourse="LCM" />
                <RESULT eventid="1196" points="499" reactiontime="+72" swimtime="00:02:21.08" resultid="1854" heatid="2339" lane="2" entrytime="00:02:19.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nina" lastname="Rocha Ribeiro Da Silva" birthdate="2010-09-22" gender="F" nation="BRA" license="367216" swrid="5588884" athleteid="1802" externalid="367216">
              <RESULTS>
                <RESULT eventid="1124" points="444" swimtime="00:01:24.06" resultid="1803" heatid="2286" lane="4" entrytime="00:01:23.50" entrycourse="LCM" />
                <RESULT eventid="1076" points="407" swimtime="00:02:32.21" resultid="1804" heatid="2253" lane="1" entrytime="00:02:38.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="381" swimtime="00:03:09.65" resultid="1805" heatid="2320" lane="8" entrytime="00:03:03.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="406" swimtime="00:01:09.78" resultid="1806" heatid="2299" lane="4" entrytime="00:01:10.67" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Guimaraes E Souza" birthdate="2008-12-21" gender="M" nation="BRA" license="376972" swrid="5600182" athleteid="1781" externalid="376972">
              <RESULTS>
                <RESULT eventid="1132" points="444" swimtime="00:01:14.52" resultid="1782" heatid="2295" lane="1" entrytime="00:01:12.45" entrycourse="LCM" />
                <RESULT eventid="1164" points="399" swimtime="00:02:50.37" resultid="1783" heatid="2324" lane="7" entrytime="00:02:41.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Rocha" birthdate="2011-08-25" gender="F" nation="BRA" license="366904" swrid="5602578" athleteid="1723" externalid="366904">
              <RESULTS>
                <RESULT eventid="1108" points="375" reactiontime="+54" swimtime="00:01:19.49" resultid="1724" heatid="2275" lane="8" entrytime="00:01:21.95" entrycourse="LCM" />
                <RESULT eventid="1076" points="459" swimtime="00:02:26.29" resultid="1725" heatid="2253" lane="3" entrytime="00:02:34.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="365" reactiontime="+71" swimtime="00:02:52.22" resultid="1726" heatid="2334" lane="3" entrytime="00:02:57.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:23.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="387" swimtime="00:11:05.13" resultid="1727" heatid="2325" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.75" />
                    <SPLIT distance="200" swimtime="00:02:45.94" />
                    <SPLIT distance="300" swimtime="00:04:11.98" />
                    <SPLIT distance="400" swimtime="00:05:37.99" />
                    <SPLIT distance="500" swimtime="00:07:03.43" />
                    <SPLIT distance="600" swimtime="00:08:27.64" />
                    <SPLIT distance="700" swimtime="00:09:51.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="436" swimtime="00:01:08.15" resultid="1728" heatid="2301" lane="1" entrytime="00:01:07.33" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Trevisan" birthdate="2000-11-28" gender="M" nation="BRA" license="346847" swrid="5600266" athleteid="1807" externalid="346847">
              <RESULTS>
                <RESULT eventid="1084" points="505" swimtime="00:02:08.01" resultid="1808" heatid="2266" lane="4" entrytime="00:02:05.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="470" swimtime="00:01:03.57" resultid="1809" heatid="2350" lane="8" entrytime="00:01:01.04" entrycourse="LCM" />
                <RESULT eventid="1148" points="602" swimtime="00:00:55.49" resultid="1810" heatid="2315" lane="8" entrytime="00:00:54.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Vitoria Kuzmann Cercal" birthdate="2009-04-10" gender="F" nation="BRA" license="339082" swrid="5600274" athleteid="1576" externalid="339082">
              <RESULTS>
                <RESULT eventid="1076" points="506" swimtime="00:02:21.61" resultid="1577" heatid="2256" lane="8" entrytime="00:02:22.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="401" swimtime="00:02:46.94" resultid="1578" heatid="2333" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinícius" lastname="Oliveira Cruz" birthdate="2005-07-02" gender="M" nation="BRA" license="298495" swrid="5653299" athleteid="1845" externalid="298495" level="ADTRISC">
              <RESULTS>
                <RESULT eventid="1084" points="737" swimtime="00:01:52.89" resultid="1846" heatid="2267" lane="4" entrytime="00:01:51.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:55.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="554" swimtime="00:01:00.18" resultid="1847" heatid="2350" lane="6" entrytime="00:00:58.17" entrycourse="LCM" />
                <RESULT eventid="1148" points="723" swimtime="00:00:52.19" resultid="1848" heatid="2315" lane="5" entrytime="00:00:51.56" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Fontes Hoshina" birthdate="2008-02-15" gender="M" nation="BRA" license="369445" swrid="5600165" athleteid="1507" externalid="369445">
              <RESULTS>
                <RESULT eventid="1100" status="DNS" swimtime="00:00:00.00" resultid="1508" heatid="2269" lane="7" />
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="1509" heatid="2350" lane="1" entrytime="00:01:00.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16131" nation="BRA" region="PR" clubid="1873" swrid="93766" name="Associação Nadar Colombo" shortname="Equipe Nadar">
          <ATHLETES>
            <ATHLETE firstname="Eduardo" lastname="Luiz Sartori" birthdate="2008-04-07" gender="M" nation="BRA" license="384742" swrid="5622287" athleteid="1885" externalid="384742">
              <RESULTS>
                <RESULT eventid="1084" points="400" swimtime="00:02:18.39" resultid="1886" heatid="2264" lane="8" entrytime="00:02:23.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="341" reactiontime="+80" swimtime="00:02:40.11" resultid="1887" heatid="2337" lane="3" entrytime="00:02:44.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Rafael D Agostin Batistao" birthdate="2008-05-13" gender="M" nation="BRA" license="384738" swrid="5622300" athleteid="1874" externalid="384738">
              <RESULTS>
                <RESULT eventid="1132" points="323" swimtime="00:01:22.87" resultid="1875" heatid="2293" lane="5" entrytime="00:01:22.96" entrycourse="LCM" />
                <RESULT eventid="1148" points="344" swimtime="00:01:06.87" resultid="1876" heatid="2310" lane="7" entrytime="00:01:06.86" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Krik" birthdate="2010-11-24" gender="F" nation="BRA" license="406702" swrid="5717277" athleteid="1896" externalid="406702">
              <RESULTS>
                <RESULT eventid="1124" points="134" swimtime="00:02:05.08" resultid="1897" heatid="2283" lane="3" />
                <RESULT eventid="1140" points="144" swimtime="00:01:38.60" resultid="1898" heatid="2297" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Felipe Glir" birthdate="2006-10-11" gender="M" nation="BRA" license="384741" swrid="5622280" athleteid="1882" externalid="384741">
              <RESULTS>
                <RESULT eventid="1212" status="DNS" swimtime="00:00:00.00" resultid="1883" heatid="2346" lane="7" />
                <RESULT eventid="1148" points="392" swimtime="00:01:04.01" resultid="1884" heatid="2312" lane="1" entrytime="00:01:02.26" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaylaine" lastname="Sofia Vargas Bueno" birthdate="2006-11-28" gender="F" nation="BRA" license="384739" swrid="5622307" athleteid="1877" externalid="384739">
              <RESULTS>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="1878" heatid="2284" lane="5" entrytime="00:01:42.66" entrycourse="LCM" />
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="1879" heatid="2251" lane="5" entrytime="00:02:57.14" entrycourse="LCM" />
                <RESULT eventid="1156" points="221" swimtime="00:03:47.28" resultid="1880" heatid="2317" lane="4" entrytime="00:03:45.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:50.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="304" swimtime="00:01:16.85" resultid="1881" heatid="2298" lane="3" entrytime="00:01:18.21" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Rosa De Souza" birthdate="2009-01-01" gender="F" nation="BRA" license="399926" swrid="5653301" athleteid="1888" externalid="399926">
              <RESULTS>
                <RESULT eventid="1124" points="221" swimtime="00:01:46.07" resultid="1889" heatid="2284" lane="3" entrytime="00:01:46.82" entrycourse="LCM" />
                <RESULT eventid="1204" points="104" swimtime="00:01:57.81" resultid="1890" heatid="2341" lane="8" />
                <RESULT eventid="1172" points="210" swimtime="00:13:34.50" resultid="1891" heatid="2326" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.45" />
                    <SPLIT distance="200" swimtime="00:03:18.68" />
                    <SPLIT distance="300" swimtime="00:05:04.14" />
                    <SPLIT distance="400" swimtime="00:06:48.98" />
                    <SPLIT distance="500" swimtime="00:08:33.90" />
                    <SPLIT distance="600" swimtime="00:10:19.59" />
                    <SPLIT distance="700" swimtime="00:12:00.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Carvalho" birthdate="2011-10-20" gender="F" nation="BRA" license="399927" swrid="5652882" athleteid="1892" externalid="399927">
              <RESULTS>
                <RESULT eventid="1124" points="241" swimtime="00:01:43.02" resultid="1893" heatid="2283" lane="2" />
                <RESULT eventid="1204" points="144" swimtime="00:01:45.68" resultid="1894" heatid="2340" lane="4" />
                <RESULT eventid="1140" points="265" swimtime="00:01:20.49" resultid="1895" heatid="2298" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2864" nation="BRA" region="PR" clubid="1221" swrid="93756" name="Associacao De Pais E Amigos Da Natacao De Ponta Gr" shortname="Apan Ponta Grossa">
          <ATHLETES>
            <ATHLETE firstname="Yoseph" lastname="Rigoni Moraes" birthdate="2006-04-17" gender="M" nation="BRA" license="295182" swrid="5622302" athleteid="1262" externalid="295182" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1132" points="431" swimtime="00:01:15.29" resultid="1263" heatid="2291" lane="7" />
                <RESULT eventid="1212" points="376" swimtime="00:01:08.51" resultid="1264" heatid="2344" lane="4" />
                <RESULT eventid="1148" points="466" swimtime="00:01:00.42" resultid="1265" heatid="2313" lane="7" entrytime="00:00:59.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fegert" birthdate="2009-04-13" gender="M" nation="BRA" license="353813" swrid="5622279" athleteid="1255" externalid="353813">
              <RESULTS>
                <RESULT eventid="1212" points="349" swimtime="00:01:10.21" resultid="1256" heatid="2344" lane="6" />
                <RESULT eventid="1148" points="446" swimtime="00:01:01.32" resultid="1257" heatid="2306" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Dolinski Thomassewski" birthdate="2006-12-15" gender="M" nation="BRA" license="400409" swrid="5653289" athleteid="1281" externalid="400409">
              <RESULTS>
                <RESULT eventid="1132" points="249" swimtime="00:01:30.30" resultid="1282" heatid="2292" lane="6" entrytime="00:01:35.57" entrycourse="LCM" />
                <RESULT eventid="1148" points="280" swimtime="00:01:11.60" resultid="1283" heatid="2308" lane="1" entrytime="00:01:16.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Campagnoli" birthdate="2009-04-13" gender="F" nation="BRA" license="366915" swrid="5600128" athleteid="1243" externalid="366915">
              <RESULTS>
                <RESULT eventid="1108" points="451" swimtime="00:01:14.74" resultid="1244" heatid="2276" lane="1" entrytime="00:01:15.12" entrycourse="LCM" />
                <RESULT eventid="1076" points="529" swimtime="00:02:19.52" resultid="1245" heatid="2254" lane="6" entrytime="00:02:31.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="436" reactiontime="+74" swimtime="00:02:42.35" resultid="1246" heatid="2335" lane="6" entrytime="00:02:42.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="508" swimtime="00:01:04.80" resultid="1247" heatid="2300" lane="6" entrytime="00:01:08.54" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Renato" lastname="Mandalozzo Tebcherani" birthdate="2004-03-16" gender="M" nation="BRA" license="279221" swrid="5622290" athleteid="1236" externalid="279221" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1132" points="407" swimtime="00:01:16.73" resultid="1237" heatid="2294" lane="5" entrytime="00:01:17.16" entrycourse="LCM" />
                <RESULT eventid="1148" points="421" swimtime="00:01:02.52" resultid="1238" heatid="2303" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Augusto" lastname="Tramontin" birthdate="2011-11-29" gender="M" nation="BRA" license="399691" swrid="5652901" athleteid="1266" externalid="399691">
              <RESULTS>
                <RESULT eventid="1132" points="236" swimtime="00:01:31.92" resultid="1267" heatid="2292" lane="7" entrytime="00:01:40.68" entrycourse="LCM" />
                <RESULT eventid="1116" points="285" reactiontime="+79" swimtime="00:01:18.33" resultid="1268" heatid="2277" lane="7" />
                <RESULT eventid="1148" points="299" swimtime="00:01:10.07" resultid="1269" heatid="2308" lane="7" entrytime="00:01:13.26" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Franca Berger" birthdate="2010-05-07" gender="F" nation="BRA" license="399692" swrid="5653290" athleteid="1270" externalid="399692">
              <RESULTS>
                <RESULT eventid="1124" points="231" swimtime="00:01:44.45" resultid="1271" heatid="2284" lane="2" entrytime="00:01:57.23" entrycourse="LCM" />
                <RESULT eventid="1156" points="200" swimtime="00:03:55.04" resultid="1272" heatid="2317" lane="3" entrytime="00:04:23.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:55.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="256" swimtime="00:01:21.34" resultid="1273" heatid="2298" lane="2" entrytime="00:01:25.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Mandalozzo Tebcherani" birthdate="2006-03-02" gender="M" nation="BRA" license="295181" swrid="5622289" athleteid="1274" externalid="295181" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1132" points="299" swimtime="00:01:25.05" resultid="1275" heatid="2289" lane="5" />
                <RESULT eventid="1148" points="381" swimtime="00:01:04.61" resultid="1276" heatid="2304" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Allana" lastname="Lacerda" birthdate="2005-03-15" gender="F" nation="BRA" license="295186" swrid="5600197" athleteid="1239" externalid="295186" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1124" points="408" swimtime="00:01:26.45" resultid="1240" heatid="2287" lane="1" entrytime="00:01:22.04" entrycourse="LCM" />
                <RESULT eventid="1204" points="312" swimtime="00:01:21.77" resultid="1241" heatid="2342" lane="5" entrytime="00:01:20.90" entrycourse="LCM" />
                <RESULT eventid="1156" points="420" swimtime="00:03:03.57" resultid="1242" heatid="2320" lane="7" entrytime="00:02:58.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:30.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Chi Kravchychyn" birthdate="2009-09-27" gender="M" nation="BRA" license="344268" swrid="5600134" athleteid="1227" externalid="344268">
              <RESULTS>
                <RESULT eventid="1132" points="497" swimtime="00:01:11.77" resultid="1228" heatid="2295" lane="6" entrytime="00:01:09.95" entrycourse="LCM" />
                <RESULT eventid="1100" points="457" swimtime="00:02:23.22" resultid="1229" heatid="2270" lane="3" entrytime="00:02:16.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="520" swimtime="00:05:01.46" resultid="1230" heatid="2248" lane="5" entrytime="00:04:51.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.69" />
                    <SPLIT distance="200" swimtime="00:02:26.13" />
                    <SPLIT distance="300" swimtime="00:03:52.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="481" swimtime="00:01:03.10" resultid="1231" heatid="2349" lane="2" entrytime="00:01:02.93" entrycourse="LCM" />
                <RESULT eventid="1164" points="520" swimtime="00:02:35.99" resultid="1232" heatid="2324" lane="5" entrytime="00:02:31.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yohan" lastname="Rigoni Moraes" birthdate="2002-04-03" gender="M" nation="BRA" license="272187" swrid="5600245" athleteid="1233" externalid="272187" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1132" points="596" swimtime="00:01:07.58" resultid="1234" heatid="2295" lane="3" entrytime="00:01:07.80" entrycourse="LCM" />
                <RESULT eventid="1164" points="520" swimtime="00:02:35.96" resultid="1235" heatid="2324" lane="6" entrytime="00:02:37.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Carolina Babiuki" birthdate="2007-02-06" gender="F" nation="BRA" license="316227" swrid="5600131" athleteid="1248" externalid="316227" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1108" points="452" reactiontime="+64" swimtime="00:01:14.67" resultid="1249" heatid="2276" lane="7" entrytime="00:01:12.40" entrycourse="LCM" />
                <RESULT eventid="1188" points="440" reactiontime="+68" swimtime="00:02:41.85" resultid="1250" heatid="2335" lane="3" entrytime="00:02:40.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="495" swimtime="00:01:05.33" resultid="1251" heatid="2302" lane="1" entrytime="00:01:04.18" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Delinski" birthdate="2009-11-28" gender="F" nation="BRA" license="385190" swrid="5600150" athleteid="1252" externalid="385190">
              <RESULTS>
                <RESULT eventid="1108" points="321" reactiontime="+84" swimtime="00:01:23.70" resultid="1253" heatid="2271" lane="5" />
                <RESULT eventid="1156" points="316" swimtime="00:03:21.86" resultid="1254" heatid="2318" lane="3" entrytime="00:03:27.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Gueiber Montes" birthdate="2009-03-09" gender="M" nation="BRA" license="342154" swrid="5600179" athleteid="1222" externalid="342154">
              <RESULTS>
                <RESULT eventid="1116" points="550" reactiontime="+62" swimtime="00:01:02.97" resultid="1223" heatid="2282" lane="3" entrytime="00:01:01.79" entrycourse="LCM" />
                <RESULT eventid="1084" points="551" swimtime="00:02:04.41" resultid="1224" heatid="2267" lane="8" entrytime="00:02:04.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:59.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="471" reactiontime="+63" swimtime="00:02:23.75" resultid="1225" heatid="2339" lane="6" entrytime="00:02:19.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="586" swimtime="00:00:55.98" resultid="1226" heatid="2314" lane="7" entrytime="00:00:57.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Sabedotti" birthdate="2011-04-20" gender="F" nation="BRA" license="390877" swrid="5602580" athleteid="1277" externalid="390877">
              <RESULTS>
                <RESULT eventid="1108" points="369" reactiontime="+74" swimtime="00:01:19.92" resultid="1278" heatid="2274" lane="4" entrytime="00:01:22.12" entrycourse="LCM" />
                <RESULT eventid="1188" points="333" reactiontime="+69" swimtime="00:02:57.64" resultid="1279" heatid="2332" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="417" swimtime="00:01:09.20" resultid="1280" heatid="2297" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Carraro Borges" birthdate="2009-05-11" gender="M" nation="BRA" license="345590" swrid="5622267" athleteid="1258" externalid="345590" level="SAGRADA FA">
              <RESULTS>
                <RESULT eventid="1084" points="422" swimtime="00:02:15.97" resultid="1259" heatid="2264" lane="5" entrytime="00:02:18.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="424" swimtime="00:10:01.46" resultid="1260" heatid="2330" lane="3" entrytime="00:10:18.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.09" />
                    <SPLIT distance="200" swimtime="00:02:22.55" />
                    <SPLIT distance="300" swimtime="00:03:37.81" />
                    <SPLIT distance="400" swimtime="00:04:54.59" />
                    <SPLIT distance="500" swimtime="00:06:10.94" />
                    <SPLIT distance="600" swimtime="00:07:28.41" />
                    <SPLIT distance="700" swimtime="00:08:46.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="397" swimtime="00:01:03.71" resultid="1261" heatid="2311" lane="1" entrytime="00:01:03.46" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13068" nation="BRA" region="PR" clubid="1941" swrid="93787" name="Sociedade Morgenau" shortname="Morgenau">
          <ATHLETES>
            <ATHLETE firstname="Bruno" lastname="Gabriel Sarmento Buski" birthdate="2010-04-05" gender="M" nation="BRA" license="399533" swrid="5717264" athleteid="1963" externalid="399533">
              <RESULTS>
                <RESULT eventid="1132" points="222" swimtime="00:01:33.87" resultid="1964" heatid="2290" lane="4" />
                <RESULT eventid="1084" points="275" swimtime="00:02:36.68" resultid="1965" heatid="2260" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="294" swimtime="00:11:19.76" resultid="1966" heatid="2329" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.07" />
                    <SPLIT distance="200" swimtime="00:02:45.45" />
                    <SPLIT distance="300" swimtime="00:04:13.48" />
                    <SPLIT distance="400" swimtime="00:05:40.65" />
                    <SPLIT distance="500" swimtime="00:07:07.54" />
                    <SPLIT distance="600" swimtime="00:08:34.38" />
                    <SPLIT distance="700" swimtime="00:09:59.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="273" swimtime="00:01:12.23" resultid="1967" heatid="2305" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="De Mello Araujo" birthdate="2010-11-03" gender="F" nation="BRA" license="406723" swrid="5717254" athleteid="2085" externalid="406723">
              <RESULTS>
                <RESULT eventid="1124" points="183" swimtime="00:01:52.84" resultid="2086" heatid="2283" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monike" lastname="Lemos Carvalho" birthdate="2008-03-28" gender="F" nation="BRA" license="307796" swrid="5600199" athleteid="2015" externalid="307796">
              <RESULTS>
                <RESULT eventid="1108" points="404" reactiontime="+69" swimtime="00:01:17.55" resultid="2016" heatid="2275" lane="7" entrytime="00:01:19.73" entrycourse="LCM" />
                <RESULT eventid="1076" points="469" swimtime="00:02:25.21" resultid="2017" heatid="2254" lane="3" entrytime="00:02:31.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="386" swimtime="00:11:05.75" resultid="2018" heatid="2325" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.22" />
                    <SPLIT distance="200" swimtime="00:02:39.71" />
                    <SPLIT distance="300" swimtime="00:04:05.40" />
                    <SPLIT distance="400" swimtime="00:05:31.39" />
                    <SPLIT distance="500" swimtime="00:06:57.60" />
                    <SPLIT distance="600" swimtime="00:08:23.31" />
                    <SPLIT distance="700" swimtime="00:09:48.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="437" swimtime="00:01:08.11" resultid="2019" heatid="2300" lane="3" entrytime="00:01:08.33" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kedny" lastname="Correa" birthdate="2004-11-05" gender="M" nation="BRA" license="383858" swrid="5600142" athleteid="2003" externalid="383858">
              <RESULTS>
                <RESULT eventid="1100" points="251" swimtime="00:02:54.78" resultid="2004" heatid="2270" lane="1" entrytime="00:02:39.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1084" points="426" swimtime="00:02:15.54" resultid="2005" heatid="2258" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="317" swimtime="00:01:12.52" resultid="2006" heatid="2348" lane="2" entrytime="00:01:08.42" entrycourse="LCM" />
                <RESULT eventid="1180" points="440" swimtime="00:09:54.19" resultid="2007" heatid="2331" lane="8" entrytime="00:09:54.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.41" />
                    <SPLIT distance="200" swimtime="00:02:17.16" />
                    <SPLIT distance="300" swimtime="00:03:31.98" />
                    <SPLIT distance="400" swimtime="00:04:47.98" />
                    <SPLIT distance="500" swimtime="00:06:04.98" />
                    <SPLIT distance="600" swimtime="00:07:21.67" />
                    <SPLIT distance="700" swimtime="00:08:38.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Rodrigues Galvao" birthdate="2007-04-19" gender="M" nation="BRA" license="376586" swrid="5600247" athleteid="1953" externalid="376586">
              <RESULTS>
                <RESULT eventid="1100" points="324" swimtime="00:02:40.63" resultid="1954" heatid="2270" lane="2" entrytime="00:02:36.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="463" swimtime="00:01:03.91" resultid="1955" heatid="2348" lane="4" entrytime="00:01:04.73" entrycourse="LCM" />
                <RESULT eventid="1148" points="516" swimtime="00:00:58.39" resultid="1956" heatid="2313" lane="6" entrytime="00:00:59.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Bilecki" birthdate="2007-05-28" gender="M" nation="BRA" license="406726" swrid="5717247" athleteid="2087" externalid="406726">
              <RESULTS>
                <RESULT eventid="1212" points="255" swimtime="00:01:17.98" resultid="2088" heatid="2346" lane="1" />
                <RESULT eventid="1180" points="249" swimtime="00:11:58.12" resultid="2089" heatid="2330" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.49" />
                    <SPLIT distance="200" swimtime="00:02:48.60" />
                    <SPLIT distance="300" swimtime="00:04:20.31" />
                    <SPLIT distance="400" swimtime="00:05:54.42" />
                    <SPLIT distance="500" swimtime="00:07:28.53" />
                    <SPLIT distance="600" swimtime="00:09:03.59" />
                    <SPLIT distance="700" swimtime="00:10:33.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" status="DSQ" swimtime="00:00:00.00" resultid="2090" heatid="2303" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benito" lastname="Alves Sant&apos;Ana" birthdate="2009-06-01" gender="M" nation="BRA" license="376585" swrid="5351951" athleteid="1957" externalid="376585">
              <RESULTS>
                <RESULT eventid="1116" points="374" reactiontime="+84" swimtime="00:01:11.59" resultid="1958" heatid="2280" lane="4" entrytime="00:01:15.08" entrycourse="LCM" />
                <RESULT eventid="1084" points="458" swimtime="00:02:12.30" resultid="1959" heatid="2258" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:05.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1068" points="438" swimtime="00:05:19.27" resultid="1960" heatid="2248" lane="2" entrytime="00:05:30.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.60" />
                    <SPLIT distance="200" swimtime="00:02:35.89" />
                    <SPLIT distance="300" swimtime="00:04:12.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="379" reactiontime="+72" swimtime="00:02:34.63" resultid="1961" heatid="2338" lane="8" entrytime="00:02:37.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="518" swimtime="00:09:22.90" resultid="1962" heatid="2331" lane="2" entrytime="00:09:42.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.59" />
                    <SPLIT distance="200" swimtime="00:02:14.88" />
                    <SPLIT distance="300" swimtime="00:03:26.47" />
                    <SPLIT distance="400" swimtime="00:04:38.30" />
                    <SPLIT distance="500" swimtime="00:05:49.78" />
                    <SPLIT distance="600" swimtime="00:07:02.55" />
                    <SPLIT distance="700" swimtime="00:08:14.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thiago" lastname="Kozera Chiarato" birthdate="2008-01-22" gender="M" nation="BRA" license="406728" swrid="5717276" athleteid="2091" externalid="406728">
              <RESULTS>
                <RESULT eventid="1100" status="DSQ" swimtime="00:03:12.39" resultid="2092" heatid="2269" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:28.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1084" points="299" swimtime="00:02:32.45" resultid="2093" heatid="2259" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="236" swimtime="00:01:19.97" resultid="2094" heatid="2345" lane="4" />
                <RESULT eventid="1148" points="351" swimtime="00:01:06.43" resultid="2095" heatid="2303" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Fernanda Pinto" birthdate="2004-09-17" gender="F" nation="BRA" license="391144" swrid="5600157" athleteid="2035" externalid="391144">
              <RESULTS>
                <RESULT eventid="1108" points="203" reactiontime="+86" swimtime="00:01:37.45" resultid="2036" heatid="2272" lane="6" entrytime="00:01:51.11" entrycourse="LCM" />
                <RESULT eventid="1076" points="310" swimtime="00:02:46.69" resultid="2037" heatid="2251" lane="6" entrytime="00:03:03.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="199" swimtime="00:01:35.00" resultid="2038" heatid="2340" lane="6" />
                <RESULT eventid="1140" points="342" swimtime="00:01:13.88" resultid="2039" heatid="2298" lane="5" entrytime="00:01:17.91" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Capoia Soares" birthdate="2011-11-07" gender="M" nation="BRA" license="393257" swrid="5616440" athleteid="2054" externalid="393257">
              <RESULTS>
                <RESULT eventid="1212" status="DSQ" swimtime="00:02:01.65" resultid="2055" heatid="2345" lane="5" />
                <RESULT eventid="1148" points="107" swimtime="00:01:38.47" resultid="2056" heatid="2307" lane="7" entrytime="00:01:49.26" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Vitor Navarro Zanini" birthdate="2008-06-30" gender="M" nation="BRA" license="369415" swrid="5600273" athleteid="1990" externalid="369415">
              <RESULTS>
                <RESULT eventid="1132" points="317" swimtime="00:01:23.36" resultid="1991" heatid="2293" lane="2" entrytime="00:01:28.54" entrycourse="LCM" />
                <RESULT eventid="1084" points="345" swimtime="00:02:25.31" resultid="1992" heatid="2259" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="292" swimtime="00:03:08.97" resultid="1993" heatid="2322" lane="4" entrytime="00:03:12.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Portella Da Silva" birthdate="2010-07-19" gender="M" nation="BRA" license="399534" swrid="5717288" athleteid="1968" externalid="399534">
              <RESULTS>
                <RESULT eventid="1132" points="163" swimtime="00:01:43.97" resultid="1969" heatid="2289" lane="4" />
                <RESULT eventid="1084" points="185" swimtime="00:02:58.95" resultid="1970" heatid="2257" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="180" swimtime="00:01:22.89" resultid="1971" heatid="2305" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stella" lastname="Magalhaes Birnbaum" birthdate="2009-05-14" gender="F" nation="BRA" license="399684" swrid="5653298" athleteid="2065" externalid="399684">
              <RESULTS>
                <RESULT eventid="1204" points="136" swimtime="00:01:47.72" resultid="2066" heatid="2341" lane="5" />
                <RESULT eventid="1188" points="271" reactiontime="+93" swimtime="00:03:10.15" resultid="2067" heatid="2332" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="332" swimtime="00:01:14.64" resultid="2068" heatid="2299" lane="7" entrytime="00:01:14.23" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabryel" lastname="Denk" birthdate="2011-05-09" gender="M" nation="BRA" license="391138" swrid="5602531" athleteid="2022" externalid="391138">
              <RESULTS>
                <RESULT eventid="1132" points="189" swimtime="00:01:38.97" resultid="2023" heatid="2289" lane="8" />
                <RESULT eventid="1116" points="244" reactiontime="+65" swimtime="00:01:22.52" resultid="2024" heatid="2278" lane="7" />
                <RESULT eventid="1084" points="295" swimtime="00:02:33.18" resultid="2025" heatid="2261" lane="4" entrytime="00:02:50.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Yoshie Kimura" birthdate="2010-07-08" gender="F" nation="BRA" license="391142" swrid="5600277" athleteid="1972" externalid="391142">
              <RESULTS>
                <RESULT eventid="1124" points="456" swimtime="00:01:23.31" resultid="1973" heatid="2286" lane="6" entrytime="00:01:26.68" entrycourse="LCM" />
                <RESULT eventid="1172" points="334" swimtime="00:11:38.09" resultid="1974" heatid="2325" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.39" />
                    <SPLIT distance="200" swimtime="00:02:48.55" />
                    <SPLIT distance="300" swimtime="00:04:17.98" />
                    <SPLIT distance="400" swimtime="00:05:47.64" />
                    <SPLIT distance="500" swimtime="00:07:17.31" />
                    <SPLIT distance="600" swimtime="00:08:48.62" />
                    <SPLIT distance="700" swimtime="00:10:17.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="382" swimtime="00:03:09.42" resultid="1975" heatid="2319" lane="6" entrytime="00:03:08.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:29.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Kozera Chiarato" birthdate="2010-05-28" gender="M" nation="BRA" license="406722" swrid="5717275" athleteid="2080" externalid="406722">
              <RESULTS>
                <RESULT eventid="1132" points="188" swimtime="00:01:39.27" resultid="2081" heatid="2291" lane="1" />
                <RESULT eventid="1084" points="222" swimtime="00:02:48.42" resultid="2082" heatid="2259" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="193" swimtime="00:01:25.50" resultid="2083" heatid="2345" lane="8" />
                <RESULT eventid="1148" points="264" swimtime="00:01:12.98" resultid="2084" heatid="2306" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauan" lastname="Araujo" birthdate="2009-12-17" gender="M" nation="BRA" license="385119" swrid="5653286" athleteid="2008" externalid="385119">
              <RESULTS>
                <RESULT eventid="1132" points="246" swimtime="00:01:30.76" resultid="2009" heatid="2292" lane="1" entrytime="00:01:42.70" entrycourse="LCM" />
                <RESULT eventid="1084" points="347" swimtime="00:02:25.04" resultid="2010" heatid="2261" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="379" swimtime="00:01:04.73" resultid="2011" heatid="2308" lane="4" entrytime="00:01:11.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Mingorance Martins" birthdate="2007-10-13" gender="M" nation="BRA" license="393920" swrid="5622295" athleteid="2057" externalid="393920">
              <RESULTS>
                <RESULT eventid="1084" points="442" swimtime="00:02:13.84" resultid="2058" heatid="2265" lane="7" entrytime="00:02:15.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="396" swimtime="00:10:15.33" resultid="2059" heatid="2329" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.06" />
                    <SPLIT distance="200" swimtime="00:02:26.91" />
                    <SPLIT distance="300" swimtime="00:03:44.65" />
                    <SPLIT distance="400" swimtime="00:05:03.07" />
                    <SPLIT distance="500" swimtime="00:06:22.08" />
                    <SPLIT distance="600" swimtime="00:07:42.70" />
                    <SPLIT distance="700" swimtime="00:09:01.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="522" swimtime="00:00:58.19" resultid="2060" heatid="2314" lane="1" entrytime="00:00:57.58" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karine" lastname="Correa" birthdate="2002-08-01" gender="F" nation="BRA" license="385191" swrid="5600141" athleteid="2012" externalid="385191">
              <RESULTS>
                <RESULT eventid="1076" points="300" swimtime="00:02:48.45" resultid="2013" heatid="2253" lane="8" entrytime="00:02:39.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="346" swimtime="00:01:13.64" resultid="2014" heatid="2299" lane="2" entrytime="00:01:12.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduarda" lastname="Azevedo Birsneek" birthdate="2010-03-31" gender="F" nation="BRA" license="391145" swrid="5389427" athleteid="2040" externalid="391145">
              <RESULTS>
                <RESULT eventid="1108" points="203" swimtime="00:01:37.48" resultid="2041" heatid="2273" lane="1" entrytime="00:01:36.29" entrycourse="LCM" />
                <RESULT eventid="1076" points="167" swimtime="00:03:24.81" resultid="2042" heatid="2250" lane="4" entrytime="00:03:40.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="113" swimtime="00:01:54.43" resultid="2043" heatid="2342" lane="1" />
                <RESULT eventid="1188" points="192" reactiontime="+70" swimtime="00:03:33.25" resultid="2044" heatid="2333" lane="3" entrytime="00:03:39.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:45.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Andreis Ramos" birthdate="2007-03-26" gender="M" nation="BRA" license="406719" swrid="5717243" athleteid="2072" externalid="406719">
              <RESULTS>
                <RESULT eventid="1084" points="262" swimtime="00:02:39.25" resultid="2073" heatid="2260" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="363" swimtime="00:01:05.69" resultid="2074" heatid="2303" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauren" lastname="Dziura" birthdate="2010-01-11" gender="F" nation="BRA" license="369416" swrid="5588668" athleteid="1994" externalid="369416">
              <RESULTS>
                <RESULT eventid="1108" points="295" reactiontime="+70" swimtime="00:01:26.04" resultid="1995" heatid="2274" lane="7" entrytime="00:01:24.45" entrycourse="LCM" />
                <RESULT eventid="1076" points="386" swimtime="00:02:34.94" resultid="1996" heatid="2252" lane="5" entrytime="00:02:42.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="374" swimtime="00:11:12.46" resultid="1997" heatid="2326" lane="5" entrytime="00:11:52.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.68" />
                    <SPLIT distance="200" swimtime="00:02:40.73" />
                    <SPLIT distance="300" swimtime="00:04:04.18" />
                    <SPLIT distance="400" swimtime="00:05:30.77" />
                    <SPLIT distance="500" swimtime="00:06:56.81" />
                    <SPLIT distance="600" swimtime="00:08:23.76" />
                    <SPLIT distance="700" swimtime="00:09:49.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="358" swimtime="00:01:12.76" resultid="1998" heatid="2299" lane="6" entrytime="00:01:12.13" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Luiz Fischer" birthdate="2009-06-07" gender="M" nation="BRA" license="400273" swrid="5653296" athleteid="2069" externalid="400273">
              <RESULTS>
                <RESULT eventid="1212" points="186" swimtime="00:01:26.50" resultid="2070" heatid="2347" lane="1" entrytime="00:01:25.84" entrycourse="LCM" />
                <RESULT eventid="1148" points="214" swimtime="00:01:18.33" resultid="2071" heatid="2307" lane="3" entrytime="00:01:19.63" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Lima" birthdate="2006-12-03" gender="M" nation="BRA" license="366749" swrid="5600201" athleteid="1999" externalid="366749">
              <RESULTS>
                <RESULT eventid="1084" points="517" swimtime="00:02:07.03" resultid="2000" heatid="2267" lane="1" entrytime="00:02:03.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:00.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="462" swimtime="00:01:03.94" resultid="2001" heatid="2349" lane="6" entrytime="00:01:02.90" entrycourse="LCM" />
                <RESULT eventid="1148" points="578" swimtime="00:00:56.25" resultid="2002" heatid="2314" lane="6" entrytime="00:00:55.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Liz Skowronski" birthdate="2008-01-24" gender="F" nation="BRA" license="358245" swrid="5600202" athleteid="1948" externalid="358245">
              <RESULTS>
                <RESULT eventid="1108" points="369" reactiontime="+66" swimtime="00:01:19.87" resultid="1949" heatid="2275" lane="2" entrytime="00:01:19.52" entrycourse="LCM" />
                <RESULT eventid="1076" points="408" swimtime="00:02:32.10" resultid="1950" heatid="2249" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="348" reactiontime="+67" swimtime="00:02:54.94" resultid="1951" heatid="2335" lane="8" entrytime="00:02:49.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1172" points="372" swimtime="00:11:13.77" resultid="1952" heatid="2327" lane="8" entrytime="00:11:24.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.74" />
                    <SPLIT distance="200" swimtime="00:02:42.45" />
                    <SPLIT distance="300" swimtime="00:04:07.77" />
                    <SPLIT distance="400" swimtime="00:05:33.03" />
                    <SPLIT distance="500" swimtime="00:06:58.98" />
                    <SPLIT distance="600" swimtime="00:08:25.21" />
                    <SPLIT distance="700" swimtime="00:09:50.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Isabel Santos" birthdate="2005-12-20" gender="F" nation="BRA" license="391141" swrid="5600191" athleteid="2026" externalid="391141">
              <RESULTS>
                <RESULT eventid="1076" points="265" swimtime="00:02:55.57" resultid="2027" heatid="2250" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="165" swimtime="00:01:40.97" resultid="2028" heatid="2341" lane="3" />
                <RESULT eventid="1140" points="299" swimtime="00:01:17.31" resultid="2029" heatid="2298" lane="4" entrytime="00:01:17.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcus" lastname="Vinicius De Almeida" birthdate="2009-06-16" gender="M" nation="BRA" license="348099" swrid="5600272" athleteid="1976" externalid="348099">
              <RESULTS>
                <RESULT eventid="1196" points="443" reactiontime="+72" swimtime="00:02:26.78" resultid="1977" heatid="2338" lane="3" entrytime="00:02:30.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="444" swimtime="00:02:44.48" resultid="1978" heatid="2324" lane="1" entrytime="00:02:45.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="483" swimtime="00:00:59.69" resultid="1979" heatid="2311" lane="6" entrytime="00:01:02.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Marcos Pinto" birthdate="2006-01-26" gender="M" nation="BRA" license="391143" swrid="5600209" athleteid="2030" externalid="391143">
              <RESULTS>
                <RESULT eventid="1132" points="209" swimtime="00:01:35.80" resultid="2031" heatid="2290" lane="7" />
                <RESULT eventid="1084" points="277" swimtime="00:02:36.29" resultid="2032" heatid="2262" lane="1" entrytime="00:02:50.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="245" swimtime="00:12:01.69" resultid="2033" heatid="2330" lane="1" entrytime="00:13:09.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.51" />
                    <SPLIT distance="200" swimtime="00:02:52.68" />
                    <SPLIT distance="300" swimtime="00:04:24.41" />
                    <SPLIT distance="400" swimtime="00:05:55.92" />
                    <SPLIT distance="500" swimtime="00:07:27.90" />
                    <SPLIT distance="600" swimtime="00:08:59.65" />
                    <SPLIT distance="700" swimtime="00:10:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="300" swimtime="00:01:09.95" resultid="2034" heatid="2308" lane="2" entrytime="00:01:12.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Geovana" lastname="Dos Santos" birthdate="2011-01-20" gender="F" nation="BRA" license="367254" swrid="5602533" athleteid="1980" externalid="367254">
              <RESULTS>
                <RESULT eventid="1108" points="258" reactiontime="+70" swimtime="00:01:30.05" resultid="1981" heatid="2273" lane="3" entrytime="00:01:29.31" entrycourse="LCM" />
                <RESULT eventid="1076" points="297" swimtime="00:02:49.04" resultid="1982" heatid="2249" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="264" reactiontime="+72" swimtime="00:03:11.82" resultid="1983" heatid="2333" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="283" swimtime="00:01:18.67" resultid="1984" heatid="2298" lane="6" entrytime="00:01:20.32" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jhenyffer" lastname="Stefany Szaida" birthdate="2006-09-16" gender="F" nation="BRA" license="369326" swrid="5600264" athleteid="1988" externalid="369326">
              <RESULTS>
                <RESULT eventid="1204" points="211" swimtime="00:01:33.11" resultid="1989" heatid="2342" lane="3" entrytime="00:01:30.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Henrique Opuchkevich" birthdate="2011-02-22" gender="M" nation="BRA" license="406720" swrid="5717273" athleteid="2075" externalid="406720">
              <RESULTS>
                <RESULT eventid="1132" points="192" swimtime="00:01:38.52" resultid="2076" heatid="2288" lane="4" />
                <RESULT eventid="1116" points="169" reactiontime="+77" swimtime="00:01:33.26" resultid="2077" heatid="2277" lane="6" />
                <RESULT eventid="1084" points="230" swimtime="00:02:46.43" resultid="2078" heatid="2261" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:20.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="228" swimtime="00:01:16.67" resultid="2079" heatid="2304" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Matos Oliveira" birthdate="2007-10-26" gender="M" nation="BRA" license="391136" swrid="5600215" athleteid="2020" externalid="391136">
              <RESULTS>
                <RESULT eventid="1180" points="321" swimtime="00:10:59.82" resultid="2021" heatid="2330" lane="7" entrytime="00:11:18.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:14.13" />
                    <SPLIT distance="200" swimtime="00:02:36.83" />
                    <SPLIT distance="300" swimtime="00:04:01.15" />
                    <SPLIT distance="400" swimtime="00:05:25.18" />
                    <SPLIT distance="500" swimtime="00:06:49.95" />
                    <SPLIT distance="600" swimtime="00:08:14.47" />
                    <SPLIT distance="700" swimtime="00:09:37.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mayara" lastname="Fieber" birthdate="2008-08-20" gender="F" nation="BRA" license="391147" swrid="5600161" athleteid="2050" externalid="391147">
              <RESULTS>
                <RESULT eventid="1108" points="275" reactiontime="+68" swimtime="00:01:28.13" resultid="2051" heatid="2273" lane="6" entrytime="00:01:30.57" entrycourse="LCM" />
                <RESULT eventid="1076" points="286" swimtime="00:02:51.26" resultid="2052" heatid="2251" lane="7" entrytime="00:03:07.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="288" swimtime="00:03:06.45" resultid="2053" heatid="2333" lane="5" entrytime="00:03:25.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaylane" lastname="Marques Ferreira" birthdate="2010-03-06" gender="F" nation="BRA" license="391146" swrid="5600211" athleteid="2045" externalid="391146">
              <RESULTS>
                <RESULT eventid="1108" points="152" reactiontime="+69" swimtime="00:01:47.27" resultid="2046" heatid="2272" lane="3" entrytime="00:01:46.10" entrycourse="LCM" />
                <RESULT eventid="1076" points="189" swimtime="00:03:16.62" resultid="2047" heatid="2251" lane="8" entrytime="00:03:22.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="153" swimtime="00:01:43.61" resultid="2048" heatid="2342" lane="6" entrytime="00:01:44.70" entrycourse="LCM" />
                <RESULT eventid="1140" points="250" swimtime="00:01:22.04" resultid="2049" heatid="2298" lane="7" entrytime="00:01:28.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Madalena De Lima" birthdate="2006-05-04" gender="M" nation="BRA" license="307786" swrid="5600206" athleteid="1945" externalid="307786">
              <RESULTS>
                <RESULT eventid="1180" points="425" swimtime="00:10:01.18" resultid="1946" heatid="2330" lane="4" entrytime="00:09:57.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.95" />
                    <SPLIT distance="200" swimtime="00:02:22.61" />
                    <SPLIT distance="300" swimtime="00:03:38.29" />
                    <SPLIT distance="400" swimtime="00:04:54.78" />
                    <SPLIT distance="500" swimtime="00:06:11.24" />
                    <SPLIT distance="600" swimtime="00:07:29.06" />
                    <SPLIT distance="700" swimtime="00:08:47.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="490" swimtime="00:00:59.40" resultid="1947" heatid="2313" lane="4" entrytime="00:00:57.82" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Luiza Rimbano De Jesus" birthdate="2008-09-02" gender="F" nation="BRA" license="366819" swrid="5653297" athleteid="2061" externalid="366819">
              <RESULTS>
                <RESULT eventid="1124" points="396" swimtime="00:01:27.31" resultid="2062" heatid="2285" lane="2" entrytime="00:01:34.59" entrycourse="LCM" />
                <RESULT eventid="1076" points="463" swimtime="00:02:25.77" resultid="2063" heatid="2253" lane="4" entrytime="00:02:33.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="491" swimtime="00:01:05.51" resultid="2064" heatid="2301" lane="2" entrytime="00:01:06.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luan" lastname="Schwarzbach Paula" birthdate="2005-07-29" gender="M" nation="BRA" license="358250" swrid="5622305" athleteid="1985" externalid="358250">
              <RESULTS>
                <RESULT eventid="1132" points="367" swimtime="00:01:19.41" resultid="1986" heatid="2294" lane="1" entrytime="00:01:20.89" entrycourse="LCM" />
                <RESULT eventid="1180" points="360" swimtime="00:10:35.00" resultid="1987" heatid="2328" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.21" />
                    <SPLIT distance="200" swimtime="00:02:35.78" />
                    <SPLIT distance="300" swimtime="00:03:57.80" />
                    <SPLIT distance="400" swimtime="00:05:19.52" />
                    <SPLIT distance="500" swimtime="00:06:39.57" />
                    <SPLIT distance="600" swimtime="00:07:59.42" />
                    <SPLIT distance="700" swimtime="00:09:18.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Barros Zagonel" birthdate="2006-06-01" gender="M" nation="BRA" license="347856" swrid="5622261" athleteid="1942" externalid="347856" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1164" points="253" swimtime="00:03:18.19" resultid="1943" heatid="2322" lane="3" entrytime="00:03:23.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:31.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="385" swimtime="00:01:04.38" resultid="1944" heatid="2310" lane="4" entrytime="00:01:04.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1007" nation="BRA" region="PR" clubid="2096" swrid="93785" name="Santa Mônica Clube De Campo" shortname="Santa Mônica">
          <ATHLETES>
            <ATHLETE firstname="Joao" lastname="Guilherme Ieger" birthdate="2009-02-20" gender="M" nation="BRA" license="356888" swrid="5600180" athleteid="2132" externalid="356888">
              <RESULTS>
                <RESULT eventid="1132" points="339" swimtime="00:01:21.57" resultid="2133" heatid="2294" lane="7" entrytime="00:01:20.41" entrycourse="LCM" />
                <RESULT eventid="1084" points="397" swimtime="00:02:18.74" resultid="2134" heatid="2264" lane="1" entrytime="00:02:23.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="463" swimtime="00:01:00.53" resultid="2135" heatid="2311" lane="4" entrytime="00:01:02.44" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Novakoski" birthdate="2009-03-05" gender="F" nation="BRA" license="339136" swrid="5600225" athleteid="2123" externalid="339136">
              <RESULTS>
                <RESULT eventid="1076" points="384" swimtime="00:02:35.20" resultid="2124" heatid="2254" lane="5" entrytime="00:02:31.41" entrycourse="LCM" />
                <RESULT eventid="1172" points="367" swimtime="00:11:16.75" resultid="2125" heatid="2326" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.65" />
                    <SPLIT distance="200" swimtime="00:02:42.22" />
                    <SPLIT distance="300" swimtime="00:04:07.98" />
                    <SPLIT distance="400" swimtime="00:05:34.47" />
                    <SPLIT distance="500" swimtime="00:07:01.50" />
                    <SPLIT distance="600" swimtime="00:08:28.47" />
                    <SPLIT distance="700" swimtime="00:09:56.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucca" lastname="Maceno Araujo" birthdate="2010-09-29" gender="M" nation="BRA" license="367056" swrid="5588788" athleteid="2151" externalid="367056">
              <RESULTS>
                <RESULT eventid="1084" points="378" swimtime="00:02:21.04" resultid="2152" heatid="2263" lane="4" entrytime="00:02:24.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="361" swimtime="00:01:09.42" resultid="2153" heatid="2348" lane="1" entrytime="00:01:15.49" entrycourse="LCM" />
                <RESULT eventid="1148" points="411" swimtime="00:01:03.01" resultid="2154" heatid="2311" lane="8" entrytime="00:01:04.94" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Augusto Vaz" birthdate="2011-06-25" gender="M" nation="BRA" license="401737" swrid="5661339" athleteid="2211" externalid="401737">
              <RESULTS>
                <RESULT eventid="1084" points="229" swimtime="00:02:46.69" resultid="2212" heatid="2261" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" status="DSQ" swimtime="00:01:26.76" resultid="2213" heatid="2346" lane="6" />
                <RESULT eventid="1148" points="287" swimtime="00:01:11.01" resultid="2214" heatid="2307" lane="4" entrytime="00:01:18.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Cavassin Ieger" birthdate="2011-08-31" gender="M" nation="BRA" license="367149" swrid="5588743" athleteid="2155" externalid="367149">
              <RESULTS>
                <RESULT eventid="1132" points="219" swimtime="00:01:34.32" resultid="2156" heatid="2292" lane="2" entrytime="00:01:37.72" entrycourse="LCM" />
                <RESULT eventid="1212" points="204" swimtime="00:01:23.97" resultid="2157" heatid="2346" lane="8" />
                <RESULT eventid="1164" points="260" swimtime="00:03:16.55" resultid="2158" heatid="2322" lane="2" entrytime="00:03:30.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathalia" lastname="Lourenco Osorio" birthdate="2007-04-14" gender="F" nation="BRA" license="307465" swrid="5600203" athleteid="2100" externalid="307465">
              <RESULTS>
                <RESULT eventid="1108" points="510" reactiontime="+66" swimtime="00:01:11.71" resultid="2101" heatid="2276" lane="5" entrytime="00:01:08.78" entrycourse="LCM" />
                <RESULT eventid="1140" points="539" swimtime="00:01:03.52" resultid="2102" heatid="2302" lane="6" entrytime="00:01:01.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Celli Schneider" birthdate="2011-02-21" gender="M" nation="BRA" license="367055" swrid="5588587" athleteid="2147" externalid="367055">
              <RESULTS>
                <RESULT eventid="1116" points="331" reactiontime="+75" swimtime="00:01:14.57" resultid="2148" heatid="2280" lane="5" entrytime="00:01:16.79" entrycourse="LCM" />
                <RESULT eventid="1196" reactiontime="+75" status="DSQ" swimtime="00:02:46.39" resultid="2149" heatid="2337" lane="7" entrytime="00:02:53.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="316" swimtime="00:01:08.74" resultid="2150" heatid="2306" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Zanatta Flizikowski" birthdate="2010-01-08" gender="F" nation="BRA" license="367051" swrid="5588969" athleteid="2225" externalid="367051">
              <RESULTS>
                <RESULT eventid="1076" points="406" swimtime="00:02:32.36" resultid="2226" heatid="2255" lane="7" entrytime="00:02:24.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="276" swimtime="00:01:25.14" resultid="2227" heatid="2343" lane="8" entrytime="00:01:18.96" entrycourse="LCM" />
                <RESULT eventid="1140" points="429" swimtime="00:01:08.56" resultid="2228" heatid="2301" lane="6" entrytime="00:01:06.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietra" lastname="Vitoria Paczrowski" birthdate="2009-08-12" gender="F" nation="BRA" license="351253" swrid="5600275" athleteid="2129" externalid="351253" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1076" points="445" swimtime="00:02:27.71" resultid="2130" heatid="2255" lane="8" entrytime="00:02:28.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="434" swimtime="00:01:08.25" resultid="2131" heatid="2301" lane="7" entrytime="00:01:07.29" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otto" lastname="Hedeke" birthdate="2011-03-24" gender="M" nation="BRA" license="372643" swrid="5588738" athleteid="2188" externalid="372643">
              <RESULTS>
                <RESULT eventid="1084" points="256" swimtime="00:02:40.44" resultid="2189" heatid="2262" lane="8" entrytime="00:02:50.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1180" points="272" swimtime="00:11:37.56" resultid="2190" heatid="2329" lane="3">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.02" />
                    <SPLIT distance="200" swimtime="00:02:53.13" />
                    <SPLIT distance="300" swimtime="00:04:24.45" />
                    <SPLIT distance="400" swimtime="00:05:53.52" />
                    <SPLIT distance="500" swimtime="00:07:21.28" />
                    <SPLIT distance="600" swimtime="00:08:48.23" />
                    <SPLIT distance="700" swimtime="00:10:15.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="241" swimtime="00:01:15.29" resultid="2191" heatid="2308" lane="8" entrytime="00:01:18.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Marques Machado" birthdate="2010-02-17" gender="M" nation="BRA" license="390918" swrid="5600212" athleteid="2200" externalid="390918">
              <RESULTS>
                <RESULT eventid="1084" points="365" swimtime="00:02:22.71" resultid="2201" heatid="2263" lane="3" entrytime="00:02:27.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="260" swimtime="00:01:17.39" resultid="2202" heatid="2347" lane="6" entrytime="00:01:23.61" entrycourse="LCM" />
                <RESULT eventid="1148" points="361" swimtime="00:01:05.77" resultid="2203" heatid="2309" lane="5" entrytime="00:01:08.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Lopes Rempel" birthdate="2010-09-25" gender="M" nation="BRA" license="399739" swrid="5653294" athleteid="2207" externalid="399739">
              <RESULTS>
                <RESULT eventid="1116" points="222" reactiontime="+74" swimtime="00:01:25.14" resultid="2208" heatid="2280" lane="8" entrytime="00:01:30.57" entrycourse="LCM" />
                <RESULT eventid="1084" points="250" swimtime="00:02:41.90" resultid="2209" heatid="2261" lane="5" entrytime="00:02:57.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="250" reactiontime="+79" swimtime="00:02:57.54" resultid="2210" heatid="2336" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:25.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Marques" birthdate="2007-06-29" gender="M" nation="BRA" license="367257" swrid="5600213" athleteid="2232" externalid="367257">
              <RESULTS>
                <RESULT eventid="1084" points="318" swimtime="00:02:29.38" resultid="2233" heatid="2264" lane="3" entrytime="00:02:19.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="366" swimtime="00:01:05.46" resultid="2234" heatid="2312" lane="7" entrytime="00:01:01.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Araujo Felix" birthdate="2010-05-27" gender="F" nation="BRA" license="393157" swrid="5622260" athleteid="2239" externalid="393157">
              <RESULTS>
                <RESULT eventid="1108" points="244" reactiontime="+83" swimtime="00:01:31.66" resultid="2240" heatid="2272" lane="5" entrytime="00:01:43.56" entrycourse="LCM" />
                <RESULT eventid="1076" points="331" swimtime="00:02:43.06" resultid="2241" heatid="2251" lane="4" entrytime="00:02:53.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:17.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="239" reactiontime="+75" swimtime="00:03:18.20" resultid="2242" heatid="2333" lane="6" entrytime="00:03:41.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:34.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Gelenski Pelaio" birthdate="2005-10-10" gender="M" nation="BRA" license="281473" swrid="5600173" athleteid="2174" externalid="281473" level="UNIDOMBOSC">
              <RESULTS>
                <RESULT eventid="1084" points="464" swimtime="00:02:11.69" resultid="2175" heatid="2266" lane="5" entrytime="00:02:07.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="509" swimtime="00:01:01.90" resultid="2176" heatid="2350" lane="7" entrytime="00:01:00.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Pinterich Almeida" birthdate="2005-03-13" gender="M" nation="BRA" license="330749" swrid="5600235" athleteid="2136" externalid="330749">
              <RESULTS>
                <RESULT eventid="1084" points="610" swimtime="00:02:00.26" resultid="2137" heatid="2267" lane="3" entrytime="00:01:56.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="615" swimtime="00:00:55.08" resultid="2138" heatid="2315" lane="2" entrytime="00:00:53.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diego" lastname="Brasil Caropreso" birthdate="2009-10-29" gender="M" nation="BRA" license="399502" swrid="5653287" athleteid="2229" externalid="399502">
              <RESULTS>
                <RESULT eventid="1084" points="333" swimtime="00:02:27.12" resultid="2230" heatid="2262" lane="4" entrytime="00:02:33.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:09.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="366" swimtime="00:01:05.51" resultid="2231" heatid="2310" lane="3" entrytime="00:01:05.92" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="F" nation="BRA" license="344301" swrid="5569976" athleteid="2097" externalid="344301">
              <RESULTS>
                <RESULT eventid="1076" points="554" swimtime="00:02:17.39" resultid="2098" heatid="2255" lane="4" entrytime="00:02:22.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="548" swimtime="00:01:07.79" resultid="2099" heatid="2343" lane="4" entrytime="00:01:04.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Garcia Reschetti Rubbo" birthdate="2011-08-06" gender="F" nation="BRA" license="367053" swrid="5588720" athleteid="2143" externalid="367053" level="DCOMP IT">
              <RESULTS>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="2144" heatid="2285" lane="8" entrytime="00:01:38.24" entrycourse="LCM" />
                <RESULT eventid="1076" status="DNS" swimtime="00:00:00.00" resultid="2145" heatid="2252" lane="1" entrytime="00:02:52.99" entrycourse="LCM" />
                <RESULT eventid="1156" status="DNS" swimtime="00:00:00.00" resultid="2146" heatid="2318" lane="2" entrytime="00:03:31.04" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Breno" lastname="Borges Piekarzievicz" birthdate="2011-11-11" gender="M" nation="BRA" license="403144" swrid="5676295" athleteid="2218" externalid="403144">
              <RESULTS>
                <RESULT eventid="1132" points="118" swimtime="00:01:55.85" resultid="2219" heatid="2289" lane="7" />
                <RESULT eventid="1084" points="141" swimtime="00:03:15.96" resultid="2220" heatid="2259" lane="1">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="141" swimtime="00:04:00.93" resultid="2221" heatid="2321" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:57.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cardim Martins" birthdate="2010-09-01" gender="F" nation="BRA" license="390920" swrid="5600130" athleteid="2235" externalid="390920">
              <RESULTS>
                <RESULT eventid="1108" points="270" reactiontime="+84" swimtime="00:01:28.63" resultid="2236" heatid="2273" lane="2" entrytime="00:01:33.83" entrycourse="LCM" />
                <RESULT eventid="1076" points="278" swimtime="00:02:52.73" resultid="2237" heatid="2251" lane="2" entrytime="00:03:04.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:22.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1188" points="269" reactiontime="+80" swimtime="00:03:10.68" resultid="2238" heatid="2332" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kethelyn" lastname="Ribeiro Rodrigues" birthdate="2009-04-24" gender="F" nation="BRA" license="367052" swrid="5600244" athleteid="2139" externalid="367052">
              <RESULTS>
                <RESULT eventid="1108" points="293" swimtime="00:01:26.29" resultid="2140" heatid="2274" lane="1" entrytime="00:01:26.55" entrycourse="LCM" />
                <RESULT eventid="1076" points="409" swimtime="00:02:31.99" resultid="2141" heatid="2254" lane="7" entrytime="00:02:32.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:12.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="415" swimtime="00:01:09.30" resultid="2142" heatid="2299" lane="3" entrytime="00:01:11.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emily" lastname="Sayuri Tangueria De Lima" birthdate="2010-06-11" gender="F" nation="BRA" license="367215" swrid="5588901" athleteid="2167" externalid="367215">
              <RESULTS>
                <RESULT eventid="1092" points="318" swimtime="00:02:58.43" resultid="2168" heatid="2268" lane="6" entrytime="00:03:07.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="346" swimtime="00:01:19.02" resultid="2169" heatid="2343" lane="1" entrytime="00:01:16.95" entrycourse="LCM" />
                <RESULT eventid="1172" points="405" swimtime="00:10:54.91" resultid="2170" heatid="2327" lane="1" entrytime="00:11:12.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:15.49" />
                    <SPLIT distance="200" swimtime="00:02:38.49" />
                    <SPLIT distance="300" swimtime="00:04:01.16" />
                    <SPLIT distance="400" swimtime="00:05:24.12" />
                    <SPLIT distance="500" swimtime="00:06:49.19" />
                    <SPLIT distance="600" swimtime="00:08:14.07" />
                    <SPLIT distance="700" swimtime="00:09:35.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Vianna" birthdate="2011-01-31" gender="M" nation="BRA" license="371380" swrid="5588947" athleteid="2177" externalid="371380">
              <RESULTS>
                <RESULT eventid="1084" points="313" swimtime="00:02:30.12" resultid="2178" heatid="2259" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="278" swimtime="00:01:15.68" resultid="2179" heatid="2347" lane="7" entrytime="00:01:25.27" entrycourse="LCM" />
                <RESULT eventid="1148" points="349" swimtime="00:01:06.52" resultid="2180" heatid="2309" lane="7" entrytime="00:01:10.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="De Castro Paiva Maciel" birthdate="2008-04-10" gender="M" nation="BRA" license="378333" swrid="5622275" athleteid="2111" externalid="378333">
              <RESULTS>
                <RESULT eventid="1084" points="386" swimtime="00:02:20.03" resultid="2112" heatid="2263" lane="6" entrytime="00:02:27.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="453" swimtime="00:01:01.00" resultid="2113" heatid="2311" lane="7" entrytime="00:01:03.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wilson" lastname="Candido Souza" birthdate="2005-04-06" gender="M" nation="BRA" license="256803" swrid="5600129" athleteid="2171" externalid="256803">
              <RESULTS>
                <RESULT eventid="1132" status="DSQ" swimtime="00:01:16.50" resultid="2172" heatid="2295" lane="8" entrytime="00:01:15.05" entrycourse="LCM" />
                <RESULT eventid="1164" points="363" swimtime="00:02:55.80" resultid="2173" heatid="2323" lane="5" entrytime="00:02:52.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carol" lastname="Nalle Bejes" birthdate="2010-04-20" gender="F" nation="BRA" license="377315" swrid="5588824" athleteid="2192" externalid="377315">
              <RESULTS>
                <RESULT eventid="1124" points="389" swimtime="00:01:27.83" resultid="2193" heatid="2286" lane="3" entrytime="00:01:26.38" entrycourse="LCM" />
                <RESULT eventid="1076" points="414" swimtime="00:02:31.35" resultid="2194" heatid="2250" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:11.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="446" swimtime="00:02:59.98" resultid="2195" heatid="2319" lane="3" entrytime="00:03:07.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:27.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Leticia Durat" birthdate="2008-02-09" gender="F" nation="BRA" license="331636" swrid="5600200" athleteid="2114" externalid="331636">
              <RESULTS>
                <RESULT eventid="1124" points="346" swimtime="00:01:31.32" resultid="2115" heatid="2286" lane="2" entrytime="00:01:27.33" entrycourse="LCM" />
                <RESULT eventid="1156" points="298" swimtime="00:03:25.79" resultid="2116" heatid="2319" lane="7" entrytime="00:03:10.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:38.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Giuseppe Bulla Lanaro" birthdate="2007-05-22" gender="M" nation="BRA" license="331630" swrid="5600174" athleteid="2103" externalid="331630">
              <RESULTS>
                <RESULT eventid="1084" points="604" swimtime="00:02:00.62" resultid="2104" heatid="2267" lane="6" entrytime="00:01:57.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:00:58.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="461" swimtime="00:01:04.01" resultid="2105" heatid="2349" lane="7" entrytime="00:01:03.69" entrycourse="LCM" />
                <RESULT eventid="1148" points="626" swimtime="00:00:54.75" resultid="2106" heatid="2315" lane="1" entrytime="00:00:54.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Bello Costa Lange" birthdate="2010-09-13" gender="M" nation="BRA" license="367152" swrid="5588547" athleteid="2163" externalid="367152">
              <RESULTS>
                <RESULT eventid="1084" points="348" swimtime="00:02:24.96" resultid="2164" heatid="2263" lane="7" entrytime="00:02:29.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" status="DSQ" swimtime="00:01:11.70" resultid="2165" heatid="2348" lane="7" entrytime="00:01:14.27" entrycourse="LCM" />
                <RESULT eventid="1164" points="259" swimtime="00:03:16.68" resultid="2166" heatid="2321" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:35.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="Moreira Furtado" birthdate="2011-01-27" gender="F" nation="BRA" license="403783" swrid="5684587" athleteid="2222" externalid="403783">
              <RESULTS>
                <RESULT eventid="1108" points="107" swimtime="00:02:00.54" resultid="2223" heatid="2272" lane="1" />
                <RESULT eventid="1140" points="206" swimtime="00:01:27.48" resultid="2224" heatid="2297" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Helena Vieira Jussen" birthdate="2011-12-29" gender="F" nation="BRA" license="372282" swrid="5588740" athleteid="2184" externalid="372282">
              <RESULTS>
                <RESULT eventid="1124" points="317" swimtime="00:01:33.96" resultid="2185" heatid="2285" lane="1" entrytime="00:01:37.98" entrycourse="LCM" />
                <RESULT eventid="1076" points="274" swimtime="00:02:53.55" resultid="2186" heatid="2251" lane="1" entrytime="00:03:07.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:24.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="294" swimtime="00:03:26.73" resultid="2187" heatid="2318" lane="7" entrytime="00:03:31.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:43.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Analyce" lastname="Nunes Porto Luz" birthdate="2006-10-29" gender="F" nation="BRA" license="369322" swrid="5600226" athleteid="2107" externalid="369322">
              <RESULTS>
                <RESULT eventid="1076" points="506" swimtime="00:02:21.59" resultid="2108" heatid="2256" lane="6" entrytime="00:02:16.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1204" points="413" swimtime="00:01:14.44" resultid="2109" heatid="2343" lane="6" entrytime="00:01:11.70" entrycourse="LCM" />
                <RESULT eventid="1140" points="507" swimtime="00:01:04.81" resultid="2110" heatid="2302" lane="7" entrytime="00:01:03.42" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabio" lastname="C Burak" birthdate="2009-08-29" gender="M" nation="BRA" license="343297" swrid="5600126" athleteid="2204" externalid="343297">
              <RESULTS>
                <RESULT eventid="1084" points="419" swimtime="00:02:16.22" resultid="2205" heatid="2260" lane="2">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1196" points="409" reactiontime="+79" swimtime="00:02:30.66" resultid="2206" heatid="2336" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Blansky Hagebock" birthdate="2008-08-15" gender="M" nation="BRA" license="339123" swrid="5455418" athleteid="2126" externalid="339123">
              <RESULTS>
                <RESULT eventid="1084" points="472" swimtime="00:02:10.97" resultid="2127" heatid="2266" lane="1" entrytime="00:02:10.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:04.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1148" points="548" swimtime="00:00:57.25" resultid="2128" heatid="2314" lane="8" entrytime="00:00:57.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Ruschel" birthdate="2009-12-28" gender="F" nation="BRA" license="371384" swrid="5600251" athleteid="2181" externalid="371384">
              <RESULTS>
                <RESULT eventid="1076" points="511" swimtime="00:02:21.15" resultid="2182" heatid="2256" lane="1" entrytime="00:02:21.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:07.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1140" points="509" swimtime="00:01:04.75" resultid="2183" heatid="2302" lane="8" entrytime="00:01:04.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Inoue Kuroda" birthdate="2009-04-18" gender="M" nation="BRA" license="324700" swrid="5600190" athleteid="2120" externalid="324700">
              <RESULTS>
                <RESULT eventid="1116" points="431" reactiontime="+73" swimtime="00:01:08.28" resultid="2121" heatid="2281" lane="4" entrytime="00:01:08.75" entrycourse="LCM" />
                <RESULT eventid="1196" points="402" reactiontime="+64" swimtime="00:02:31.60" resultid="2122" heatid="2339" lane="8" entrytime="00:02:27.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Nalle Bejes" birthdate="2010-04-20" gender="F" nation="BRA" license="377323" swrid="5588826" athleteid="2196" externalid="377323">
              <RESULTS>
                <RESULT eventid="1124" points="373" swimtime="00:01:29.05" resultid="2197" heatid="2285" lane="4" entrytime="00:01:30.30" entrycourse="LCM" />
                <RESULT eventid="1188" points="280" reactiontime="+89" swimtime="00:03:08.15" resultid="2198" heatid="2333" lane="4" entrytime="00:03:14.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1156" points="381" swimtime="00:03:09.63" resultid="2199" heatid="2319" lane="8" entrytime="00:03:12.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wagner" lastname="Junior Cabral Gama" birthdate="2007-07-22" gender="M" nation="BRA" license="345334" athleteid="2243" externalid="345334">
              <RESULTS>
                <RESULT eventid="1116" points="393" reactiontime="+60" swimtime="00:01:10.44" resultid="2244" heatid="2279" lane="5" />
                <RESULT eventid="1148" points="433" swimtime="00:01:01.90" resultid="2245" heatid="2306" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabrizio" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="M" nation="BRA" license="344303" swrid="5559846" athleteid="2117" externalid="344303">
              <RESULTS>
                <RESULT eventid="1084" points="426" swimtime="00:02:15.51" resultid="2118" heatid="2264" lane="4" entrytime="00:02:18.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:06.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1212" points="447" swimtime="00:01:04.64" resultid="2119" heatid="2349" lane="8" entrytime="00:01:04.40" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Fontoura Barros" birthdate="2011-08-04" gender="F" nation="BRA" license="403143" swrid="5676298" athleteid="2215" externalid="403143">
              <RESULTS>
                <RESULT eventid="1124" points="157" swimtime="00:01:58.84" resultid="2216" heatid="2284" lane="8" />
                <RESULT eventid="1156" points="168" swimtime="00:04:09.21" resultid="2217" heatid="2317" lane="6">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:02.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Nogueira Silva" birthdate="2011-08-13" gender="M" nation="BRA" license="367150" swrid="5588832" athleteid="2159" externalid="367150">
              <RESULTS>
                <RESULT eventid="1132" points="237" swimtime="00:01:31.86" resultid="2160" heatid="2289" lane="6" />
                <RESULT eventid="1084" points="329" swimtime="00:02:27.74" resultid="2161" heatid="2262" lane="6" entrytime="00:02:37.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:10.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1164" points="258" swimtime="00:03:17.05" resultid="2162" heatid="2322" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:36.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
