<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.79911">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Campo Mourão" name="70º Jogos Escolares do Paraná (12/14 Anos) 2024" course="SCM" deadline="1969-12-31" hostclub="Secretaria do Esporte, Governo do Estado do Paraná" hostclub.url="https://www.esporte.pr.gov.br/" number="38311" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/newInterface/eventos/38311" startmethod="1" timing="AUTOMATIC" touchpad="ONESIDE" masters="F" state="PR" nation="BRA">
      <AGEDATE value="2024-01-01" type="YEAR" />
      <POOL name="Complexo Esportivo Roberto Brzezinski" lanemin="1" lanemax="8" />
      <FACILITY city="Campo Mourão" name="Complexo Esportivo Roberto Brzezinski" nation="BRA" state="PR" street="Rua Miguel Luís Pereira" street2="Bela Vista" zip="87302-140" />
      <POINTTABLE pointtableid="3016" name="FINA Point Scoring" version="2023" />
      <QUALIFY from="2023-01-01" until="2024-07-12" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-07-13" daytime="09:10" endtime="11:43" number="1" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1061" daytime="09:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1062" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1449" />
                    <RANKING order="2" place="2" resultid="1621" />
                    <RANKING order="3" place="3" resultid="1667" />
                    <RANKING order="4" place="4" resultid="1625" />
                    <RANKING order="5" place="5" resultid="1180" />
                    <RANKING order="6" place="6" resultid="2012" />
                    <RANKING order="7" place="7" resultid="1677" />
                    <RANKING order="8" place="8" resultid="1441" />
                    <RANKING order="9" place="9" resultid="1990" />
                    <RANKING order="10" place="10" resultid="1639" />
                    <RANKING order="11" place="11" resultid="1175" />
                    <RANKING order="12" place="-1" resultid="1211" />
                    <RANKING order="13" place="-1" resultid="1252" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2067" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2068" daytime="09:18" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1063" daytime="09:26" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1064" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1682" />
                    <RANKING order="2" place="2" resultid="1826" />
                    <RANKING order="3" place="3" resultid="1372" />
                    <RANKING order="4" place="4" resultid="1428" />
                    <RANKING order="5" place="5" resultid="1398" />
                    <RANKING order="6" place="6" resultid="1502" />
                    <RANKING order="7" place="7" resultid="1879" />
                    <RANKING order="8" place="8" resultid="1960" />
                    <RANKING order="9" place="9" resultid="1838" />
                    <RANKING order="10" place="10" resultid="1507" />
                    <RANKING order="11" place="11" resultid="1783" />
                    <RANKING order="12" place="12" resultid="1347" />
                    <RANKING order="13" place="13" resultid="1754" />
                    <RANKING order="14" place="14" resultid="1698" />
                    <RANKING order="15" place="15" resultid="1436" />
                    <RANKING order="16" place="16" resultid="1204" />
                    <RANKING order="17" place="17" resultid="1797" />
                    <RANKING order="18" place="18" resultid="1476" />
                    <RANKING order="19" place="19" resultid="1921" />
                    <RANKING order="20" place="20" resultid="1467" />
                    <RANKING order="21" place="21" resultid="1353" />
                    <RANKING order="22" place="22" resultid="1842" />
                    <RANKING order="23" place="23" resultid="1511" />
                    <RANKING order="24" place="24" resultid="2017" />
                    <RANKING order="25" place="25" resultid="1433" />
                    <RANKING order="26" place="25" resultid="1834" />
                    <RANKING order="27" place="27" resultid="1401" />
                    <RANKING order="28" place="28" resultid="1809" />
                    <RANKING order="29" place="29" resultid="1386" />
                    <RANKING order="30" place="30" resultid="1268" />
                    <RANKING order="31" place="31" resultid="1139" />
                    <RANKING order="32" place="31" resultid="1942" />
                    <RANKING order="33" place="33" resultid="1945" />
                    <RANKING order="34" place="34" resultid="1322" />
                    <RANKING order="35" place="35" resultid="1118" />
                    <RANKING order="36" place="36" resultid="1157" />
                    <RANKING order="37" place="37" resultid="1310" />
                    <RANKING order="38" place="38" resultid="1526" />
                    <RANKING order="39" place="39" resultid="1975" />
                    <RANKING order="40" place="40" resultid="1350" />
                    <RANKING order="41" place="41" resultid="1306" />
                    <RANKING order="42" place="42" resultid="1861" />
                    <RANKING order="43" place="43" resultid="1240" />
                    <RANKING order="44" place="44" resultid="2003" />
                    <RANKING order="45" place="45" resultid="1651" />
                    <RANKING order="46" place="46" resultid="1672" />
                    <RANKING order="47" place="47" resultid="1168" />
                    <RANKING order="48" place="48" resultid="1298" />
                    <RANKING order="49" place="49" resultid="1162" />
                    <RANKING order="50" place="50" resultid="1143" />
                    <RANKING order="51" place="51" resultid="1273" />
                    <RANKING order="52" place="52" resultid="1147" />
                    <RANKING order="53" place="53" resultid="1719" />
                    <RANKING order="54" place="54" resultid="2045" />
                    <RANKING order="55" place="55" resultid="1716" />
                    <RANKING order="56" place="56" resultid="2041" />
                    <RANKING order="57" place="-1" resultid="1662" />
                    <RANKING order="58" place="-1" resultid="1114" />
                    <RANKING order="59" place="-1" resultid="1124" />
                    <RANKING order="60" place="-1" resultid="1126" />
                    <RANKING order="61" place="-1" resultid="1224" />
                    <RANKING order="62" place="-1" resultid="1419" />
                    <RANKING order="63" place="-1" resultid="1831" />
                    <RANKING order="64" place="-1" resultid="1207" />
                    <RANKING order="65" place="-1" resultid="1303" />
                    <RANKING order="66" place="-1" resultid="1925" />
                    <RANKING order="67" place="-1" resultid="1851" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2069" daytime="09:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2070" daytime="09:28" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2071" daytime="09:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2072" daytime="09:32" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2073" daytime="09:34" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2074" daytime="09:36" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2075" daytime="09:38" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="2076" daytime="09:40" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1065" daytime="09:42" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1066" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1536" />
                    <RANKING order="2" place="2" resultid="1736" />
                    <RANKING order="3" place="3" resultid="1424" />
                    <RANKING order="4" place="4" resultid="1817" />
                    <RANKING order="5" place="5" resultid="1516" />
                    <RANKING order="6" place="6" resultid="1445" />
                    <RANKING order="7" place="7" resultid="1461" />
                    <RANKING order="8" place="8" resultid="2036" />
                    <RANKING order="9" place="9" resultid="1692" />
                    <RANKING order="10" place="10" resultid="1480" />
                    <RANKING order="11" place="11" resultid="1343" />
                    <RANKING order="12" place="12" resultid="1198" />
                    <RANKING order="13" place="13" resultid="1668" />
                    <RANKING order="14" place="14" resultid="1916" />
                    <RANKING order="15" place="15" resultid="1287" />
                    <RANKING order="16" place="16" resultid="1367" />
                    <RANKING order="17" place="17" resultid="1998" />
                    <RANKING order="18" place="18" resultid="1130" />
                    <RANKING order="19" place="19" resultid="1965" />
                    <RANKING order="20" place="20" resultid="1256" />
                    <RANKING order="21" place="21" resultid="1640" />
                    <RANKING order="22" place="22" resultid="1787" />
                    <RANKING order="23" place="23" resultid="1237" />
                    <RANKING order="24" place="24" resultid="1407" />
                    <RANKING order="25" place="25" resultid="1728" />
                    <RANKING order="26" place="26" resultid="2060" />
                    <RANKING order="27" place="27" resultid="1410" />
                    <RANKING order="28" place="28" resultid="2008" />
                    <RANKING order="29" place="29" resultid="1134" />
                    <RANKING order="30" place="30" resultid="1968" />
                    <RANKING order="31" place="31" resultid="1261" />
                    <RANKING order="32" place="32" resultid="1929" />
                    <RANKING order="33" place="33" resultid="1740" />
                    <RANKING order="34" place="34" resultid="1711" />
                    <RANKING order="35" place="35" resultid="1745" />
                    <RANKING order="36" place="36" resultid="1338" />
                    <RANKING order="37" place="37" resultid="1933" />
                    <RANKING order="38" place="38" resultid="1647" />
                    <RANKING order="39" place="39" resultid="2022" />
                    <RANKING order="40" place="40" resultid="1294" />
                    <RANKING order="41" place="41" resultid="1290" />
                    <RANKING order="42" place="42" resultid="1937" />
                    <RANKING order="43" place="43" resultid="1750" />
                    <RANKING order="44" place="-1" resultid="1122" />
                    <RANKING order="45" place="-1" resultid="1212" />
                    <RANKING order="46" place="-1" resultid="1232" />
                    <RANKING order="47" place="-1" resultid="1635" />
                    <RANKING order="48" place="-1" resultid="1769" />
                    <RANKING order="49" place="-1" resultid="1778" />
                    <RANKING order="50" place="-1" resultid="2049" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2077" daytime="09:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2078" daytime="09:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2079" daytime="09:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2080" daytime="09:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2081" daytime="09:50" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2082" daytime="09:52" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2083" daytime="09:54" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1067" daytime="09:56" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1068" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1590" />
                    <RANKING order="2" place="2" resultid="1377" />
                    <RANKING order="3" place="3" resultid="1546" />
                    <RANKING order="4" place="4" resultid="1907" />
                    <RANKING order="5" place="5" resultid="1657" />
                    <RANKING order="6" place="6" resultid="1397" />
                    <RANKING order="7" place="7" resultid="1371" />
                    <RANKING order="8" place="8" resultid="1878" />
                    <RANKING order="9" place="9" resultid="1576" />
                    <RANKING order="10" place="10" resultid="1795" />
                    <RANKING order="11" place="11" resultid="1220" />
                    <RANKING order="12" place="12" resultid="1189" />
                    <RANKING order="13" place="13" resultid="1782" />
                    <RANKING order="14" place="14" resultid="1202" />
                    <RANKING order="15" place="15" resultid="1893" />
                    <RANKING order="16" place="16" resultid="1466" />
                    <RANKING order="17" place="17" resultid="1643" />
                    <RANKING order="18" place="18" resultid="1956" />
                    <RANKING order="19" place="19" resultid="1244" />
                    <RANKING order="20" place="20" resultid="1272" />
                    <RANKING order="21" place="-1" resultid="1580" />
                    <RANKING order="22" place="-1" resultid="1897" />
                    <RANKING order="23" place="-1" resultid="1902" />
                    <RANKING order="24" place="-1" resultid="1151" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2084" daytime="09:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2085" daytime="10:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2086" daytime="10:04" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1069" daytime="10:22" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1070" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1572" />
                    <RANKING order="2" place="2" resultid="1382" />
                    <RANKING order="3" place="3" resultid="1448" />
                    <RANKING order="4" place="4" resultid="2027" />
                    <RANKING order="5" place="5" resultid="1773" />
                    <RANKING order="6" place="6" resultid="1497" />
                    <RANKING order="7" place="7" resultid="1415" />
                    <RANKING order="8" place="8" resultid="1732" />
                    <RANKING order="9" place="9" resultid="1193" />
                    <RANKING order="10" place="10" resultid="1444" />
                    <RANKING order="11" place="11" resultid="1687" />
                    <RANKING order="12" place="12" resultid="1216" />
                    <RANKING order="13" place="13" resultid="1764" />
                    <RANKING order="14" place="14" resultid="1521" />
                    <RANKING order="15" place="15" resultid="1286" />
                    <RANKING order="16" place="16" resultid="1440" />
                    <RANKING order="17" place="17" resultid="1330" />
                    <RANKING order="18" place="18" resultid="1888" />
                    <RANKING order="19" place="19" resultid="1952" />
                    <RANKING order="20" place="20" resultid="1723" />
                    <RANKING order="21" place="21" resultid="1129" />
                    <RANKING order="22" place="22" resultid="1236" />
                    <RANKING order="23" place="23" resultid="1989" />
                    <RANKING order="24" place="-1" resultid="1260" />
                    <RANKING order="25" place="-1" resultid="1706" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2087" daytime="10:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2088" daytime="10:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2089" daytime="10:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2090" daytime="10:34" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1071" daytime="10:36" gender="M" number="6" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1072" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1883" />
                    <RANKING order="2" place="2" resultid="1825" />
                    <RANKING order="3" place="3" resultid="1594" />
                    <RANKING order="4" place="4" resultid="1994" />
                    <RANKING order="5" place="5" resultid="1185" />
                    <RANKING order="6" place="6" resultid="1697" />
                    <RANKING order="7" place="7" resultid="1791" />
                    <RANKING order="8" place="8" resultid="1796" />
                    <RANKING order="9" place="9" resultid="1559" />
                    <RANKING order="10" place="9" resultid="1563" />
                    <RANKING order="11" place="11" resultid="1248" />
                    <RANKING order="12" place="12" resultid="1813" />
                    <RANKING order="13" place="13" resultid="1346" />
                    <RANKING order="14" place="14" resultid="1808" />
                    <RANKING order="15" place="15" resultid="1475" />
                    <RANKING order="16" place="16" resultid="1245" />
                    <RANKING order="17" place="17" resultid="1941" />
                    <RANKING order="18" place="18" resultid="1432" />
                    <RANKING order="19" place="19" resultid="1613" />
                    <RANKING order="20" place="20" resultid="1799" />
                    <RANKING order="21" place="21" resultid="1161" />
                    <RANKING order="22" place="-1" resultid="1830" />
                    <RANKING order="23" place="-1" resultid="1206" />
                    <RANKING order="24" place="-1" resultid="1302" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2091" daytime="10:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2092" daytime="10:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2093" daytime="10:40" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1073" daytime="10:42" gender="F" number="7" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1074" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1531" />
                    <RANKING order="2" place="2" resultid="1866" />
                    <RANKING order="3" place="3" resultid="2028" />
                    <RANKING order="4" place="4" resultid="1342" />
                    <RANKING order="5" place="5" resultid="1911" />
                    <RANKING order="6" place="6" resultid="1847" />
                    <RANKING order="7" place="7" resultid="1366" />
                    <RANKING order="8" place="8" resultid="2013" />
                    <RANKING order="9" place="9" resultid="1584" />
                    <RANKING order="10" place="10" resultid="1678" />
                    <RANKING order="11" place="11" resultid="1406" />
                    <RANKING order="12" place="12" resultid="1971" />
                    <RANKING order="13" place="13" resultid="1554" />
                    <RANKING order="14" place="14" resultid="1964" />
                    <RANKING order="15" place="15" resultid="2007" />
                    <RANKING order="16" place="-1" resultid="1253" />
                    <RANKING order="17" place="-1" resultid="1456" />
                    <RANKING order="18" place="-1" resultid="1707" />
                    <RANKING order="19" place="-1" resultid="1759" />
                    <RANKING order="20" place="-1" resultid="1768" />
                    <RANKING order="21" place="-1" resultid="1777" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2094" daytime="10:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2095" daytime="10:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2096" daytime="10:48" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1075" daytime="10:50" gender="M" number="8" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1076" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1591" />
                    <RANKING order="2" place="2" resultid="1378" />
                    <RANKING order="3" place="3" resultid="1541" />
                    <RANKING order="4" place="4" resultid="1617" />
                    <RANKING order="5" place="5" resultid="1547" />
                    <RANKING order="6" place="6" resultid="1908" />
                    <RANKING order="7" place="7" resultid="1493" />
                    <RANKING order="8" place="8" resultid="1489" />
                    <RANKING order="9" place="9" resultid="1506" />
                    <RANKING order="10" place="10" resultid="1228" />
                    <RANKING order="11" place="11" resultid="1894" />
                    <RANKING order="12" place="12" resultid="1203" />
                    <RANKING order="13" place="13" resultid="1392" />
                    <RANKING order="14" place="14" resultid="1948" />
                    <RANKING order="15" place="15" resultid="1874" />
                    <RANKING order="16" place="16" resultid="1550" />
                    <RANKING order="17" place="17" resultid="1598" />
                    <RANKING order="18" place="-1" resultid="1567" />
                    <RANKING order="19" place="-1" resultid="1156" />
                    <RANKING order="20" place="-1" resultid="1898" />
                    <RANKING order="21" place="-1" resultid="1608" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2097" daytime="10:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2098" daytime="10:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2099" daytime="11:00" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1077" daytime="11:20" gender="X" number="9" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1078" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1453" />
                    <RANKING order="2" place="2" resultid="1587" />
                    <RANKING order="3" place="3" resultid="1632" />
                    <RANKING order="4" place="4" resultid="1279" />
                    <RANKING order="5" place="5" resultid="1363" />
                    <RANKING order="6" place="6" resultid="1982" />
                    <RANKING order="7" place="7" resultid="1315" />
                    <RANKING order="8" place="-1" resultid="1654" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2100" daytime="11:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-07-13" daytime="16:10" endtime="18:19" number="2" officialmeeting="15:10" teamleadermeeting="15:20" warmupfrom="15:00" warmupuntil="16:00">
          <EVENTS>
            <EVENT eventid="1079" daytime="16:10" gender="M" number="10" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1080" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1543" />
                    <RANKING order="2" place="2" resultid="1592" />
                    <RANKING order="3" place="3" resultid="1430" />
                    <RANKING order="4" place="4" resultid="1187" />
                    <RANKING order="5" place="5" resultid="1595" />
                    <RANKING order="6" place="6" resultid="1663" />
                    <RANKING order="7" place="7" resultid="1318" />
                    <RANKING order="8" place="8" resultid="1508" />
                    <RANKING order="9" place="9" resultid="1560" />
                    <RANKING order="10" place="10" resultid="1839" />
                    <RANKING order="11" place="11" resultid="1792" />
                    <RANKING order="12" place="12" resultid="1393" />
                    <RANKING order="13" place="13" resultid="1348" />
                    <RANKING order="14" place="14" resultid="1551" />
                    <RANKING order="15" place="15" resultid="1645" />
                    <RANKING order="16" place="16" resultid="1949" />
                    <RANKING order="17" place="17" resultid="1312" />
                    <RANKING order="18" place="18" resultid="1170" />
                    <RANKING order="19" place="19" resultid="1300" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2101" daytime="16:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2102" daytime="16:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2103" daytime="16:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2153" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1081" daytime="16:32" gender="F" number="11" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1082" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1282" />
                    <RANKING order="2" place="2" resultid="1848" />
                    <RANKING order="3" place="3" resultid="1327" />
                    <RANKING order="4" place="4" resultid="1194" />
                    <RANKING order="5" place="5" resultid="1485" />
                    <RANKING order="6" place="6" resultid="2037" />
                    <RANKING order="7" place="7" resultid="1774" />
                    <RANKING order="8" place="8" resultid="1416" />
                    <RANKING order="9" place="9" resultid="1604" />
                    <RANKING order="10" place="10" resultid="1918" />
                    <RANKING order="11" place="11" resultid="1630" />
                    <RANKING order="12" place="12" resultid="1200" />
                    <RANKING order="13" place="13" resultid="1821" />
                    <RANKING order="14" place="14" resultid="1972" />
                    <RANKING order="15" place="15" resultid="2032" />
                    <RANKING order="16" place="16" resultid="1966" />
                    <RANKING order="17" place="17" resultid="2056" />
                    <RANKING order="18" place="18" resultid="1265" />
                    <RANKING order="19" place="19" resultid="1472" />
                    <RANKING order="20" place="20" resultid="1934" />
                    <RANKING order="21" place="21" resultid="1339" />
                    <RANKING order="22" place="22" resultid="1649" />
                    <RANKING order="23" place="-1" resultid="2023" />
                    <RANKING order="24" place="-1" resultid="1296" />
                    <RANKING order="25" place="-1" resultid="1233" />
                    <RANKING order="26" place="-1" resultid="1262" />
                    <RANKING order="27" place="-1" resultid="1457" />
                    <RANKING order="28" place="-1" resultid="1637" />
                    <RANKING order="29" place="-1" resultid="1770" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2104" daytime="16:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2105" daytime="16:34" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2106" daytime="16:36" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2107" daytime="16:38" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1083" daytime="16:42" gender="M" number="12" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1084" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1755" />
                    <RANKING order="2" place="2" resultid="1804" />
                    <RANKING order="3" place="3" resultid="1618" />
                    <RANKING order="4" place="4" resultid="1494" />
                    <RANKING order="5" place="5" resultid="1961" />
                    <RANKING order="6" place="6" resultid="1437" />
                    <RANKING order="7" place="7" resultid="1319" />
                    <RANKING order="8" place="8" resultid="1568" />
                    <RANKING order="9" place="9" resultid="1229" />
                    <RANKING order="10" place="10" resultid="1858" />
                    <RANKING order="11" place="11" resultid="1922" />
                    <RANKING order="12" place="12" resultid="1985" />
                    <RANKING order="13" place="13" resultid="1249" />
                    <RANKING order="14" place="14" resultid="1323" />
                    <RANKING order="15" place="15" resultid="1358" />
                    <RANKING order="16" place="16" resultid="1875" />
                    <RANKING order="17" place="17" resultid="1388" />
                    <RANKING order="18" place="18" resultid="1141" />
                    <RANKING order="19" place="19" resultid="2019" />
                    <RANKING order="20" place="20" resultid="1402" />
                    <RANKING order="21" place="21" resultid="1599" />
                    <RANKING order="22" place="22" resultid="1614" />
                    <RANKING order="23" place="23" resultid="1354" />
                    <RANKING order="24" place="24" resultid="1862" />
                    <RANKING order="25" place="25" resultid="1119" />
                    <RANKING order="26" place="26" resultid="1242" />
                    <RANKING order="27" place="27" resultid="1976" />
                    <RANKING order="28" place="28" resultid="1673" />
                    <RANKING order="29" place="29" resultid="1145" />
                    <RANKING order="30" place="-1" resultid="1720" />
                    <RANKING order="31" place="-1" resultid="2046" />
                    <RANKING order="32" place="-1" resultid="1226" />
                    <RANKING order="33" place="-1" resultid="1609" />
                    <RANKING order="34" place="-1" resultid="1853" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2108" daytime="16:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2109" daytime="16:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2110" daytime="16:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2111" daytime="16:48" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1085" daytime="16:50" gender="F" number="13" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1086" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1425" />
                    <RANKING order="2" place="2" resultid="1537" />
                    <RANKING order="3" place="3" resultid="1867" />
                    <RANKING order="4" place="4" resultid="1737" />
                    <RANKING order="5" place="5" resultid="1383" />
                    <RANKING order="6" place="6" resultid="1498" />
                    <RANKING order="7" place="7" resultid="1733" />
                    <RANKING order="8" place="8" resultid="1344" />
                    <RANKING order="9" place="9" resultid="1818" />
                    <RANKING order="10" place="10" resultid="1446" />
                    <RANKING order="11" place="11" resultid="1517" />
                    <RANKING order="12" place="12" resultid="1669" />
                    <RANKING order="13" place="13" resultid="1693" />
                    <RANKING order="14" place="14" resultid="1199" />
                    <RANKING order="15" place="15" resultid="1765" />
                    <RANKING order="16" place="16" resultid="1217" />
                    <RANKING order="17" place="17" resultid="1679" />
                    <RANKING order="18" place="18" resultid="1889" />
                    <RANKING order="19" place="19" resultid="1288" />
                    <RANKING order="20" place="20" resultid="1331" />
                    <RANKING order="21" place="21" resultid="1442" />
                    <RANKING order="22" place="22" resultid="1257" />
                    <RANKING order="23" place="23" resultid="1953" />
                    <RANKING order="24" place="24" resultid="1991" />
                    <RANKING order="25" place="25" resultid="1238" />
                    <RANKING order="26" place="26" resultid="1917" />
                    <RANKING order="27" place="27" resultid="1724" />
                    <RANKING order="28" place="28" resultid="1641" />
                    <RANKING order="29" place="29" resultid="2009" />
                    <RANKING order="30" place="30" resultid="1135" />
                    <RANKING order="31" place="31" resultid="1411" />
                    <RANKING order="32" place="32" resultid="1264" />
                    <RANKING order="33" place="33" resultid="1702" />
                    <RANKING order="34" place="34" resultid="1471" />
                    <RANKING order="35" place="35" resultid="1741" />
                    <RANKING order="36" place="36" resultid="1712" />
                    <RANKING order="37" place="37" resultid="1746" />
                    <RANKING order="38" place="38" resultid="1291" />
                    <RANKING order="39" place="39" resultid="1648" />
                    <RANKING order="40" place="40" resultid="1295" />
                    <RANKING order="41" place="-1" resultid="1213" />
                    <RANKING order="42" place="-1" resultid="1636" />
                    <RANKING order="43" place="-1" resultid="1708" />
                    <RANKING order="44" place="-1" resultid="1999" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2112" daytime="16:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2113" daytime="16:54" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2114" daytime="16:56" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2115" daytime="17:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2116" daytime="17:02" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2117" daytime="17:04" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1087" daytime="17:22" gender="M" number="14" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1088" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1884" />
                    <RANKING order="2" place="2" resultid="1429" />
                    <RANKING order="3" place="2" resultid="1542" />
                    <RANKING order="4" place="4" resultid="1658" />
                    <RANKING order="5" place="5" resultid="1503" />
                    <RANKING order="6" place="6" resultid="1186" />
                    <RANKING order="7" place="7" resultid="1683" />
                    <RANKING order="8" place="8" resultid="1548" />
                    <RANKING order="9" place="9" resultid="1880" />
                    <RANKING order="10" place="10" resultid="1995" />
                    <RANKING order="11" place="11" resultid="1490" />
                    <RANKING order="12" place="12" resultid="1784" />
                    <RANKING order="13" place="13" resultid="1564" />
                    <RANKING order="14" place="14" resultid="1190" />
                    <RANKING order="15" place="15" resultid="1857" />
                    <RANKING order="16" place="16" resultid="1895" />
                    <RANKING order="17" place="17" resultid="1434" />
                    <RANKING order="18" place="18" resultid="1512" />
                    <RANKING order="19" place="19" resultid="1835" />
                    <RANKING order="20" place="20" resultid="1870" />
                    <RANKING order="21" place="21" resultid="1246" />
                    <RANKING order="22" place="22" resultid="1814" />
                    <RANKING order="23" place="23" resultid="1843" />
                    <RANKING order="24" place="24" resultid="1810" />
                    <RANKING order="25" place="25" resultid="2018" />
                    <RANKING order="26" place="26" resultid="1357" />
                    <RANKING order="27" place="27" resultid="1269" />
                    <RANKING order="28" place="28" resultid="1387" />
                    <RANKING order="29" place="29" resultid="1957" />
                    <RANKING order="30" place="30" resultid="1140" />
                    <RANKING order="31" place="31" resultid="1527" />
                    <RANKING order="32" place="32" resultid="1644" />
                    <RANKING order="33" place="33" resultid="1311" />
                    <RANKING order="34" place="34" resultid="1334" />
                    <RANKING order="35" place="35" resultid="1800" />
                    <RANKING order="36" place="36" resultid="1652" />
                    <RANKING order="37" place="37" resultid="1307" />
                    <RANKING order="38" place="38" resultid="1241" />
                    <RANKING order="39" place="39" resultid="1351" />
                    <RANKING order="40" place="40" resultid="1169" />
                    <RANKING order="41" place="41" resultid="2004" />
                    <RANKING order="42" place="42" resultid="1299" />
                    <RANKING order="43" place="43" resultid="1163" />
                    <RANKING order="44" place="44" resultid="1144" />
                    <RANKING order="45" place="45" resultid="1148" />
                    <RANKING order="46" place="-1" resultid="1477" />
                    <RANKING order="47" place="-1" resultid="1581" />
                    <RANKING order="48" place="-1" resultid="1225" />
                    <RANKING order="49" place="-1" resultid="1420" />
                    <RANKING order="50" place="-1" resultid="1903" />
                    <RANKING order="51" place="-1" resultid="1208" />
                    <RANKING order="52" place="-1" resultid="1304" />
                    <RANKING order="53" place="-1" resultid="1152" />
                    <RANKING order="54" place="-1" resultid="1852" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2118" daytime="17:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2119" daytime="17:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2120" daytime="17:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2121" daytime="17:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2122" daytime="17:34" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2123" daytime="17:36" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="2124" daytime="17:38" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1089" daytime="17:42" gender="F" number="15" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1090" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1532" />
                    <RANKING order="2" place="2" resultid="1573" />
                    <RANKING order="3" place="3" resultid="1481" />
                    <RANKING order="4" place="4" resultid="1622" />
                    <RANKING order="5" place="5" resultid="1603" />
                    <RANKING order="6" place="6" resultid="1626" />
                    <RANKING order="7" place="7" resultid="1462" />
                    <RANKING order="8" place="8" resultid="1326" />
                    <RANKING order="9" place="9" resultid="1181" />
                    <RANKING order="10" place="10" resultid="1585" />
                    <RANKING order="11" place="11" resultid="1629" />
                    <RANKING order="12" place="12" resultid="1688" />
                    <RANKING order="13" place="13" resultid="1912" />
                    <RANKING order="14" place="14" resultid="1555" />
                    <RANKING order="15" place="15" resultid="1788" />
                    <RANKING order="16" place="16" resultid="1703" />
                    <RANKING order="17" place="-1" resultid="2031" />
                    <RANKING order="18" place="-1" resultid="1176" />
                    <RANKING order="19" place="-1" resultid="1760" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2125" daytime="17:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2126" daytime="17:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2127" daytime="17:52" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1091" daytime="18:12" gender="M" number="16" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1092" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1277" />
                    <RANKING order="2" place="2" resultid="1361" />
                    <RANKING order="3" place="3" resultid="1980" />
                    <RANKING order="4" place="-1" resultid="1313" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2128" daytime="18:12" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1093" daytime="18:16" gender="F" number="17" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1094" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1359" />
                    <RANKING order="2" place="2" resultid="1275" />
                    <RANKING order="3" place="3" resultid="1978" />
                    <RANKING order="4" place="-1" resultid="1451" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2129" daytime="18:16" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-07-14" daytime="09:10" endtime="10:42" number="3" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1095" daytime="09:10" gender="F" number="18" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1096" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1533" />
                    <RANKING order="2" place="2" resultid="1450" />
                    <RANKING order="3" place="3" resultid="1868" />
                    <RANKING order="4" place="4" resultid="1623" />
                    <RANKING order="5" place="5" resultid="1586" />
                    <RANKING order="6" place="6" resultid="1463" />
                    <RANKING order="7" place="7" resultid="1913" />
                    <RANKING order="8" place="8" resultid="1689" />
                    <RANKING order="9" place="9" resultid="2014" />
                    <RANKING order="10" place="10" resultid="1766" />
                    <RANKING order="11" place="11" resultid="1368" />
                    <RANKING order="12" place="12" resultid="1408" />
                    <RANKING order="13" place="13" resultid="1177" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2130" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2131" daytime="09:14" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1097" daytime="09:16" gender="M" number="19" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1098" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1885" />
                    <RANKING order="2" place="2" resultid="1379" />
                    <RANKING order="3" place="3" resultid="1596" />
                    <RANKING order="4" place="4" resultid="1996" />
                    <RANKING order="5" place="5" resultid="1699" />
                    <RANKING order="6" place="6" resultid="1561" />
                    <RANKING order="7" place="7" resultid="1565" />
                    <RANKING order="8" place="8" resultid="1491" />
                    <RANKING order="9" place="9" resultid="1221" />
                    <RANKING order="10" place="10" resultid="1871" />
                    <RANKING order="11" place="11" resultid="1664" />
                    <RANKING order="12" place="12" resultid="1513" />
                    <RANKING order="13" place="13" resultid="1250" />
                    <RANKING order="14" place="14" resultid="1552" />
                    <RANKING order="15" place="15" resultid="1950" />
                    <RANKING order="16" place="16" resultid="1600" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2132" daytime="09:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2133" daytime="09:20" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1099" daytime="09:22" gender="F" number="20" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1100" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1574" />
                    <RANKING order="2" place="2" resultid="2029" />
                    <RANKING order="3" place="3" resultid="1775" />
                    <RANKING order="4" place="4" resultid="1384" />
                    <RANKING order="5" place="4" resultid="1538" />
                    <RANKING order="6" place="6" resultid="1426" />
                    <RANKING order="7" place="7" resultid="1734" />
                    <RANKING order="8" place="8" resultid="1523" />
                    <RANKING order="9" place="9" resultid="1417" />
                    <RANKING order="10" place="10" resultid="1195" />
                    <RANKING order="11" place="11" resultid="1819" />
                    <RANKING order="12" place="12" resultid="1218" />
                    <RANKING order="13" place="13" resultid="1789" />
                    <RANKING order="14" place="14" resultid="1890" />
                    <RANKING order="15" place="15" resultid="1729" />
                    <RANKING order="16" place="16" resultid="1332" />
                    <RANKING order="17" place="17" resultid="1258" />
                    <RANKING order="18" place="18" resultid="1973" />
                    <RANKING order="19" place="19" resultid="2000" />
                    <RANKING order="20" place="20" resultid="1725" />
                    <RANKING order="21" place="21" resultid="1136" />
                    <RANKING order="22" place="22" resultid="1131" />
                    <RANKING order="23" place="23" resultid="2024" />
                    <RANKING order="24" place="24" resultid="1412" />
                    <RANKING order="25" place="25" resultid="1473" />
                    <RANKING order="26" place="26" resultid="1969" />
                    <RANKING order="27" place="27" resultid="1930" />
                    <RANKING order="28" place="28" resultid="1935" />
                    <RANKING order="29" place="29" resultid="1292" />
                    <RANKING order="30" place="30" resultid="1713" />
                    <RANKING order="31" place="31" resultid="1751" />
                    <RANKING order="32" place="-1" resultid="1747" />
                    <RANKING order="33" place="-1" resultid="1938" />
                    <RANKING order="34" place="-1" resultid="1254" />
                    <RANKING order="35" place="-1" resultid="1742" />
                    <RANKING order="36" place="-1" resultid="1761" />
                    <RANKING order="37" place="-1" resultid="2050" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2134" daytime="09:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2135" daytime="09:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2136" daytime="09:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2137" daytime="09:32" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2138" daytime="09:36" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1101" daytime="09:38" gender="M" number="21" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1102" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1374" />
                    <RANKING order="2" place="2" resultid="1684" />
                    <RANKING order="3" place="3" resultid="1827" />
                    <RANKING order="4" place="4" resultid="1659" />
                    <RANKING order="5" place="5" resultid="1399" />
                    <RANKING order="6" place="6" resultid="1909" />
                    <RANKING order="7" place="7" resultid="1578" />
                    <RANKING order="8" place="8" resultid="1222" />
                    <RANKING order="9" place="9" resultid="1840" />
                    <RANKING order="10" place="10" resultid="1899" />
                    <RANKING order="11" place="11" resultid="1962" />
                    <RANKING order="12" place="12" resultid="1793" />
                    <RANKING order="13" place="13" resultid="1582" />
                    <RANKING order="14" place="14" resultid="1468" />
                    <RANKING order="15" place="15" resultid="1923" />
                    <RANKING order="16" place="16" resultid="1191" />
                    <RANKING order="17" place="17" resultid="1987" />
                    <RANKING order="18" place="18" resultid="1403" />
                    <RANKING order="19" place="19" resultid="1844" />
                    <RANKING order="20" place="20" resultid="1832" />
                    <RANKING order="21" place="21" resultid="1815" />
                    <RANKING order="22" place="22" resultid="1270" />
                    <RANKING order="23" place="23" resultid="1158" />
                    <RANKING order="24" place="24" resultid="1528" />
                    <RANKING order="25" place="25" resultid="1336" />
                    <RANKING order="26" place="26" resultid="1977" />
                    <RANKING order="27" place="27" resultid="1801" />
                    <RANKING order="28" place="28" resultid="1653" />
                    <RANKING order="29" place="29" resultid="1274" />
                    <RANKING order="30" place="-1" resultid="1717" />
                    <RANKING order="31" place="-1" resultid="2042" />
                    <RANKING order="32" place="-1" resultid="1115" />
                    <RANKING order="33" place="-1" resultid="1308" />
                    <RANKING order="34" place="-1" resultid="1421" />
                    <RANKING order="35" place="-1" resultid="1904" />
                    <RANKING order="36" place="-1" resultid="1926" />
                    <RANKING order="37" place="-1" resultid="1153" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2139" daytime="09:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2140" daytime="09:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2141" daytime="09:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2142" daytime="09:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2143" daytime="09:50" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1103" daytime="09:52" gender="F" number="22" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1104" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1283" />
                    <RANKING order="2" place="2" resultid="1328" />
                    <RANKING order="3" place="3" resultid="2066" />
                    <RANKING order="4" place="4" resultid="1486" />
                    <RANKING order="5" place="5" resultid="1849" />
                    <RANKING order="6" place="6" resultid="1605" />
                    <RANKING order="7" place="7" resultid="2038" />
                    <RANKING order="8" place="8" resultid="1631" />
                    <RANKING order="9" place="9" resultid="1499" />
                    <RANKING order="10" place="10" resultid="1627" />
                    <RANKING order="11" place="11" resultid="1738" />
                    <RANKING order="12" place="12" resultid="1694" />
                    <RANKING order="13" place="13" resultid="1822" />
                    <RANKING order="14" place="14" resultid="1182" />
                    <RANKING order="15" place="15" resultid="1522" />
                    <RANKING order="16" place="16" resultid="1518" />
                    <RANKING order="17" place="17" resultid="1779" />
                    <RANKING order="18" place="18" resultid="2033" />
                    <RANKING order="19" place="19" resultid="1556" />
                    <RANKING order="20" place="20" resultid="1954" />
                    <RANKING order="21" place="21" resultid="2059" />
                    <RANKING order="22" place="22" resultid="1266" />
                    <RANKING order="23" place="23" resultid="1704" />
                    <RANKING order="24" place="-1" resultid="1340" />
                    <RANKING order="25" place="-1" resultid="1234" />
                    <RANKING order="26" place="-1" resultid="1458" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2144" daytime="09:52" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2145" daytime="09:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2146" daytime="10:00" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2147" daytime="10:02" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1105" daytime="10:06" gender="M" number="23" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1106" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1756" />
                    <RANKING order="2" place="2" resultid="1619" />
                    <RANKING order="3" place="3" resultid="1805" />
                    <RANKING order="4" place="4" resultid="1495" />
                    <RANKING order="5" place="5" resultid="1569" />
                    <RANKING order="6" place="6" resultid="1504" />
                    <RANKING order="7" place="7" resultid="1320" />
                    <RANKING order="8" place="8" resultid="1230" />
                    <RANKING order="9" place="9" resultid="1577" />
                    <RANKING order="10" place="10" resultid="1438" />
                    <RANKING order="11" place="11" resultid="1859" />
                    <RANKING order="12" place="12" resultid="1872" />
                    <RANKING order="13" place="13" resultid="1324" />
                    <RANKING order="14" place="14" resultid="1394" />
                    <RANKING order="15" place="15" resultid="1355" />
                    <RANKING order="16" place="16" resultid="1615" />
                    <RANKING order="17" place="17" resultid="1958" />
                    <RANKING order="18" place="18" resultid="1863" />
                    <RANKING order="19" place="19" resultid="1335" />
                    <RANKING order="20" place="20" resultid="1674" />
                    <RANKING order="21" place="-1" resultid="1986" />
                    <RANKING order="22" place="-1" resultid="1876" />
                    <RANKING order="23" place="-1" resultid="1610" />
                    <RANKING order="24" place="-1" resultid="1854" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2148" daytime="10:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2149" daytime="10:08" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2150" daytime="10:12" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1107" daytime="10:28" gender="F" number="24" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1108" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1360" />
                    <RANKING order="2" place="2" resultid="1276" />
                    <RANKING order="3" place="3" resultid="1979" />
                    <RANKING order="4" place="-1" resultid="2154" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2151" daytime="10:28" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1109" daytime="10:34" gender="M" number="25" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="4" stroke="MEDLEY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1110" agemax="-1" agemin="-1">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1278" />
                    <RANKING order="2" place="2" resultid="1362" />
                    <RANKING order="3" place="3" resultid="1981" />
                    <RANKING order="4" place="-1" resultid="1314" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2152" daytime="10:34" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="17693" nation="BRA" region="PR" clubid="2043" name="7º Colégio Da Polícia Militar, União Da Vitória" shortname="Unvt-7ºcpm,C">
          <ATHLETES>
            <ATHLETE firstname="Joao" lastname="Pedro Da Silva Souza" birthdate="2010-11-10" gender="M" nation="BRA" license="V413932" athleteid="2044" externalid="V413932">
              <RESULTS>
                <RESULT eventid="1063" points="46" swimtime="00:00:56.19" resultid="2045" heatid="2075" lane="7" />
                <RESULT eventid="1083" status="DSQ" swimtime="00:01:31.06" resultid="2046" heatid="2108" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15595" nation="BRA" region="PR" clubid="1762" name="Colégio Adventista De Maringá" shortname="Mrga-Adventista,C">
          <ATHLETES>
            <ATHLETE firstname="Yasmin" lastname="Ghelere" birthdate="2011-04-03" gender="F" nation="BRA" license="368146" swrid="5603843" athleteid="1763" externalid="368146">
              <RESULTS>
                <RESULT eventid="1069" points="303" swimtime="00:01:21.65" resultid="1764" heatid="2089" lane="2" entrytime="00:01:23.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="355" swimtime="00:01:10.95" resultid="1765" heatid="2115" lane="3" entrytime="00:01:12.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="228" swimtime="00:01:28.37" resultid="1766" heatid="2130" lane="5" entrytime="00:01:36.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Sales" birthdate="2011-02-28" gender="F" nation="BRA" license="374103" swrid="5616410" athleteid="1767" externalid="374103">
              <RESULTS>
                <RESULT eventid="1073" status="DNS" swimtime="00:00:00.00" resultid="1768" heatid="2096" lane="5" entrytime="00:00:32.99" entrycourse="SCM" />
                <RESULT eventid="1065" status="DNS" swimtime="00:00:00.00" resultid="1769" heatid="2083" lane="2" entrytime="00:00:30.42" entrycourse="SCM" />
                <RESULT eventid="1081" status="DNS" swimtime="00:00:00.00" resultid="1770" heatid="2107" lane="1" entrytime="00:00:40.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="9735" nation="BRA" region="PR" clubid="1823" name="Colégio São Francisco Xavier, Maringá" shortname="Mrga-Franci.Xavier,C">
          <ATHLETES>
            <ATHLETE firstname="Pedro" lastname="Henrique Campelo" birthdate="2011-09-12" gender="M" nation="BRA" license="366963" swrid="5588742" athleteid="1824" externalid="366963">
              <RESULTS>
                <RESULT eventid="1071" points="365" swimtime="00:00:30.43" resultid="1825" heatid="2093" lane="5" entrytime="00:00:31.79" entrycourse="SCM" />
                <RESULT eventid="1063" points="432" swimtime="00:00:26.65" resultid="1826" heatid="2076" lane="7" entrytime="00:00:28.67" entrycourse="SCM" />
                <RESULT eventid="1101" points="358" swimtime="00:00:31.13" resultid="1827" heatid="2143" lane="2" entrytime="00:00:34.05" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6525" nation="BRA" region="PR" clubid="1611" name="Colégio Santa Maria, Cascavel" shortname="Cvel-Santa Maria, C">
          <ATHLETES>
            <ATHLETE firstname="Breno" lastname="Zanella Janke" birthdate="2011-04-26" gender="M" nation="BRA" license="365697" swrid="5588970" athleteid="1616" externalid="365697">
              <RESULTS>
                <RESULT eventid="1075" points="405" swimtime="00:02:28.15" resultid="1617" heatid="2099" lane="2" entrytime="00:02:32.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:12.01" />
                    <SPLIT distance="150" swimtime="00:01:54.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="343" swimtime="00:00:35.63" resultid="1618" heatid="2111" lane="3" entrytime="00:00:37.79" entrycourse="SCM" />
                <RESULT eventid="1105" points="348" swimtime="00:01:18.52" resultid="1619" heatid="2150" lane="6" entrytime="00:01:22.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Bertelli Weirich" birthdate="2011-03-18" gender="F" nation="BRA" license="369534" swrid="5588552" athleteid="1620" externalid="369534">
              <RESULTS>
                <RESULT eventid="1061" points="452" swimtime="00:05:01.24" resultid="1621" heatid="2068" lane="5" entrytime="00:05:03.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:10.74" />
                    <SPLIT distance="150" swimtime="00:01:48.68" />
                    <SPLIT distance="200" swimtime="00:02:27.51" />
                    <SPLIT distance="250" swimtime="00:03:06.36" />
                    <SPLIT distance="300" swimtime="00:03:45.37" />
                    <SPLIT distance="350" swimtime="00:04:24.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1089" points="408" swimtime="00:02:44.30" resultid="1622" heatid="2127" lane="7" entrytime="00:02:50.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                    <SPLIT distance="100" swimtime="00:01:19.69" />
                    <SPLIT distance="150" swimtime="00:02:07.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="328" swimtime="00:01:18.32" resultid="1623" heatid="2131" lane="6" entrytime="00:01:19.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Colaco Da Conceicao" birthdate="2011-05-25" gender="F" nation="BRA" license="369535" swrid="5588601" athleteid="1624" externalid="369535">
              <RESULTS>
                <RESULT eventid="1061" points="447" swimtime="00:05:02.42" resultid="1625" heatid="2068" lane="7" entrytime="00:05:28.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                    <SPLIT distance="100" swimtime="00:01:12.29" />
                    <SPLIT distance="150" swimtime="00:01:50.48" />
                    <SPLIT distance="200" swimtime="00:02:29.34" />
                    <SPLIT distance="250" swimtime="00:03:08.29" />
                    <SPLIT distance="300" swimtime="00:03:46.67" />
                    <SPLIT distance="350" swimtime="00:04:25.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1089" points="388" swimtime="00:02:47.02" resultid="1626" heatid="2127" lane="2" entrytime="00:02:49.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                    <SPLIT distance="100" swimtime="00:01:22.56" />
                    <SPLIT distance="150" swimtime="00:02:10.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="329" swimtime="00:01:30.27" resultid="1627" heatid="2145" lane="4" entrytime="00:01:36.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Luisa Lottermann" birthdate="2011-08-26" gender="F" nation="BRA" license="382238" swrid="5596909" athleteid="1628" externalid="382238">
              <RESULTS>
                <RESULT eventid="1089" points="301" swimtime="00:03:01.64" resultid="1629" heatid="2126" lane="5" entrytime="00:03:05.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.72" />
                    <SPLIT distance="100" swimtime="00:01:34.26" />
                    <SPLIT distance="150" swimtime="00:02:21.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="311" swimtime="00:00:41.83" resultid="1630" heatid="2106" lane="3" entrytime="00:00:43.72" entrycourse="SCM" />
                <RESULT eventid="1103" points="346" swimtime="00:01:28.78" resultid="1631" heatid="2146" lane="4" entrytime="00:01:30.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Vieira Rohnelt" birthdate="2012-05-03" gender="M" nation="BRA" license="365692" swrid="5588952" athleteid="1612" externalid="365692">
              <RESULTS>
                <RESULT eventid="1071" points="145" swimtime="00:00:41.35" resultid="1613" heatid="2092" lane="6" entrytime="00:00:40.19" entrycourse="SCM" />
                <RESULT eventid="1083" points="155" swimtime="00:00:46.44" resultid="1614" heatid="2110" lane="7" entrytime="00:00:48.53" entrycourse="SCM" />
                <RESULT eventid="1105" points="153" swimtime="00:01:43.30" resultid="1615" heatid="2149" lane="7" entrytime="00:01:41.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="CVEL-SANTA MARIA, C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1077" points="284" swimtime="00:02:24.71" resultid="1632" heatid="2100" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                    <SPLIT distance="100" swimtime="00:01:13.53" />
                    <SPLIT distance="150" swimtime="00:01:50.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1620" number="1" />
                    <RELAYPOSITION athleteid="1616" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1624" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1612" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="15560" nation="BRA" region="PR" clubid="1164" name="Colégio Adventista Centenário, Curitiba" shortname="Ctba-Adven.Centen.,C">
          <ATHLETES>
            <ATHLETE firstname="Benjamin" lastname="Leao Silva" birthdate="2011-08-25" gender="M" nation="BRA" license="V413870" athleteid="1165" externalid="V413870">
              <RESULTS>
                <RESULT eventid="1075" status="RJC" swimtime="00:00:00.00" resultid="1166" />
                <RESULT eventid="1071" status="RJC" swimtime="00:00:00.00" resultid="1167" />
                <RESULT eventid="1063" points="124" swimtime="00:00:40.35" resultid="1168" heatid="2073" lane="8" />
                <RESULT eventid="1087" points="103" swimtime="00:01:35.63" resultid="1169" heatid="2119" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="99" swimtime="00:07:38.11" resultid="1170" heatid="2102" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                    <SPLIT distance="100" swimtime="00:01:36.96" />
                    <SPLIT distance="150" swimtime="00:02:36.92" />
                    <SPLIT distance="200" swimtime="00:03:37.71" />
                    <SPLIT distance="250" swimtime="00:04:38.74" />
                    <SPLIT distance="300" swimtime="00:05:39.08" />
                    <SPLIT distance="350" swimtime="00:06:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" status="RJC" swimtime="00:00:00.00" resultid="1171" />
                <RESULT eventid="1101" status="RJC" swimtime="00:00:00.00" resultid="1172" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="12397" nation="BRA" region="PR" clubid="1700" name="Colégio Imperatriz Dona Leopoldina, Guarapuava" shortname="Grpa-Imp.Leopoldi.,C">
          <ATHLETES>
            <ATHLETE firstname="Ana" lastname="Teresa Leh Sander" birthdate="2010-02-16" gender="F" nation="BRA" license="V399525" athleteid="1701" externalid="V399525">
              <RESULTS>
                <RESULT eventid="1085" points="178" swimtime="00:01:29.18" resultid="1702" heatid="2113" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1089" points="163" swimtime="00:03:42.63" resultid="1703" heatid="2125" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.19" />
                    <SPLIT distance="100" swimtime="00:01:42.82" />
                    <SPLIT distance="150" swimtime="00:02:47.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="145" swimtime="00:01:58.59" resultid="1704" heatid="2144" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Moreira Malucelli" birthdate="2012-08-09" gender="F" nation="BRA" license="V413842" athleteid="1705" externalid="V413842">
              <RESULTS>
                <RESULT eventid="1069" status="DNS" swimtime="00:00:00.00" resultid="1706" heatid="2087" lane="4" />
                <RESULT eventid="1073" status="DNS" swimtime="00:00:00.00" resultid="1707" heatid="2094" lane="2" />
                <RESULT eventid="1085" status="DNS" swimtime="00:00:00.00" resultid="1708" heatid="2113" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18858" nation="BRA" region="PR" clubid="2001" name="Escola Brasileirinho, Santa Cruz De Monte Castelo" shortname="Scmc-Brasileirinho,E">
          <ATHLETES>
            <ATHLETE firstname="Vitor" lastname="Verone Neto" birthdate="2011-11-30" gender="M" nation="BRA" license="V413930" athleteid="2002" externalid="V413930">
              <RESULTS>
                <RESULT eventid="1063" points="134" swimtime="00:00:39.32" resultid="2003" heatid="2072" lane="4" />
                <RESULT eventid="1087" points="95" swimtime="00:01:37.97" resultid="2004" heatid="2121" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17690" nation="BRA" region="PR" clubid="1931" name="6º Colégio Da Polícia Militar, Pato Branco" shortname="Pcbo-6ºcpm,C">
          <ATHLETES>
            <ATHLETE firstname="Isadora" lastname="Scariot Amorim" birthdate="2012-02-16" gender="F" nation="BRA" license="V413864" athleteid="1932" externalid="V413864">
              <RESULTS>
                <RESULT eventid="1065" points="160" swimtime="00:00:42.17" resultid="1933" heatid="2078" lane="2" />
                <RESULT eventid="1081" points="148" swimtime="00:00:53.53" resultid="1934" heatid="2104" lane="6" />
                <RESULT eventid="1099" points="128" swimtime="00:00:50.07" resultid="1935" heatid="2136" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Paula" lastname="Piassa" birthdate="2012-07-18" gender="F" nation="BRA" license="V413865" athleteid="1936" externalid="V413865">
              <RESULTS>
                <RESULT eventid="1065" points="115" swimtime="00:00:47.03" resultid="1937" heatid="2080" lane="1" />
                <RESULT eventid="1099" status="DSQ" swimtime="00:00:53.38" resultid="1938" heatid="2136" lane="1" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="877" nation="BRA" region="PR" clubid="1209" name="Colégio Bom Jesus Divina Providência, Curitiba" shortname="Ctba-Bj Divina,C">
          <ATHLETES>
            <ATHLETE firstname="Antonia" lastname="Adam  Fracaro" birthdate="2010-04-27" gender="F" nation="BRA" license="382212" swrid="5588512" athleteid="1210" externalid="382212">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="1211" heatid="2068" lane="8" entrytime="00:05:37.79" entrycourse="SCM" />
                <RESULT eventid="1065" status="DNS" swimtime="00:00:00.00" resultid="1212" heatid="2078" lane="3" entrytime="00:00:33.28" entrycourse="SCM" />
                <RESULT eventid="1085" status="DNS" swimtime="00:00:00.00" resultid="1213" heatid="2116" lane="6" entrytime="00:01:12.04" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15625" nation="BRA" region="PR" clubid="1655" name="Colégio Estadual Dr Arnaldo Busatto, Foz Do Iguaçu" shortname="Fozi-Arnaldo Bus.,Ce">
          <ATHLETES>
            <ATHLETE firstname="Pedro" lastname="Resende Ames" birthdate="2010-02-02" gender="M" nation="BRA" license="365505" swrid="5588876" athleteid="1656" externalid="365505" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1067" points="343" swimtime="00:01:08.98" resultid="1657" heatid="2086" lane="4" entrytime="00:01:05.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="427" swimtime="00:00:59.51" resultid="1658" heatid="2124" lane="2" entrytime="00:01:02.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="357" swimtime="00:00:31.15" resultid="1659" heatid="2143" lane="4" entrytime="00:00:32.52" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15627" nation="BRA" region="PR" clubid="1685" name="Colégio Estadual Profº Flávio Warken, Foz Do Iguaç" shortname="Fozi-Flávio Wark.,Ce">
          <ATHLETES>
            <ATHLETE firstname="Leticia" lastname="Marques Lima" birthdate="2010-04-30" gender="F" nation="BRA" license="383051" swrid="5596913" athleteid="1686" externalid="383051">
              <RESULTS>
                <RESULT eventid="1069" points="318" swimtime="00:01:20.40" resultid="1687" heatid="2089" lane="3" entrytime="00:01:19.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1089" points="299" swimtime="00:03:02.20" resultid="1688" heatid="2126" lane="3" entrytime="00:03:08.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                    <SPLIT distance="100" swimtime="00:01:22.79" />
                    <SPLIT distance="150" swimtime="00:02:18.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="245" swimtime="00:01:26.27" resultid="1689" heatid="2131" lane="7" entrytime="00:01:26.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1921" nation="BRA" region="PR" clubid="1881" name="Colégio Objetivo, Maringá" shortname="Mrga-Objetivo,C">
          <ATHLETES>
            <ATHLETE firstname="Tiago" lastname="Ficher Delmont Pais" birthdate="2010-07-15" gender="M" nation="BRA" license="338533" swrid="5588701" athleteid="1882" externalid="338533">
              <RESULTS>
                <RESULT eventid="1071" points="504" swimtime="00:00:27.33" resultid="1883" heatid="2093" lane="4" entrytime="00:00:27.98" entrycourse="SCM" />
                <RESULT eventid="1087" points="521" swimtime="00:00:55.70" resultid="1884" heatid="2124" lane="4" entrytime="00:00:56.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="470" swimtime="00:01:01.42" resultid="1885" heatid="2133" lane="4" entrytime="00:01:02.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17708" nation="BRA" region="PR" clubid="1478" name="Colégio Positivo Água Verde, Curitiba" shortname="Ctba-Posi. A.Verde,C">
          <ATHLETES>
            <ATHLETE firstname="Isabela" lastname="Mattioli" birthdate="2011-10-22" gender="F" nation="BRA" license="366896" swrid="5602559" athleteid="1479" externalid="366896">
              <RESULTS>
                <RESULT eventid="1065" points="397" swimtime="00:00:31.18" resultid="1480" heatid="2083" lane="8" entrytime="00:00:31.64" entrycourse="SCM" />
                <RESULT eventid="1089" points="409" swimtime="00:02:44.10" resultid="1481" heatid="2127" lane="1" entrytime="00:02:51.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.20" />
                    <SPLIT distance="100" swimtime="00:01:21.69" />
                    <SPLIT distance="150" swimtime="00:02:07.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="431" swimtime="00:01:22.54" resultid="2066" heatid="2146" lane="5" entrytime="00:01:31.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6577" nation="BRA" region="PR" clubid="1811" name="Colégio Dom Bosco, Maringá" shortname="Mrga-Dom Bosco,C">
          <ATHLETES>
            <ATHLETE firstname="Rafael" lastname="Pacheco" birthdate="2012-10-03" gender="M" nation="BRA" license="370663" swrid="5603883" athleteid="1812" externalid="370663">
              <RESULTS>
                <RESULT eventid="1071" points="253" swimtime="00:00:34.37" resultid="1813" heatid="2092" lane="5" entrytime="00:00:37.83" entrycourse="SCM" />
                <RESULT eventid="1087" points="228" swimtime="00:01:13.39" resultid="1814" heatid="2122" lane="4" entrytime="00:01:14.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="163" swimtime="00:00:40.43" resultid="1815" heatid="2142" lane="7" entrytime="00:00:41.22" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Sol Reolon Gomes" birthdate="2011-02-28" gender="F" nation="BRA" license="392100" swrid="5603914" athleteid="1816" externalid="392100">
              <RESULTS>
                <RESULT eventid="1065" points="435" swimtime="00:00:30.25" resultid="1817" heatid="2083" lane="1" entrytime="00:00:31.13" entrycourse="SCM" />
                <RESULT eventid="1085" points="391" swimtime="00:01:08.71" resultid="1818" heatid="2116" lane="3" entrytime="00:01:11.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="338" swimtime="00:00:36.24" resultid="1819" heatid="2138" lane="8" entrytime="00:00:38.80" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Furuchi Martins" birthdate="2011-10-05" gender="F" nation="BRA" license="367001" swrid="5602616" athleteid="1820" externalid="367001">
              <RESULTS>
                <RESULT eventid="1081" points="266" swimtime="00:00:44.08" resultid="1821" heatid="2106" lane="8" entrytime="00:00:45.33" entrycourse="SCM" />
                <RESULT eventid="1103" points="276" swimtime="00:01:35.76" resultid="1822" heatid="2146" lane="3" entrytime="00:01:34.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2653" nation="BRA" region="PR" clubid="1529" name="Escola Seb Dom Bosco Batel, Curitiba" shortname="Ctba-Seb Batel,E">
          <ATHLETES>
            <ATHLETE firstname="Gabriela" lastname="Cristina Ferreira" birthdate="2011-08-24" gender="F" nation="BRA" license="358334" swrid="5588611" athleteid="1530" externalid="358334">
              <RESULTS>
                <RESULT eventid="1073" points="573" swimtime="00:00:29.35" resultid="1531" heatid="2096" lane="4" entrytime="00:00:30.01" entrycourse="SCM" />
                <RESULT eventid="1089" points="583" swimtime="00:02:25.83" resultid="1532" heatid="2127" lane="4" entrytime="00:02:32.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                    <SPLIT distance="100" swimtime="00:01:08.68" />
                    <SPLIT distance="150" swimtime="00:01:51.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="617" swimtime="00:01:03.46" resultid="1533" heatid="2131" lane="4" entrytime="00:01:04.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18819" nation="BRA" region="PR" clubid="2005" name="Colégio Estadual Maurício Ferraz Da Costa, Sjpi" shortname="Sjpi-M.Ferraz,Ce">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Tomaz Zmievski" birthdate="2012-09-20" gender="F" nation="BRA" license="406725" swrid="5717300" athleteid="2006" externalid="406725">
              <RESULTS>
                <RESULT eventid="1073" points="109" swimtime="00:00:50.98" resultid="2007" heatid="2095" lane="7" entrytime="00:00:48.12" entrycourse="SCM" />
                <RESULT eventid="1065" points="219" swimtime="00:00:38.00" resultid="2008" heatid="2080" lane="3" entrytime="00:00:39.51" entrycourse="SCM" />
                <RESULT eventid="1085" points="213" swimtime="00:01:24.11" resultid="2009" heatid="2114" lane="3" entrytime="00:01:25.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3699" nation="BRA" region="PR" clubid="1524" name="Escola Seb Dom Bosco Ahú, Curitiba" shortname="Ctba-Seb Ahú,E">
          <ATHLETES>
            <ATHLETE firstname="Leonardo" lastname="Bernardi Iurk" birthdate="2012-04-14" gender="M" nation="BRA" license="406940" swrid="5717245" athleteid="1525" externalid="406940">
              <RESULTS>
                <RESULT eventid="1063" points="182" swimtime="00:00:35.55" resultid="1526" heatid="2074" lane="1" entrytime="00:00:34.65" entrycourse="SCM" />
                <RESULT eventid="1087" points="175" swimtime="00:01:20.11" resultid="1527" heatid="2122" lane="6" entrytime="00:01:19.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="120" swimtime="00:00:44.79" resultid="1528" heatid="2141" lane="4" entrytime="00:00:45.48" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16305" nation="BRA" region="PR" clubid="1178" name="Colégio Amplação, Curitiba" shortname="Ctba-Amplação,C">
          <ATHLETES>
            <ATHLETE firstname="Lauren" lastname="Dziura" birthdate="2010-01-11" gender="F" nation="BRA" license="369416" swrid="5588668" athleteid="1179" externalid="369416">
              <RESULTS>
                <RESULT eventid="1061" points="403" swimtime="00:05:12.94" resultid="1180" heatid="2068" lane="3" entrytime="00:05:21.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:14.15" />
                    <SPLIT distance="150" swimtime="00:01:52.92" />
                    <SPLIT distance="200" swimtime="00:02:32.43" />
                    <SPLIT distance="250" swimtime="00:03:12.36" />
                    <SPLIT distance="300" swimtime="00:03:53.21" />
                    <SPLIT distance="350" swimtime="00:04:33.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1089" points="342" swimtime="00:02:54.14" resultid="1181" heatid="2126" lane="4" entrytime="00:02:57.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                    <SPLIT distance="100" swimtime="00:01:24.02" />
                    <SPLIT distance="150" swimtime="00:02:15.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="258" swimtime="00:01:37.91" resultid="1182" heatid="2145" lane="6" entrytime="00:01:41.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="799" nation="BRA" region="PR" clubid="1855" name="Colégio Mater Dei, Maringá" shortname="Mrga-Mater Dei,C">
          <ATHLETES>
            <ATHLETE firstname="Caio" lastname="Garcia Cavalcante" birthdate="2011-11-21" gender="M" nation="BRA" license="378200" swrid="5603840" athleteid="1856" externalid="378200">
              <RESULTS>
                <RESULT eventid="1087" points="264" swimtime="00:01:09.87" resultid="1857" heatid="2122" lane="5" entrytime="00:01:15.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="240" swimtime="00:00:40.11" resultid="1858" heatid="2111" lane="1" entrytime="00:00:41.15" entrycourse="SCM" />
                <RESULT eventid="1105" points="238" swimtime="00:01:29.13" resultid="1859" heatid="2150" lane="1" entrytime="00:01:25.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diogo" lastname="Sanchez" birthdate="2012-11-29" gender="M" nation="BRA" license="370658" swrid="5603906" athleteid="1860" externalid="370658">
              <RESULTS>
                <RESULT eventid="1063" points="136" swimtime="00:00:39.16" resultid="1861" heatid="2073" lane="5" entrytime="00:00:36.70" entrycourse="SCM" />
                <RESULT eventid="1083" points="142" swimtime="00:00:47.75" resultid="1862" heatid="2110" lane="2" entrytime="00:00:45.67" entrycourse="SCM" />
                <RESULT eventid="1105" points="144" swimtime="00:01:45.40" resultid="1863" heatid="2149" lane="1" entrytime="00:01:42.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13349" nation="BRA" region="PR" clubid="1196" name="Colégio Bom Jesus Centro, Curitiba" shortname="Ctba-Bj Centro,C">
          <ATHLETES>
            <ATHLETE firstname="Luiza" lastname="Muxfeldt" birthdate="2011-05-13" gender="F" nation="BRA" license="366903" swrid="5602563" athleteid="1197" externalid="366903">
              <RESULTS>
                <RESULT eventid="1065" points="350" swimtime="00:00:32.53" resultid="1198" heatid="2082" lane="7" entrytime="00:00:33.87" entrycourse="SCM" />
                <RESULT eventid="1085" points="362" swimtime="00:01:10.45" resultid="1199" heatid="2116" lane="5" entrytime="00:01:09.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="299" swimtime="00:00:42.38" resultid="1200" heatid="2106" lane="7" entrytime="00:00:45.20" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rene" lastname="Osternack Erbe" birthdate="2011-04-03" gender="M" nation="BRA" license="366907" swrid="5588842" athleteid="1201" externalid="366907">
              <RESULTS>
                <RESULT eventid="1067" points="231" swimtime="00:01:18.70" resultid="1202" heatid="2085" lane="8" entrytime="00:01:20.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="214" swimtime="00:03:03.05" resultid="1203" heatid="2098" lane="3" entrytime="00:03:00.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.98" />
                    <SPLIT distance="100" swimtime="00:01:28.55" />
                    <SPLIT distance="150" swimtime="00:02:23.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="285" swimtime="00:00:30.60" resultid="1204" heatid="2075" lane="1" entrytime="00:00:31.14" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isaac" lastname="Moreira Cury De Deus" birthdate="2012-06-19" gender="M" nation="BRA" license="V413898" athleteid="1205" externalid="V413898">
              <RESULTS>
                <RESULT eventid="1071" status="WDR" swimtime="00:00:00.00" resultid="1206" />
                <RESULT eventid="1063" status="WDR" swimtime="00:00:00.00" resultid="1207" />
                <RESULT eventid="1087" status="WDR" swimtime="00:00:00.00" resultid="1208" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13940" nation="BRA" region="PR" clubid="1404" name="Colégio Madalena Sofia, Curitiba/Pr" shortname="Ctba-Madalena Sof.,C">
          <ATHLETES>
            <ATHLETE firstname="Bianca" lastname="Zanchetta Silva" birthdate="2010-08-05" gender="F" nation="BRA" license="406865" swrid="5717308" athleteid="1409" externalid="406865">
              <RESULTS>
                <RESULT eventid="1065" points="221" swimtime="00:00:37.87" resultid="1410" heatid="2080" lane="2" entrytime="00:00:42.17" entrycourse="SCM" />
                <RESULT eventid="1085" points="193" swimtime="00:01:26.89" resultid="1411" heatid="2114" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="173" swimtime="00:00:45.24" resultid="1412" heatid="2136" lane="4" entrytime="00:00:54.13" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Sieck" birthdate="2011-01-20" gender="F" nation="BRA" license="382234" swrid="5602584" athleteid="1405" externalid="382234">
              <RESULTS>
                <RESULT eventid="1073" points="182" swimtime="00:00:42.97" resultid="1406" heatid="2095" lane="3" entrytime="00:00:46.85" entrycourse="SCM" />
                <RESULT eventid="1065" points="238" swimtime="00:00:36.99" resultid="1407" heatid="2081" lane="1" entrytime="00:00:38.10" entrycourse="SCM" />
                <RESULT eventid="1095" points="153" swimtime="00:01:40.91" resultid="1408" heatid="2130" lane="6" entrytime="00:01:48.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15591" nation="BRA" region="PR" clubid="1752" name="Colégio Vila Militar (Feitep), Maringá" shortname="Mgra-Vila Militar,C">
          <ATHLETES>
            <ATHLETE firstname="Caio" lastname="Braga" birthdate="2010-05-07" gender="M" nation="BRA" license="378345" swrid="5343953" athleteid="1753" externalid="378345">
              <RESULTS>
                <RESULT eventid="1063" points="300" swimtime="00:00:30.10" resultid="1754" heatid="2075" lane="4" entrytime="00:00:29.36" entrycourse="SCM" />
                <RESULT eventid="1083" points="406" swimtime="00:00:33.67" resultid="1755" heatid="2111" lane="4" entrytime="00:00:35.12" entrycourse="SCM" />
                <RESULT eventid="1105" points="429" swimtime="00:01:13.25" resultid="1756" heatid="2150" lane="4" entrytime="00:01:13.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17664" nation="BRA" region="PR" clubid="1601" name="Colégio Passo Certo Growing, Cascavel" shortname="Cvel-Passo Certo G,C">
          <ATHLETES>
            <ATHLETE firstname="Laura" lastname="Assakura" birthdate="2010-06-29" gender="F" nation="BRA" license="376473" swrid="5596868" athleteid="1602" externalid="376473">
              <RESULTS>
                <RESULT eventid="1089" points="406" swimtime="00:02:44.51" resultid="1603" heatid="2127" lane="5" entrytime="00:02:42.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.61" />
                    <SPLIT distance="100" swimtime="00:01:20.85" />
                    <SPLIT distance="150" swimtime="00:02:05.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="348" swimtime="00:00:40.33" resultid="1604" heatid="2106" lane="4" entrytime="00:00:41.39" entrycourse="SCM" />
                <RESULT eventid="1103" points="387" swimtime="00:01:25.55" resultid="1605" heatid="2147" lane="6" entrytime="00:01:24.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18809" nation="BRA" region="PR" clubid="2010" name="Colégio Adventista De Toledo" shortname="Tole-Adventista,C">
          <ATHLETES>
            <ATHLETE firstname="Heloisa" lastname="Welter Levandowski" birthdate="2011-05-06" gender="F" nation="BRA" license="380286" swrid="5652626" athleteid="2011" externalid="380286">
              <RESULTS>
                <RESULT eventid="1061" points="357" swimtime="00:05:26.05" resultid="2012" heatid="2067" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.86" />
                    <SPLIT distance="100" swimtime="00:01:15.24" />
                    <SPLIT distance="150" swimtime="00:01:55.83" />
                    <SPLIT distance="200" swimtime="00:02:37.41" />
                    <SPLIT distance="250" swimtime="00:03:19.64" />
                    <SPLIT distance="300" swimtime="00:04:01.53" />
                    <SPLIT distance="350" swimtime="00:04:44.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1073" points="315" swimtime="00:00:35.82" resultid="2013" heatid="2095" lane="4" entrytime="00:00:38.90" entrycourse="SCM" />
                <RESULT eventid="1095" points="230" swimtime="00:01:28.17" resultid="2014" heatid="2131" lane="1" entrytime="00:01:26.75" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4221" nation="BRA" region="PR" clubid="1670" name="Colégio Estadual Cataratas Do Iguaçu" shortname="Fozi-Cataratas, Ce">
          <ATHLETES>
            <ATHLETE firstname="Paulo" lastname="Antonio Sousa" birthdate="2012-03-17" gender="M" nation="BRA" license="407497" swrid="5721498" athleteid="1671" externalid="407497">
              <RESULTS>
                <RESULT eventid="1063" points="127" swimtime="00:00:40.08" resultid="1672" heatid="2073" lane="3" entrytime="00:00:38.23" entrycourse="SCM" />
                <RESULT eventid="1083" points="98" swimtime="00:00:54.04" resultid="1673" heatid="2110" lane="8" entrytime="00:00:51.56" entrycourse="SCM" />
                <RESULT eventid="1105" points="97" swimtime="00:02:00.20" resultid="1674" heatid="2149" lane="8" entrytime="00:01:55.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="623" nation="BRA" region="PR" clubid="1159" name="Colégio Vicentino Santa Cruz, Campo Mourão" shortname="Cmou-Vicen.St.Cruz,C">
          <ATHLETES>
            <ATHLETE firstname="Matheus" lastname="Franca Rebollo" birthdate="2012-09-26" gender="M" nation="BRA" license="385780" swrid="5538081" athleteid="1160" externalid="385780">
              <RESULTS>
                <RESULT eventid="1071" points="67" swimtime="00:00:53.47" resultid="1161" heatid="2091" lane="4" />
                <RESULT eventid="1063" points="101" swimtime="00:00:43.18" resultid="1162" heatid="2072" lane="5" />
                <RESULT eventid="1087" points="83" swimtime="00:01:42.42" resultid="1163" heatid="2121" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3976" nation="BRA" region="PR" clubid="1695" name="Colégio Estadual Ulysses Guimarães, Foz Do Iguaçu" shortname="Fozi-Ulysses Gui.,Ce">
          <ATHLETES>
            <ATHLETE firstname="Leonardo" lastname="Carvalho Carelli" birthdate="2011-10-15" gender="M" nation="BRA" license="403146" swrid="5676300" athleteid="1696" externalid="403146" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1071" points="292" swimtime="00:00:32.78" resultid="1697" heatid="2092" lane="4" entrytime="00:00:37.38" entrycourse="SCM" />
                <RESULT eventid="1063" points="296" swimtime="00:00:30.25" resultid="1698" heatid="2074" lane="4" entrytime="00:00:31.73" entrycourse="SCM" />
                <RESULT eventid="1097" points="294" swimtime="00:01:11.81" resultid="1699" heatid="2133" lane="2" entrytime="00:01:14.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18856" nation="BRA" region="PR" clubid="1390" name="Escola Interativa, Curitiba" shortname="Ctba-Interativa,E">
          <ATHLETES>
            <ATHLETE firstname="Otto" lastname="Hedeke" birthdate="2011-03-24" gender="M" nation="BRA" license="372643" swrid="5588738" athleteid="1391" externalid="372643">
              <RESULTS>
                <RESULT eventid="1075" points="189" swimtime="00:03:10.94" resultid="1392" heatid="2098" lane="1" entrytime="00:03:13.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.61" />
                    <SPLIT distance="100" swimtime="00:01:32.96" />
                    <SPLIT distance="150" swimtime="00:02:29.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="249" swimtime="00:05:37.11" resultid="1393" heatid="2103" lane="8" entrytime="00:05:35.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                    <SPLIT distance="100" swimtime="00:01:20.33" />
                    <SPLIT distance="150" swimtime="00:02:03.35" />
                    <SPLIT distance="200" swimtime="00:02:46.48" />
                    <SPLIT distance="250" swimtime="00:03:29.92" />
                    <SPLIT distance="300" swimtime="00:04:14.50" />
                    <SPLIT distance="350" swimtime="00:04:58.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="175" swimtime="00:01:38.73" resultid="1394" heatid="2148" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18850" nation="BRA" region="PR" clubid="1828" name="Colégio Interação, Maringá" shortname="Mrga-Interação,C">
          <ATHLETES>
            <ATHLETE firstname="Theo" lastname="Rossi" birthdate="2012-05-21" gender="M" nation="BRA" license="378346" swrid="5603901" athleteid="1829" externalid="378346">
              <RESULTS>
                <RESULT eventid="1071" status="DNS" swimtime="00:00:00.00" resultid="1830" heatid="2092" lane="7" />
                <RESULT eventid="1063" status="DNS" swimtime="00:00:00.00" resultid="1831" heatid="2074" lane="2" entrytime="00:00:33.12" entrycourse="SCM" />
                <RESULT eventid="1101" points="180" swimtime="00:00:39.11" resultid="1832" heatid="2142" lane="5" entrytime="00:00:38.49" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edgar" lastname="Romero" birthdate="2011-05-12" gender="M" nation="BRA" license="V413920" athleteid="1833" externalid="V413920">
              <RESULTS>
                <RESULT eventid="1063" points="233" swimtime="00:00:32.74" resultid="1834" heatid="2070" lane="4" />
                <RESULT eventid="1087" points="241" swimtime="00:01:12.02" resultid="1835" heatid="2120" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18822" nation="BRA" region="PR" clubid="1112" name="Colégio Presbiteriano Chamberlain, Apucarana" shortname="Apuc-Chamberlain,C">
          <ATHLETES>
            <ATHLETE firstname="Jesse" lastname="Duarte Luchtemberg" birthdate="2010-11-05" gender="M" nation="BRA" license="V413929" athleteid="1113" externalid="V413929">
              <RESULTS>
                <RESULT eventid="1063" status="DNS" swimtime="00:00:00.00" resultid="1114" heatid="2072" lane="7" />
                <RESULT eventid="1101" status="DNS" swimtime="00:00:00.00" resultid="1115" heatid="2139" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18863" nation="BRA" region="PR" clubid="2015" name="Colégio Estadual Jardim Gisella, Toledo" shortname="Tole-Jard. Gisella,C">
          <ATHLETES>
            <ATHLETE firstname="Kawan" lastname="Gustavo Klein Ladeia" birthdate="2010-04-19" gender="M" nation="BRA" license="V413943" athleteid="2016" externalid="V413943">
              <RESULTS>
                <RESULT eventid="1063" points="235" swimtime="00:00:32.63" resultid="2017" heatid="2072" lane="8" />
                <RESULT eventid="1087" points="200" swimtime="00:01:16.64" resultid="2018" heatid="2118" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="166" swimtime="00:00:45.34" resultid="2019" heatid="2108" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2632" nation="BRA" region="PR" clubid="1459" name="Colégio Nossa Senhora Medianeira, Curitiba" shortname="Ctba-Medianeira,C">
          <ATHLETES>
            <ATHLETE firstname="Martina" lastname="Mayer Paludetto" birthdate="2012-10-30" gender="F" nation="BRA" license="369264" swrid="5588811" athleteid="1460" externalid="369264">
              <RESULTS>
                <RESULT eventid="1065" points="410" swimtime="00:00:30.85" resultid="1461" heatid="2083" lane="3" entrytime="00:00:29.80" entrycourse="SCM" />
                <RESULT eventid="1089" points="354" swimtime="00:02:52.14" resultid="1462" heatid="2127" lane="6" entrytime="00:02:48.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                    <SPLIT distance="100" swimtime="00:01:22.26" />
                    <SPLIT distance="150" swimtime="00:02:13.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="254" swimtime="00:01:25.24" resultid="1463" heatid="2131" lane="8" entrytime="00:01:29.57" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1994" nation="BRA" region="PR" clubid="1633" name="Colégio Anglo Americano, Foz Do Iguaçu" shortname="Fozi-Ang.Americano,C">
          <ATHLETES>
            <ATHLETE firstname="Katherine" lastname="Kotz" birthdate="2012-05-18" gender="F" nation="BRA" license="390810" swrid="5596907" athleteid="1634" externalid="390810" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1065" status="DNS" swimtime="00:00:00.00" resultid="1635" heatid="2082" lane="6" entrytime="00:00:32.56" entrycourse="SCM" />
                <RESULT eventid="1085" status="DNS" swimtime="00:00:00.00" resultid="1636" heatid="2115" lane="4" entrytime="00:01:12.81" entrycourse="SCM" />
                <RESULT eventid="1081" status="DNS" swimtime="00:00:00.00" resultid="1637" heatid="2106" lane="1" entrytime="00:00:45.32" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Leticia Sbardelatti" birthdate="2011-07-28" gender="F" nation="BRA" license="403147" swrid="5676303" athleteid="1638" externalid="403147" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1061" points="234" swimtime="00:06:15.21" resultid="1639" heatid="2067" lane="3" entrytime="00:07:39.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                    <SPLIT distance="100" swimtime="00:01:28.15" />
                    <SPLIT distance="150" swimtime="00:02:15.99" />
                    <SPLIT distance="200" swimtime="00:03:03.76" />
                    <SPLIT distance="250" swimtime="00:03:51.98" />
                    <SPLIT distance="300" swimtime="00:04:40.54" />
                    <SPLIT distance="350" swimtime="00:05:29.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="264" swimtime="00:00:35.73" resultid="1640" heatid="2081" lane="3" entrytime="00:00:36.77" entrycourse="SCM" />
                <RESULT eventid="1085" points="227" swimtime="00:01:22.33" resultid="1641" heatid="2115" lane="1" entrytime="00:01:22.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Gabriel Dreher" birthdate="2011-12-05" gender="M" nation="BRA" license="403148" swrid="5676302" athleteid="1642" externalid="403148" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1067" points="163" swimtime="00:01:28.46" resultid="1643" heatid="2084" lane="5" entrytime="00:01:35.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="166" swimtime="00:01:21.47" resultid="1644" heatid="2122" lane="7" entrytime="00:01:24.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="200" swimtime="00:06:02.61" resultid="1645" heatid="2101" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.31" />
                    <SPLIT distance="100" swimtime="00:01:25.97" />
                    <SPLIT distance="150" swimtime="00:02:13.57" />
                    <SPLIT distance="200" swimtime="00:03:01.39" />
                    <SPLIT distance="250" swimtime="00:03:44.00" />
                    <SPLIT distance="300" swimtime="00:04:30.26" />
                    <SPLIT distance="350" swimtime="00:05:17.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Lima Belo" birthdate="2012-10-07" gender="F" nation="BRA" license="407799" swrid="5721502" athleteid="1646" externalid="407799">
              <RESULTS>
                <RESULT eventid="1065" points="156" swimtime="00:00:42.58" resultid="1647" heatid="2080" lane="8" />
                <RESULT eventid="1085" points="122" swimtime="00:01:41.27" resultid="1648" heatid="2114" lane="7" entrytime="00:01:54.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="89" swimtime="00:01:03.42" resultid="1649" heatid="2105" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Marcio Peixoto" birthdate="2012-10-22" gender="M" nation="BRA" license="411994" swrid="5740013" athleteid="1650" externalid="411994">
              <RESULTS>
                <RESULT eventid="1063" points="130" swimtime="00:00:39.70" resultid="1651" heatid="2071" lane="5" />
                <RESULT eventid="1087" points="127" swimtime="00:01:29.05" resultid="1652" heatid="2120" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="79" swimtime="00:00:51.48" resultid="1653" heatid="2140" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="FOZI-ANG.AMERICANO,C" number="1">
              <RESULTS>
                <RESULT eventid="1077" status="DSQ" swimtime="00:03:07.44" resultid="1654" heatid="2100" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.73" />
                    <SPLIT distance="100" swimtime="00:01:43.30" />
                    <SPLIT distance="150" swimtime="00:02:27.80" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1642" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="1646" number="2" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1638" number="3" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1650" number="4" reactiontime="0" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="6593" nation="BRA" region="PR" clubid="1864" name="Escola Notre Dame, Maringá" shortname="Mrga-Notre Dame,E">
          <ATHLETES>
            <ATHLETE firstname="Isadora" lastname="Mochiutti Carneiro" birthdate="2010-04-22" gender="F" nation="BRA" license="370670" swrid="5588817" athleteid="1865" externalid="370670">
              <RESULTS>
                <RESULT eventid="1073" points="443" swimtime="00:00:31.98" resultid="1866" heatid="2096" lane="3" entrytime="00:00:33.29" entrycourse="SCM" />
                <RESULT eventid="1085" points="487" swimtime="00:01:03.84" resultid="1867" heatid="2117" lane="3" entrytime="00:01:05.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="409" swimtime="00:01:12.77" resultid="1868" heatid="2131" lane="3" entrytime="00:01:13.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Kenji Yamaguchi" birthdate="2011-08-25" gender="M" nation="BRA" license="385708" swrid="5603862" athleteid="1869" externalid="385708">
              <RESULTS>
                <RESULT eventid="1087" points="237" swimtime="00:01:12.43" resultid="1870" heatid="2123" lane="8" entrytime="00:01:11.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="262" swimtime="00:01:14.63" resultid="1871" heatid="2132" lane="3" entrytime="00:01:19.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="222" swimtime="00:01:31.24" resultid="1872" heatid="2149" lane="6" entrytime="00:01:31.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Moreschi" birthdate="2012-08-09" gender="M" nation="BRA" license="385715" swrid="5603876" athleteid="1873" externalid="385715">
              <RESULTS>
                <RESULT eventid="1075" points="177" swimtime="00:03:15.10" resultid="1874" heatid="2098" lane="2" entrytime="00:03:04.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.52" />
                    <SPLIT distance="100" swimtime="00:01:35.99" />
                    <SPLIT distance="150" swimtime="00:02:31.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="171" swimtime="00:00:44.89" resultid="1875" heatid="2110" lane="5" entrytime="00:00:43.33" entrycourse="SCM" />
                <RESULT eventid="1105" status="DNS" swimtime="00:00:00.00" resultid="1876" heatid="2149" lane="2" entrytime="00:01:34.81" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Jacobsen Donati" birthdate="2011-07-14" gender="M" nation="BRA" license="391851" swrid="5615735" athleteid="1877" externalid="391851">
              <RESULTS>
                <RESULT eventid="1067" points="294" swimtime="00:01:12.62" resultid="1878" heatid="2086" lane="8" entrytime="00:01:12.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="359" swimtime="00:00:28.34" resultid="1879" heatid="2076" lane="8" entrytime="00:00:29.34" entrycourse="SCM" />
                <RESULT eventid="1087" points="376" swimtime="00:01:02.11" resultid="1880" heatid="2124" lane="7" entrytime="00:01:03.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18861" nation="BRA" region="PR" clubid="1714" name="Colégio Estadual Presidente Roosevelt, Guaira" shortname="Guai-Roosevelt,Ce">
          <ATHLETES>
            <ATHLETE firstname="Leonardo" lastname="Makoto Isigaki" birthdate="2011-04-09" gender="M" nation="BRA" license="V413945" athleteid="1718" externalid="V413945">
              <RESULTS>
                <RESULT eventid="1063" points="52" swimtime="00:00:53.84" resultid="1719" heatid="2071" lane="2" />
                <RESULT eventid="1083" status="DSQ" swimtime="00:01:08.17" resultid="1720" heatid="2109" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose" lastname="Antonio Moreira Souza" birthdate="2012-11-08" gender="M" nation="BRA" license="V413944" athleteid="1715" externalid="V413944">
              <RESULTS>
                <RESULT eventid="1063" points="42" swimtime="00:00:57.89" resultid="1716" heatid="2070" lane="3" />
                <RESULT eventid="1101" status="DSQ" swimtime="00:01:16.39" resultid="1717" heatid="2140" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="319" nation="BRA" region="PR" clubid="1116" name="Colégio São José, Apucarana" shortname="Apuc-São José,C">
          <ATHLETES>
            <ATHLETE firstname="Gustavo" lastname="Murakami Niyme" birthdate="2010-01-28" gender="M" nation="BRA" license="V413950" athleteid="1117" externalid="V413950">
              <RESULTS>
                <RESULT eventid="1063" points="188" swimtime="00:00:35.16" resultid="1118" heatid="2072" lane="2" />
                <RESULT eventid="1083" points="141" swimtime="00:00:47.87" resultid="1119" heatid="2108" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13350" nation="BRA" region="PR" clubid="1214" name="Colégio Bom Jesus Nossa Srª. De Lourdes, Curitiba" shortname="Ctba-Bj Lourdes,C">
          <ATHLETES>
            <ATHLETE firstname="Rafaelle" lastname="Matos De Souza" birthdate="2011-04-24" gender="F" nation="BRA" license="367146" athleteid="1255" externalid="367146">
              <RESULTS>
                <RESULT eventid="1065" points="266" swimtime="00:00:35.62" resultid="1256" heatid="2080" lane="5" entrytime="00:00:38.85" entrycourse="SCM" />
                <RESULT eventid="1085" points="267" swimtime="00:01:18.02" resultid="1257" heatid="2112" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="221" swimtime="00:00:41.73" resultid="1258" heatid="2137" lane="8" entrytime="00:00:46.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Iglesias Prado" birthdate="2010-06-15" gender="M" nation="BRA" license="408052" swrid="5723025" athleteid="1243" externalid="408052">
              <RESULTS>
                <RESULT eventid="1067" points="149" swimtime="00:01:31.07" resultid="1244" heatid="2084" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="203" swimtime="00:00:36.99" resultid="1245" heatid="2092" lane="8" />
                <RESULT eventid="1087" points="228" swimtime="00:01:13.30" resultid="1246" heatid="2120" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Fontoura Barros" birthdate="2011-08-04" gender="F" nation="BRA" license="403143" swrid="5676298" athleteid="1231" externalid="403143">
              <RESULTS>
                <RESULT eventid="1065" status="DNS" swimtime="00:00:00.00" resultid="1232" heatid="2080" lane="7" entrytime="00:00:43.14" entrycourse="SCM" />
                <RESULT eventid="1081" status="DNS" swimtime="00:00:00.00" resultid="1233" heatid="2104" lane="4" />
                <RESULT eventid="1103" status="DNS" swimtime="00:00:00.00" resultid="1234" heatid="2145" lane="1" entrytime="00:01:58.87" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Celli Schneider" birthdate="2011-02-21" gender="M" nation="BRA" license="367055" swrid="5588587" athleteid="1219" externalid="367055">
              <RESULTS>
                <RESULT eventid="1067" points="251" swimtime="00:01:16.55" resultid="1220" heatid="2085" lane="3" entrytime="00:01:15.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="262" swimtime="00:01:14.61" resultid="1221" heatid="2132" lane="6" entrytime="00:01:24.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="280" swimtime="00:00:33.78" resultid="1222" heatid="2143" lane="3" entrytime="00:00:33.93" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabel" lastname="Martinez Tarnowski" birthdate="2010-09-20" gender="F" nation="BRA" license="V413871" athleteid="1263" externalid="V413871">
              <RESULTS>
                <RESULT eventid="1085" points="182" swimtime="00:01:28.53" resultid="1264" heatid="2113" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="176" swimtime="00:00:50.55" resultid="1265" heatid="2104" lane="5" />
                <RESULT eventid="1103" points="164" swimtime="00:01:53.78" resultid="1266" heatid="2144" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabele" lastname="Veiga Reis" birthdate="2010-04-22" gender="F" nation="BRA" license="V383046" athleteid="1251" externalid="V383046">
              <RESULTS>
                <RESULT eventid="1061" status="DNS" swimtime="00:00:00.00" resultid="1252" heatid="2067" lane="2" />
                <RESULT eventid="1073" status="DNS" swimtime="00:00:00.00" resultid="1253" heatid="2095" lane="1" entrytime="00:00:48.69" entrycourse="SCM" />
                <RESULT eventid="1099" status="DNS" swimtime="00:00:00.00" resultid="1254" heatid="2135" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cristopher" lastname="Ribas Pinto" birthdate="2011-01-27" gender="M" nation="BRA" license="V399519" athleteid="1239" externalid="V399519">
              <RESULTS>
                <RESULT eventid="1063" points="135" swimtime="00:00:39.22" resultid="1240" heatid="2073" lane="7" entrytime="00:00:41.28" entrycourse="SCM" />
                <RESULT eventid="1087" points="121" swimtime="00:01:30.57" resultid="1241" heatid="2119" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="134" swimtime="00:00:48.65" resultid="1242" heatid="2109" lane="4" entrytime="00:00:52.49" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Cavassin Ieger" birthdate="2011-08-31" gender="M" nation="BRA" license="367149" swrid="5588743" athleteid="1227" externalid="367149">
              <RESULTS>
                <RESULT eventid="1075" points="240" swimtime="00:02:56.28" resultid="1228" heatid="2098" lane="8" entrytime="00:03:16.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:25.49" />
                    <SPLIT distance="150" swimtime="00:02:14.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="262" swimtime="00:00:38.96" resultid="1229" heatid="2111" lane="7" entrytime="00:00:40.56" entrycourse="SCM" />
                <RESULT eventid="1105" points="260" swimtime="00:01:26.61" resultid="1230" heatid="2149" lane="5" entrytime="00:01:29.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giuseppe" lastname="Marquardt Ditterich" birthdate="2012-09-27" gender="M" nation="BRA" license="V413902" athleteid="1271" externalid="V413902">
              <RESULTS>
                <RESULT eventid="1067" points="75" swimtime="00:01:54.22" resultid="1272" heatid="2084" lane="1" />
                <RESULT eventid="1063" points="79" swimtime="00:00:46.80" resultid="1273" heatid="2071" lane="1" />
                <RESULT eventid="1101" points="76" swimtime="00:00:52.17" resultid="1274" heatid="2140" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Luisa Formagini Da Silva" birthdate="2011-04-20" gender="F" nation="BRA" license="V413869" athleteid="1259" externalid="V413869">
              <RESULTS>
                <RESULT eventid="1069" status="DSQ" swimtime="00:00:00.00" resultid="1260" heatid="2087" lane="3" />
                <RESULT eventid="1065" points="186" swimtime="00:00:40.16" resultid="1261" heatid="2079" lane="5" />
                <RESULT eventid="1081" status="DNS" swimtime="00:00:00.00" resultid="1262" heatid="2105" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Kozera Chiarato" birthdate="2010-05-28" gender="M" nation="BRA" license="406722" swrid="5717275" athleteid="1247" externalid="406722">
              <RESULTS>
                <RESULT eventid="1071" points="262" swimtime="00:00:33.97" resultid="1248" heatid="2093" lane="1" entrytime="00:00:34.84" entrycourse="SCM" />
                <RESULT eventid="1083" points="202" swimtime="00:00:42.48" resultid="1249" heatid="2110" lane="4" entrytime="00:00:42.98" entrycourse="SCM" />
                <RESULT eventid="1097" points="223" swimtime="00:01:18.69" resultid="1250" heatid="2132" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="Moreira Furtado" birthdate="2011-01-27" gender="F" nation="BRA" license="403783" swrid="5684587" athleteid="1235" externalid="403783">
              <RESULTS>
                <RESULT eventid="1069" points="174" swimtime="00:01:38.32" resultid="1236" heatid="2087" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="246" swimtime="00:00:36.55" resultid="1237" heatid="2080" lane="6" entrytime="00:00:40.90" entrycourse="SCM" />
                <RESULT eventid="1085" points="255" swimtime="00:01:19.15" resultid="1238" heatid="2114" lane="2" entrytime="00:01:29.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Edward" lastname="Luiz Santiago" birthdate="2012-02-02" gender="M" nation="BRA" license="V413901" athleteid="1267" externalid="V413901">
              <RESULTS>
                <RESULT eventid="1063" points="217" swimtime="00:00:33.52" resultid="1268" heatid="2070" lane="6" />
                <RESULT eventid="1087" points="191" swimtime="00:01:17.86" resultid="1269" heatid="2121" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="153" swimtime="00:00:41.25" resultid="1270" heatid="2140" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Carneiro Silva" birthdate="2011-02-21" gender="F" nation="BRA" license="390924" swrid="5602522" athleteid="1215" externalid="390924">
              <RESULTS>
                <RESULT eventid="1069" points="305" swimtime="00:01:21.49" resultid="1216" heatid="2089" lane="6" entrytime="00:01:22.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="353" swimtime="00:01:11.10" resultid="1217" heatid="2115" lane="5" entrytime="00:01:12.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="319" swimtime="00:00:36.94" resultid="1218" heatid="2138" lane="1" entrytime="00:00:37.76" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Guizun Jannuzzi" birthdate="2011-12-27" gender="M" nation="BRA" license="367148" swrid="5588732" athleteid="1223" externalid="367148">
              <RESULTS>
                <RESULT eventid="1063" status="DNS" swimtime="00:00:00.00" resultid="1224" heatid="2074" lane="8" entrytime="00:00:34.66" entrycourse="SCM" />
                <RESULT eventid="1087" status="DNS" swimtime="00:00:00.00" resultid="1225" heatid="2121" lane="6" />
                <RESULT eventid="1083" status="DNS" swimtime="00:00:00.00" resultid="1226" heatid="2109" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CTBA-BJ LOURDES,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1091" points="288" swimtime="00:02:03.74" resultid="1277" heatid="2128" lane="4" entrytime="00:01:55.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                    <SPLIT distance="100" swimtime="00:01:03.33" />
                    <SPLIT distance="150" swimtime="00:01:34.75" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1243" number="1" />
                    <RELAYPOSITION athleteid="1227" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1247" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1219" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1109" points="247" swimtime="00:02:22.97" resultid="1278" heatid="2152" lane="4" entrytime="00:02:10.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.53" />
                    <SPLIT distance="100" swimtime="00:01:18.47" />
                    <SPLIT distance="150" swimtime="00:01:50.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1267" number="1" />
                    <RELAYPOSITION athleteid="1227" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1219" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1243" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="CTBA-BJ LOURDES,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1093" points="280" swimtime="00:02:21.32" resultid="1275" heatid="2129" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:07.89" />
                    <SPLIT distance="150" swimtime="00:01:43.91" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1215" number="1" />
                    <RELAYPOSITION athleteid="1255" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1235" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1263" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1107" points="237" swimtime="00:02:45.21" resultid="1276" heatid="2151" lane="4" entrytime="00:02:29.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:01:31.92" />
                    <SPLIT distance="150" swimtime="00:02:09.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1255" number="1" />
                    <RELAYPOSITION athleteid="1263" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1215" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1235" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="CTBA-BJ LOURDES,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1077" points="283" swimtime="00:02:24.92" resultid="1279" heatid="2100" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                    <SPLIT distance="100" swimtime="00:01:17.55" />
                    <SPLIT distance="150" swimtime="00:01:49.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1215" number="1" />
                    <RELAYPOSITION athleteid="1227" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1219" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1255" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="17655" nation="BRA" region="PR" clubid="1375" name="Colégio Imaculada Conceição, Curitiba" shortname="Ctba-IMC.Conceição,C">
          <ATHLETES>
            <ATHLETE firstname="Jhon" lastname="Caleb Dos Santos" birthdate="2010-03-02" gender="M" nation="BRA" license="359020" swrid="5588574" athleteid="1376" externalid="359020">
              <RESULTS>
                <RESULT eventid="1067" points="406" swimtime="00:01:05.22" resultid="1377" heatid="2086" lane="6" entrytime="00:01:07.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="475" swimtime="00:02:20.46" resultid="1378" heatid="2099" lane="5" entrytime="00:02:26.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                    <SPLIT distance="100" swimtime="00:01:07.26" />
                    <SPLIT distance="150" swimtime="00:01:48.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="448" swimtime="00:01:02.41" resultid="1379" heatid="2133" lane="5" entrytime="00:01:04.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16331" nation="BRA" region="PR" clubid="1757" name="4º Colégio Da Polícia Militar, Maringá" shortname="Mrga-4ºcpmpr,C">
          <ATHLETES>
            <ATHLETE firstname="Sophia" lastname="Stephany" birthdate="2012-07-27" gender="F" nation="BRA" license="382210" swrid="5603917" athleteid="1758" externalid="382210">
              <RESULTS>
                <RESULT eventid="1073" status="DNS" swimtime="00:00:00.00" resultid="1759" heatid="2095" lane="6" entrytime="00:00:46.92" entrycourse="SCM" />
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="1760" heatid="2126" lane="1" entrytime="00:03:38.27" entrycourse="SCM" />
                <RESULT eventid="1099" status="DNS" swimtime="00:00:00.00" resultid="1761" heatid="2137" lane="1" entrytime="00:00:45.29" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18838" nation="BRA" region="PR" clubid="2047" name="Colégio Estadual Pedro Marcondes Ribas, Ventania" shortname="Vent-Pedro Ribas,Ce">
          <ATHLETES>
            <ATHLETE firstname="Ana" lastname="Flavia Pinheiro De Oliveira" birthdate="2012-12-11" gender="F" nation="BRA" license="V413888" athleteid="2048" externalid="V413888">
              <RESULTS>
                <RESULT eventid="1065" status="DNS" swimtime="00:00:00.00" resultid="2049" heatid="2079" lane="8" />
                <RESULT eventid="1099" status="DNS" swimtime="00:00:00.00" resultid="2050" heatid="2136" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="739" nation="BRA" region="PR" clubid="1149" name="CCM Marechal Rondon, Campo Mourão" shortname="Cmou-Mar. Rondon,CCM">
          <ATHLETES>
            <ATHLETE firstname="Enzo" lastname="Garcia Goulart" birthdate="2010-11-29" gender="M" nation="BRA" license="V413933" athleteid="1150" externalid="V413933">
              <RESULTS>
                <RESULT eventid="1067" status="SICK" swimtime="00:00:00.00" resultid="1151" />
                <RESULT eventid="1087" status="SICK" swimtime="00:00:00.00" resultid="1152" />
                <RESULT eventid="1101" status="SICK" swimtime="00:00:00.00" resultid="1153" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6544" nation="BRA" region="PR" clubid="1132" name="CCM Dr Osvaldo Cruz, Campo Mourão" shortname="Cmou-Dr Osv.Cruz,CC">
          <ATHLETES>
            <ATHLETE firstname="Yasmin" lastname="Ferreira Batista" birthdate="2012-03-29" gender="F" nation="BRA" license="385779" swrid="5532525" athleteid="1133" externalid="385779">
              <RESULTS>
                <RESULT eventid="1065" points="217" swimtime="00:00:38.12" resultid="1134" heatid="2079" lane="1" />
                <RESULT eventid="1085" points="206" swimtime="00:01:24.99" resultid="1135" heatid="2113" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="184" swimtime="00:00:44.39" resultid="1136" heatid="2136" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="10546" nation="BRA" region="PR" clubid="1483" name="Colégio Positivo Jardim Ambiental, Curitiba" shortname="Ctba-Posi. Ambien.,C">
          <ATHLETES>
            <ATHLETE firstname="Laura" lastname="Zaroni" birthdate="2010-03-03" gender="F" nation="BRA" license="356345" swrid="5600282" athleteid="1484" externalid="356345">
              <RESULTS>
                <RESULT eventid="1081" points="400" swimtime="00:00:38.48" resultid="1485" heatid="2107" lane="5" entrytime="00:00:38.14" entrycourse="SCM" />
                <RESULT eventid="1103" points="417" swimtime="00:01:23.44" resultid="1486" heatid="2147" lane="5" entrytime="00:01:21.61" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2661" nation="BRA" region="PR" clubid="1785" name="Colégio Estadual Branca Da Mota Fernandes, Maringá" shortname="Mrga-Branca,Ce">
          <ATHLETES>
            <ATHLETE firstname="Arthur" lastname="Ayres" birthdate="2012-05-05" gender="M" nation="BRA" license="378035" swrid="5208079" athleteid="1794" externalid="378035">
              <RESULTS>
                <RESULT eventid="1067" points="269" swimtime="00:01:14.85" resultid="1795" heatid="2085" lane="5" entrytime="00:01:14.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1071" points="274" swimtime="00:00:33.48" resultid="1796" heatid="2093" lane="6" entrytime="00:00:33.20" entrycourse="SCM" />
                <RESULT eventid="1063" points="273" swimtime="00:00:31.05" resultid="1797" heatid="2075" lane="8" entrytime="00:00:31.27" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Muniz" birthdate="2012-09-03" gender="M" nation="BRA" license="392106" swrid="5603877" athleteid="1798" externalid="392106">
              <RESULTS>
                <RESULT eventid="1071" points="99" swimtime="00:00:46.95" resultid="1799" heatid="2092" lane="2" entrytime="00:00:50.79" entrycourse="SCM" />
                <RESULT eventid="1087" points="145" swimtime="00:01:25.17" resultid="1800" heatid="2122" lane="8" entrytime="00:01:29.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="100" swimtime="00:00:47.51" resultid="1801" heatid="2141" lane="5" entrytime="00:00:52.84" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Pavão" birthdate="2012-04-04" gender="F" nation="BRA" license="377259" swrid="5603888" athleteid="1786" externalid="377259">
              <RESULTS>
                <RESULT eventid="1065" points="262" swimtime="00:00:35.79" resultid="1787" heatid="2081" lane="6" entrytime="00:00:36.79" entrycourse="SCM" />
                <RESULT eventid="1089" points="228" swimtime="00:03:19.45" resultid="1788" heatid="2126" lane="2" entrytime="00:03:23.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.07" />
                    <SPLIT distance="100" swimtime="00:01:34.85" />
                    <SPLIT distance="150" swimtime="00:02:33.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="228" swimtime="00:00:41.32" resultid="1789" heatid="2137" lane="4" entrytime="00:00:41.41" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raphael" lastname="Piai Pellegrini" birthdate="2012-03-24" gender="M" nation="BRA" license="377261" swrid="5603894" athleteid="1790" externalid="377261">
              <RESULTS>
                <RESULT eventid="1071" points="287" swimtime="00:00:32.96" resultid="1791" heatid="2093" lane="3" entrytime="00:00:33.17" entrycourse="SCM" />
                <RESULT eventid="1079" points="256" swimtime="00:05:34.22" resultid="1792" heatid="2153" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:18.71" />
                    <SPLIT distance="150" swimtime="00:02:03.37" />
                    <SPLIT distance="200" swimtime="00:02:45.51" />
                    <SPLIT distance="250" swimtime="00:03:28.90" />
                    <SPLIT distance="300" swimtime="00:04:12.89" />
                    <SPLIT distance="350" swimtime="00:04:57.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="239" swimtime="00:00:35.58" resultid="1793" heatid="2141" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2603" nation="BRA" region="PR" clubid="1946" name="Colégio Sagrada Família, Ponta Grossa" shortname="Pgro-Sagrada Fami.,C">
          <ATHLETES>
            <ATHLETE firstname="Isis" lastname="Maria Simoes" birthdate="2012-10-22" gender="F" nation="BRA" license="V413868" athleteid="1970" externalid="V413868">
              <RESULTS>
                <RESULT eventid="1073" points="162" swimtime="00:00:44.66" resultid="1971" heatid="2094" lane="6" />
                <RESULT eventid="1081" points="224" swimtime="00:00:46.68" resultid="1972" heatid="2105" lane="3" />
                <RESULT eventid="1099" points="218" swimtime="00:00:41.92" resultid="1973" heatid="2136" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Derick" lastname="Vinicius Garbuio Santana" birthdate="2011-09-12" gender="M" nation="BRA" license="V413925" athleteid="1974" externalid="V413925">
              <RESULTS>
                <RESULT eventid="1063" points="158" swimtime="00:00:37.27" resultid="1975" heatid="2072" lane="3" />
                <RESULT eventid="1083" points="105" swimtime="00:00:52.73" resultid="1976" heatid="2109" lane="3" />
                <RESULT eventid="1101" points="105" swimtime="00:00:46.79" resultid="1977" heatid="2140" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Franca Berger" birthdate="2010-05-07" gender="F" nation="BRA" license="399692" swrid="5653290" athleteid="1963" externalid="399692">
              <RESULTS>
                <RESULT eventid="1073" points="134" swimtime="00:00:47.55" resultid="1964" heatid="2094" lane="5" />
                <RESULT eventid="1065" points="268" swimtime="00:00:35.54" resultid="1965" heatid="2081" lane="5" entrytime="00:00:35.83" entrycourse="SCM" />
                <RESULT eventid="1081" points="203" swimtime="00:00:48.26" resultid="1966" heatid="2106" lane="6" entrytime="00:00:44.95" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Brenda" lastname="Gabriele Carvalho" birthdate="2010-04-11" gender="F" nation="BRA" license="399557" swrid="5658060" athleteid="1951" externalid="399557">
              <RESULTS>
                <RESULT eventid="1069" points="217" swimtime="00:01:31.33" resultid="1952" heatid="2088" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="265" swimtime="00:01:18.19" resultid="1953" heatid="2115" lane="8" entrytime="00:01:22.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="179" swimtime="00:01:50.59" resultid="1954" heatid="2145" lane="3" entrytime="00:01:40.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Augusto" lastname="Tramontin" birthdate="2011-11-29" gender="M" nation="BRA" license="399691" swrid="5652901" athleteid="1959" externalid="399691">
              <RESULTS>
                <RESULT eventid="1063" points="338" swimtime="00:00:28.93" resultid="1960" heatid="2075" lane="5" entrytime="00:00:29.87" entrycourse="SCM" />
                <RESULT eventid="1083" points="274" swimtime="00:00:38.39" resultid="1961" heatid="2111" lane="8" entrytime="00:00:41.66" entrycourse="SCM" />
                <RESULT eventid="1101" points="243" swimtime="00:00:35.39" resultid="1962" heatid="2142" lane="4" entrytime="00:00:37.69" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Rodrigues Neto" birthdate="2010-07-30" gender="M" nation="BRA" license="V387186" athleteid="1947" externalid="V387186">
              <RESULTS>
                <RESULT eventid="1075" points="177" swimtime="00:03:14.93" resultid="1948" heatid="2097" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.83" />
                    <SPLIT distance="100" swimtime="00:01:30.13" />
                    <SPLIT distance="150" swimtime="00:02:31.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="199" swimtime="00:06:03.41" resultid="1949" heatid="2102" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:01:18.93" />
                    <SPLIT distance="150" swimtime="00:02:03.38" />
                    <SPLIT distance="200" swimtime="00:02:51.29" />
                    <SPLIT distance="250" swimtime="00:03:39.70" />
                    <SPLIT distance="300" swimtime="00:04:27.92" />
                    <SPLIT distance="350" swimtime="00:05:15.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="110" swimtime="00:01:39.50" resultid="1950" heatid="2132" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Fernanda Mileo" birthdate="2012-09-17" gender="F" nation="BRA" license="V413860" athleteid="1967" externalid="V413860">
              <RESULTS>
                <RESULT eventid="1065" points="188" swimtime="00:00:40.02" resultid="1968" heatid="2079" lane="4" />
                <RESULT eventid="1099" points="153" swimtime="00:00:47.13" resultid="1969" heatid="2134" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Viechineski Bernardes" birthdate="2011-02-26" gender="M" nation="BRA" license="390879" swrid="5602588" athleteid="1955" externalid="390879">
              <RESULTS>
                <RESULT eventid="1067" points="150" swimtime="00:01:30.88" resultid="1956" heatid="2084" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="185" swimtime="00:01:18.65" resultid="1957" heatid="2120" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="147" swimtime="00:01:44.65" resultid="1958" heatid="2148" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="PGRO-SAGRADA FAMIL,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1091" points="237" swimtime="00:02:12.11" resultid="1980" heatid="2128" lane="5" entrytime="00:02:23.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                    <SPLIT distance="100" swimtime="00:01:08.93" />
                    <SPLIT distance="150" swimtime="00:01:43.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1947" number="1" />
                    <RELAYPOSITION athleteid="1974" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1955" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1959" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1109" points="182" swimtime="00:02:38.25" resultid="1981" heatid="2152" lane="5" entrytime="00:02:31.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.23" />
                    <SPLIT distance="100" swimtime="00:01:24.50" />
                    <SPLIT distance="150" swimtime="00:02:03.81" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1974" number="1" />
                    <RELAYPOSITION athleteid="1959" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1947" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1955" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="PGRO-SAGRADA FAMIL,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1093" points="238" swimtime="00:02:29.09" resultid="1978" heatid="2129" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:14.09" />
                    <SPLIT distance="150" swimtime="00:01:54.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1970" number="1" />
                    <RELAYPOSITION athleteid="1951" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1967" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1963" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1107" points="204" swimtime="00:02:53.80" resultid="1979" heatid="2151" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.71" />
                    <SPLIT distance="100" swimtime="00:01:28.90" />
                    <SPLIT distance="150" swimtime="00:02:13.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1951" number="1" />
                    <RELAYPOSITION athleteid="1963" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1970" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1967" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="PGRO-SAGRADA FAMIL,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1077" points="225" swimtime="00:02:36.33" resultid="1982" heatid="2100" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.01" />
                    <SPLIT distance="100" swimtime="00:01:28.05" />
                    <SPLIT distance="150" swimtime="00:02:07.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1951" number="1" />
                    <RELAYPOSITION athleteid="1963" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1947" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1959" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="15580" nation="BRA" region="PR" clubid="1469" name="Colégio Nossa Senhora Do Rosário, Curitiba" shortname="Ctba-N.Srª.Rosário,C">
          <ATHLETES>
            <ATHLETE firstname="Daniel" lastname="Cravcenco Marcondes" birthdate="2011-05-06" gender="M" nation="BRA" license="406867" swrid="5723023" athleteid="1474" externalid="406867">
              <RESULTS>
                <RESULT eventid="1071" points="217" swimtime="00:00:36.16" resultid="1475" heatid="2091" lane="5" />
                <RESULT eventid="1063" points="263" swimtime="00:00:31.46" resultid="1476" heatid="2070" lane="8" />
                <RESULT eventid="1087" status="DSQ" swimtime="00:01:13.77" resultid="1477" heatid="2120" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Cravcenco Marcondes" birthdate="2012-06-23" gender="F" nation="BRA" license="406866" swrid="5725987" athleteid="1470" externalid="406866">
              <RESULTS>
                <RESULT eventid="1085" points="175" swimtime="00:01:29.74" resultid="1471" heatid="2114" lane="5" entrytime="00:01:23.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="166" swimtime="00:00:51.53" resultid="1472" heatid="2105" lane="4" entrytime="00:00:48.19" entrycourse="SCM" />
                <RESULT eventid="1099" points="155" swimtime="00:00:46.93" resultid="1473" heatid="2137" lane="2" entrytime="00:00:44.16" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13953" nation="BRA" region="PR" clubid="1606" name="Escola Saber, Cascavel" shortname="Cvel-Saber,E">
          <ATHLETES>
            <ATHLETE firstname="Guilherme" lastname="Cordeiro Silva" birthdate="2011-09-04" gender="M" nation="BRA" license="380664" swrid="5596877" athleteid="1607" externalid="380664">
              <RESULTS>
                <RESULT eventid="1075" status="SICK" swimtime="00:00:00.00" resultid="1608" entrytime="00:02:57.90" entrycourse="SCM" />
                <RESULT eventid="1083" status="SICK" swimtime="00:00:00.00" resultid="1609" entrytime="00:00:40.73" entrycourse="SCM" />
                <RESULT eventid="1105" status="SICK" swimtime="00:00:00.00" resultid="1610" entrytime="00:01:29.78" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17684" nation="BRA" region="PR" clubid="1369" name="Colégio Estadual Gelvira Correa Pacheco, Curitiba" shortname="Ctba-Gelvira Corre,C">
          <ATHLETES>
            <ATHLETE firstname="Leonardo" lastname="Fernandes" birthdate="2010-03-13" gender="M" nation="BRA" license="339266" swrid="5588695" athleteid="1370" externalid="339266">
              <RESULTS>
                <RESULT eventid="1067" points="299" swimtime="00:01:12.22" resultid="1371" heatid="2086" lane="3" entrytime="00:01:06.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="409" swimtime="00:00:27.15" resultid="1372" heatid="2076" lane="4" entrytime="00:00:26.41" entrycourse="SCM" />
                <RESULT eventid="1087" status="RJC" swimtime="00:00:00.00" resultid="1373" entrytime="00:00:58.19" entrycourse="SCM" />
                <RESULT eventid="1101" points="386" swimtime="00:00:30.36" resultid="1374" heatid="2141" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16304" nation="BRA" region="PR" clubid="1173" name="Escola Estadual Aline Picheth, Curitiba" shortname="Ctba-Alinepicheth,Ee">
          <ATHLETES>
            <ATHLETE firstname="Eduarda" lastname="Azevedo Birsneek" birthdate="2010-03-31" gender="F" nation="BRA" license="391145" swrid="5389427" athleteid="1174" externalid="391145">
              <RESULTS>
                <RESULT eventid="1061" points="183" swimtime="00:06:47.12" resultid="1175" heatid="2067" lane="5" entrytime="00:07:02.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.06" />
                    <SPLIT distance="100" swimtime="00:01:31.82" />
                    <SPLIT distance="150" swimtime="00:02:23.61" />
                    <SPLIT distance="200" swimtime="00:03:14.35" />
                    <SPLIT distance="250" swimtime="00:04:06.17" />
                    <SPLIT distance="300" swimtime="00:04:59.52" />
                    <SPLIT distance="350" swimtime="00:05:53.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1089" status="DSQ" swimtime="00:03:42.89" resultid="1176" heatid="2126" lane="8" entrytime="00:03:53.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.53" />
                    <SPLIT distance="100" swimtime="00:01:39.94" />
                    <SPLIT distance="150" swimtime="00:02:53.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="128" swimtime="00:01:47.06" resultid="1177" heatid="2130" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18834" nation="BRA" region="PR" clubid="2020" name="Colégio Estadual João Arnaldo Ritt, Toledo" shortname="Tole-João Ritt,Ce">
          <ATHLETES>
            <ATHLETE firstname="Yasmin" lastname="Pauly Follmann" birthdate="2011-04-19" gender="F" nation="BRA" license="V413886" athleteid="2021" externalid="V413886">
              <RESULTS>
                <RESULT eventid="1065" points="146" swimtime="00:00:43.45" resultid="2022" heatid="2077" lane="5" />
                <RESULT eventid="1081" status="DSQ" swimtime="00:00:50.65" resultid="2023" heatid="2105" lane="8" />
                <RESULT eventid="1099" points="176" swimtime="00:00:45.04" resultid="2024" heatid="2135" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="14773" nation="BRA" region="PR" clubid="1364" name="Escola Estadual Profº Elias Abrahão, Curitiba" shortname="Ctba-E.Abrahão,Ee">
          <ATHLETES>
            <ATHLETE firstname="Kaylane" lastname="Marques Ferreira" birthdate="2010-03-06" gender="F" nation="BRA" license="391146" swrid="5600211" athleteid="1365" externalid="391146">
              <RESULTS>
                <RESULT eventid="1073" points="317" swimtime="00:00:35.73" resultid="1366" heatid="2095" lane="5" entrytime="00:00:39.07" entrycourse="SCM" />
                <RESULT eventid="1065" points="289" swimtime="00:00:34.66" resultid="1367" heatid="2081" lane="2" entrytime="00:00:36.87" entrycourse="SCM" />
                <RESULT eventid="1095" points="217" swimtime="00:01:29.83" resultid="1368" heatid="2130" lane="3" entrytime="00:01:38.41" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6517" nation="BRA" region="PR" clubid="1900" name="Colégio Regina Mundi, Maringá" shortname="Mrga-Regina Mundi,C">
          <ATHLETES>
            <ATHLETE firstname="Felipe" lastname="Lima Coelho" birthdate="2012-12-12" gender="M" nation="BRA" license="393775" swrid="5615959" athleteid="1901" externalid="393775">
              <RESULTS>
                <RESULT eventid="1067" status="DNS" swimtime="00:00:00.00" resultid="1902" heatid="2084" lane="3" />
                <RESULT eventid="1087" status="DNS" swimtime="00:00:00.00" resultid="1903" heatid="2122" lane="1" entrytime="00:01:26.02" entrycourse="SCM" />
                <RESULT eventid="1101" status="DNS" swimtime="00:00:00.00" resultid="1904" heatid="2142" lane="1" entrytime="00:00:42.35" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6500" nation="BRA" region="PR" clubid="1500" name="Colégio Sagrado Coração De Jesus, Curitiba" shortname="Ctba-Sag.Cor.Jesus,C">
          <ATHLETES>
            <ATHLETE firstname="Miguel" lastname="Fernandes  Dos Reis" birthdate="2012-09-18" gender="M" nation="BRA" license="369279" swrid="5588696" athleteid="1510" externalid="369279">
              <RESULTS>
                <RESULT eventid="1063" points="236" swimtime="00:00:32.58" resultid="1511" heatid="2074" lane="3" entrytime="00:00:32.13" entrycourse="SCM" />
                <RESULT eventid="1087" points="251" swimtime="00:01:11.00" resultid="1512" heatid="2123" lane="3" entrytime="00:01:09.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="224" swimtime="00:01:18.60" resultid="1513" heatid="2132" lane="4" entrytime="00:01:18.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Ribeiro Melo" birthdate="2011-07-01" gender="F" nation="BRA" license="390923" swrid="5602577" athleteid="1514" externalid="390923">
              <RESULTS>
                <RESULT eventid="1069" status="RJC" swimtime="00:00:00.00" resultid="1515" />
                <RESULT eventid="1065" points="420" swimtime="00:00:30.60" resultid="1516" heatid="2082" lane="3" entrytime="00:00:31.95" entrycourse="SCM" />
                <RESULT eventid="1085" points="379" swimtime="00:01:09.38" resultid="1517" heatid="2116" lane="2" entrytime="00:01:12.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="250" swimtime="00:01:38.95" resultid="1518" heatid="2146" lane="1" entrytime="00:01:35.91" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Magalhaes Dos Reis" birthdate="2010-05-05" gender="M" nation="BRA" license="356361" swrid="5600207" athleteid="1501" externalid="356361">
              <RESULTS>
                <RESULT eventid="1063" points="378" swimtime="00:00:27.86" resultid="1502" heatid="2076" lane="2" entrytime="00:00:27.78" entrycourse="SCM" />
                <RESULT eventid="1087" points="408" swimtime="00:01:00.44" resultid="1503" heatid="2124" lane="6" entrytime="00:01:02.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="295" swimtime="00:01:22.97" resultid="1504" heatid="2150" lane="5" entrytime="00:01:19.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Leao" birthdate="2011-09-18" gender="M" nation="BRA" license="366880" swrid="5602553" athleteid="1505" externalid="366880">
              <RESULTS>
                <RESULT eventid="1075" points="292" swimtime="00:02:45.13" resultid="1506" heatid="2098" lane="4" entrytime="00:02:54.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.91" />
                    <SPLIT distance="100" swimtime="00:01:19.07" />
                    <SPLIT distance="150" swimtime="00:02:09.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="316" swimtime="00:00:29.57" resultid="1507" heatid="2075" lane="2" entrytime="00:00:30.71" entrycourse="SCM" />
                <RESULT eventid="1079" points="360" swimtime="00:04:58.27" resultid="1508" heatid="2103" lane="7" entrytime="00:05:02.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                    <SPLIT distance="100" swimtime="00:01:10.22" />
                    <SPLIT distance="150" swimtime="00:01:47.74" />
                    <SPLIT distance="200" swimtime="00:02:25.61" />
                    <SPLIT distance="250" swimtime="00:03:03.89" />
                    <SPLIT distance="300" swimtime="00:03:42.61" />
                    <SPLIT distance="350" swimtime="00:04:21.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" status="RJC" swimtime="00:00:00.00" resultid="1509" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4194" nation="BRA" region="PR" clubid="1154" name="Colégio Estadual Unidade Polo, Campo Mourão" shortname="Cmou-Un.Polo,Ce">
          <ATHLETES>
            <ATHLETE firstname="Gabriel" lastname="Giroldo Santos" birthdate="2011-05-16" gender="M" nation="BRA" license="V399602" athleteid="1155" externalid="V399602">
              <RESULTS>
                <RESULT eventid="1075" status="DSQ" swimtime="00:03:29.52" resultid="1156" heatid="2097" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.60" />
                    <SPLIT distance="100" swimtime="00:01:41.05" />
                    <SPLIT distance="150" swimtime="00:02:40.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="186" swimtime="00:00:35.31" resultid="1157" heatid="2073" lane="1" entrytime="00:00:44.25" entrycourse="SCM" />
                <RESULT eventid="1101" points="128" swimtime="00:00:43.79" resultid="1158" heatid="2140" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18826" nation="BRA" region="PR" clubid="1395" name="Escola Municipal Júlia Amaral DI Lenna" shortname="Ctba-Júlia.Lenna,Em">
          <ATHLETES>
            <ATHLETE firstname="Davi" lastname="Da Reginalda" birthdate="2012-11-09" gender="M" nation="BRA" license="400275" swrid="5717253" athleteid="1400" externalid="400275">
              <RESULTS>
                <RESULT eventid="1063" points="231" swimtime="00:00:32.85" resultid="1401" heatid="2074" lane="6" entrytime="00:00:32.43" entrycourse="SCM" />
                <RESULT eventid="1083" points="165" swimtime="00:00:45.45" resultid="1402" heatid="2108" lane="3" />
                <RESULT eventid="1101" points="189" swimtime="00:00:38.50" resultid="1403" heatid="2143" lane="8" entrytime="00:00:37.59" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="De Reginalda" birthdate="2011-07-22" gender="M" nation="BRA" license="400323" swrid="5717257" athleteid="1396" externalid="400323">
              <RESULTS>
                <RESULT eventid="1067" points="330" swimtime="00:01:09.87" resultid="1397" heatid="2085" lane="4" entrytime="00:01:13.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="389" swimtime="00:00:27.61" resultid="1398" heatid="2073" lane="6" entrytime="00:00:39.22" entrycourse="SCM" />
                <RESULT eventid="1101" points="344" swimtime="00:00:31.54" resultid="1399" heatid="2143" lane="5" entrytime="00:00:33.48" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17659" nation="BRA" region="PR" clubid="1380" name="Escola Internacional De Curitiba" shortname="Ctba-Inernacional,E">
          <ATHLETES>
            <ATHLETE firstname="Sophie" lastname="Kraemer Geremia" birthdate="2011-07-20" gender="F" nation="BRA" license="366908" swrid="5588763" athleteid="1381" externalid="366908">
              <RESULTS>
                <RESULT eventid="1069" points="438" swimtime="00:01:12.23" resultid="1382" heatid="2090" lane="6" entrytime="00:01:15.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="434" swimtime="00:01:06.35" resultid="1383" heatid="2117" lane="1" entrytime="00:01:06.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="388" swimtime="00:00:34.61" resultid="1384" heatid="2138" lane="2" entrytime="00:00:36.99" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ian" lastname="Thierbach Ruiz" birthdate="2011-10-12" gender="M" nation="BRA" license="V413946" athleteid="1385" externalid="V413946">
              <RESULTS>
                <RESULT eventid="1063" points="224" swimtime="00:00:33.19" resultid="1386" heatid="2072" lane="1" />
                <RESULT eventid="1087" points="190" swimtime="00:01:17.92" resultid="1387" heatid="2119" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="170" swimtime="00:00:44.96" resultid="1388" heatid="2109" lane="8" />
                <RESULT eventid="1105" status="RJC" swimtime="00:00:00.00" resultid="1389" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="14010" nation="BRA" region="PR" clubid="1557" name="Colégio Expressão, Cascavel" shortname="Cvel-Expressão,C">
          <ATHLETES>
            <ATHLETE firstname="Danilo" lastname="Rodrigues" birthdate="2011-05-23" gender="M" nation="BRA" license="370763" swrid="5596934" athleteid="1562" externalid="370763">
              <RESULTS>
                <RESULT eventid="1071" points="270" swimtime="00:00:33.63" resultid="1563" heatid="2093" lane="7" entrytime="00:00:34.02" entrycourse="SCM" />
                <RESULT eventid="1087" points="292" swimtime="00:01:07.58" resultid="1564" heatid="2119" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="266" swimtime="00:01:14.23" resultid="1565" heatid="2133" lane="7" entrytime="00:01:15.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ramirez Vasconcelos" birthdate="2011-04-06" gender="M" nation="BRA" license="392013" swrid="4863662" athleteid="1566" externalid="392013">
              <RESULTS>
                <RESULT eventid="1075" status="DSQ" swimtime="00:02:41.19" resultid="1567" heatid="2099" lane="1" entrytime="00:02:53.12" entrycourse="SCM" />
                <RESULT eventid="1083" points="263" swimtime="00:00:38.91" resultid="1568" heatid="2109" lane="1" />
                <RESULT eventid="1105" points="308" swimtime="00:01:21.79" resultid="1569" heatid="2150" lane="8" entrytime="00:01:28.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Claudio" lastname="Rohnelt" birthdate="2010-03-08" gender="M" nation="BRA" license="357954" swrid="5596935" athleteid="1558" externalid="357954">
              <RESULTS>
                <RESULT eventid="1071" points="270" swimtime="00:00:33.63" resultid="1559" heatid="2093" lane="8" entrytime="00:00:35.78" entrycourse="SCM" />
                <RESULT eventid="1079" points="356" swimtime="00:04:59.39" resultid="1560" heatid="2103" lane="1" entrytime="00:05:06.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                    <SPLIT distance="100" swimtime="00:01:10.92" />
                    <SPLIT distance="150" swimtime="00:01:49.13" />
                    <SPLIT distance="200" swimtime="00:02:27.29" />
                    <SPLIT distance="250" swimtime="00:03:05.14" />
                    <SPLIT distance="300" swimtime="00:03:43.63" />
                    <SPLIT distance="350" swimtime="00:04:21.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="280" swimtime="00:01:13.00" resultid="1561" heatid="2133" lane="1" entrytime="00:01:15.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13979" nation="BRA" region="PR" clubid="1127" name="Colégio Conexão, Campo Mourão" shortname="Cmou-Conexão,C">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Gabrieli Oliveira" birthdate="2010-09-23" gender="F" nation="BRA" license="403428" swrid="5676288" athleteid="1128" externalid="403428">
              <RESULTS>
                <RESULT eventid="1069" points="193" swimtime="00:01:34.91" resultid="1129" heatid="2088" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="271" swimtime="00:00:35.41" resultid="1130" heatid="2078" lane="6" />
                <RESULT eventid="1099" points="182" swimtime="00:00:44.54" resultid="1131" heatid="2136" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15636" nation="BRA" region="PR" clubid="1588" name="CCM Professora Júlia Wanderley, Cascavel" shortname="Cvel-J.Wanderley,CCM">
          <ATHLETES>
            <ATHLETE firstname="Guilherme" lastname="Zimmermann" birthdate="2010-01-19" gender="M" nation="BRA" license="357160" swrid="5588977" athleteid="1589" externalid="357160">
              <RESULTS>
                <RESULT eventid="1067" points="417" swimtime="00:01:04.69" resultid="1590" heatid="2086" lane="5" entrytime="00:01:05.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="476" swimtime="00:02:20.32" resultid="1591" heatid="2099" lane="4" entrytime="00:02:20.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:08.80" />
                    <SPLIT distance="150" swimtime="00:01:49.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="538" swimtime="00:04:20.92" resultid="1592" heatid="2103" lane="5" entrytime="00:04:21.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                    <SPLIT distance="100" swimtime="00:01:03.77" />
                    <SPLIT distance="150" swimtime="00:01:37.15" />
                    <SPLIT distance="200" swimtime="00:02:10.74" />
                    <SPLIT distance="250" swimtime="00:02:44.15" />
                    <SPLIT distance="300" swimtime="00:03:17.80" />
                    <SPLIT distance="350" swimtime="00:03:50.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hendrik" lastname="Alteiro Groenwold" birthdate="2011-03-23" gender="M" nation="BRA" license="365756" swrid="5588520" athleteid="1593" externalid="365756">
              <RESULTS>
                <RESULT eventid="1071" points="358" swimtime="00:00:30.61" resultid="1594" heatid="2091" lane="7" />
                <RESULT eventid="1079" points="421" swimtime="00:04:43.13" resultid="1595" heatid="2103" lane="6" entrytime="00:04:44.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:04.98" />
                    <SPLIT distance="150" swimtime="00:01:40.03" />
                    <SPLIT distance="200" swimtime="00:02:16.50" />
                    <SPLIT distance="250" swimtime="00:02:53.57" />
                    <SPLIT distance="300" swimtime="00:03:30.17" />
                    <SPLIT distance="350" swimtime="00:04:07.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="395" swimtime="00:01:05.08" resultid="1596" heatid="2133" lane="3" entrytime="00:01:10.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Macedo Medeiros" birthdate="2012-05-12" gender="M" nation="BRA" license="392015" swrid="4697574" athleteid="1597" externalid="392015">
              <RESULTS>
                <RESULT eventid="1075" points="167" swimtime="00:03:18.99" resultid="1598" heatid="2097" lane="5" entrytime="00:03:46.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.93" />
                    <SPLIT distance="100" swimtime="00:01:43.84" />
                    <SPLIT distance="150" swimtime="00:02:36.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="163" swimtime="00:00:45.66" resultid="1599" heatid="2110" lane="1" entrytime="00:00:48.99" entrycourse="SCM" />
                <RESULT eventid="1097" points="107" swimtime="00:01:40.52" resultid="1600" heatid="2132" lane="2" entrytime="00:01:48.79" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15564" nation="BRA" region="PR" clubid="1939" name="Colégio Alfa Rede De Ensino, Ponta Grossa" shortname="Pgro-Alfa Ensino,C">
          <ATHLETES>
            <ATHLETE firstname="Guilherme" lastname="Novassat Paula" birthdate="2010-03-29" gender="M" nation="BRA" license="V413872" athleteid="1940" externalid="V413872">
              <RESULTS>
                <RESULT eventid="1071" points="196" swimtime="00:00:37.43" resultid="1941" heatid="2092" lane="1" />
                <RESULT eventid="1063" points="215" swimtime="00:00:33.62" resultid="1942" heatid="2069" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15570" nation="BRA" region="PR" clubid="1280" name="Colégio Bom Jesus Seminário, Curitiba" shortname="Ctba-Bj Seminário,C">
          <ATHLETES>
            <ATHLETE firstname="Nina" lastname="Rocha Ribeiro Da Silva" birthdate="2010-09-22" gender="F" nation="BRA" license="367216" swrid="5588884" athleteid="1281" externalid="367216">
              <RESULTS>
                <RESULT eventid="1081" points="463" swimtime="00:00:36.67" resultid="1282" heatid="2105" lane="7" />
                <RESULT eventid="1103" points="432" swimtime="00:01:22.43" resultid="1283" heatid="2147" lane="4" entrytime="00:01:20.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2617" nation="BRA" region="PR" clubid="2025" name="Colégio La Salle, Toledo" shortname="Tole-La Salle,C">
          <ATHLETES>
            <ATHLETE firstname="Isabela" lastname="Torres Romancini" birthdate="2010-05-28" gender="F" nation="BRA" license="347218" swrid="5622309" athleteid="2026" externalid="347218">
              <RESULTS>
                <RESULT eventid="1069" points="414" swimtime="00:01:13.60" resultid="2027" heatid="2090" lane="1" entrytime="00:01:17.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1073" points="380" swimtime="00:00:33.64" resultid="2028" heatid="2096" lane="8" entrytime="00:00:37.00" entrycourse="SCM" />
                <RESULT eventid="1099" points="421" swimtime="00:00:33.68" resultid="2029" heatid="2138" lane="7" entrytime="00:00:37.54" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lavinia" lastname="Martins Paludo" birthdate="2010-09-30" gender="F" nation="BRA" license="347217" swrid="5652624" athleteid="2030" externalid="347217">
              <RESULTS>
                <RESULT eventid="1089" status="DSQ" swimtime="00:03:24.05" resultid="2031" heatid="2125" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.71" />
                    <SPLIT distance="100" swimtime="00:01:43.21" />
                    <SPLIT distance="150" swimtime="00:02:38.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="221" swimtime="00:00:46.87" resultid="2032" heatid="2106" lane="2" entrytime="00:00:44.97" entrycourse="SCM" />
                <RESULT eventid="1103" points="217" swimtime="00:01:43.76" resultid="2033" heatid="2145" lane="5" entrytime="00:01:38.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2647" nation="BRA" region="PR" clubid="1983" name="Colégio Sepam, Ponta Grossa" shortname="Pgro-Sepam,C">
          <ATHLETES>
            <ATHLETE firstname="Luiz" lastname="Miguel Rodrigues Neto" birthdate="2010-05-12" gender="M" nation="BRA" license="V399583" athleteid="1984" externalid="V399583">
              <RESULTS>
                <RESULT eventid="1083" points="210" swimtime="00:00:41.94" resultid="1985" heatid="2110" lane="6" entrytime="00:00:45.44" entrycourse="SCM" />
                <RESULT eventid="1105" status="DSQ" swimtime="00:01:40.33" resultid="1986" heatid="2148" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="205" reactiontime="+750" swimtime="00:00:37.47" resultid="1987" heatid="2142" lane="8" entrytime="00:00:43.60" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Clara Domingues" birthdate="2012-01-19" gender="F" nation="BRA" license="377291" swrid="5588599" athleteid="1988" externalid="377291">
              <RESULTS>
                <RESULT eventid="1069" points="170" swimtime="00:01:38.95" resultid="1989" heatid="2088" lane="5" entrytime="00:01:36.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1061" points="234" swimtime="00:06:14.83" resultid="1990" heatid="2067" lane="4" entrytime="00:06:19.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:26.49" />
                    <SPLIT distance="150" swimtime="00:02:13.87" />
                    <SPLIT distance="200" swimtime="00:03:03.60" />
                    <SPLIT distance="250" swimtime="00:03:52.95" />
                    <SPLIT distance="300" swimtime="00:04:41.89" />
                    <SPLIT distance="350" swimtime="00:05:30.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="262" swimtime="00:01:18.44" resultid="1991" heatid="2115" lane="7" entrytime="00:01:19.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16332" nation="BRA" region="PR" clubid="1771" name="Colégio Alfa Tesla, Maringá" shortname="Mrga-Alfa Tesla,C">
          <ATHLETES>
            <ATHLETE firstname="Bianca" lastname="Corsine Ferreira" birthdate="2010-03-10" gender="F" nation="BRA" license="353591" swrid="5588608" athleteid="1772" externalid="353591">
              <RESULTS>
                <RESULT eventid="1069" points="398" swimtime="00:01:14.62" resultid="1773" heatid="2090" lane="4" entrytime="00:01:13.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="353" swimtime="00:00:40.13" resultid="1774" heatid="2106" lane="5" entrytime="00:00:42.04" entrycourse="SCM" />
                <RESULT eventid="1099" points="407" swimtime="00:00:34.06" resultid="1775" heatid="2138" lane="4" entrytime="00:00:34.15" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eloah" lastname="Juvedi Trindade" birthdate="2011-03-05" gender="F" nation="BRA" license="396829" swrid="5641768" athleteid="1776" externalid="396829">
              <RESULTS>
                <RESULT eventid="1073" status="DNS" swimtime="00:00:00.00" resultid="1777" heatid="2094" lane="3" />
                <RESULT eventid="1065" status="DNS" swimtime="00:00:00.00" resultid="1778" heatid="2081" lane="7" entrytime="00:00:36.87" entrycourse="SCM" />
                <RESULT eventid="1103" points="249" swimtime="00:01:39.10" resultid="1779" heatid="2146" lane="8" entrytime="00:01:36.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17666" nation="BRA" region="PR" clubid="1721" name="Colégio Integrado Sônia Marcondes, Ibiporã" shortname="Ibip-Sonia Marcon.,C">
          <ATHLETES>
            <ATHLETE firstname="Gabriela" lastname="Gomes" birthdate="2011-12-03" gender="F" nation="BRA" license="382051" swrid="5603846" athleteid="1722" externalid="382051">
              <RESULTS>
                <RESULT eventid="1069" points="204" swimtime="00:01:33.12" resultid="1723" heatid="2088" lane="3" entrytime="00:01:38.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="227" swimtime="00:01:22.27" resultid="1724" heatid="2114" lane="4" entrytime="00:01:22.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="198" swimtime="00:00:43.29" resultid="1725" heatid="2137" lane="7" entrytime="00:00:45.25" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6498" nation="BRA" region="PR" clubid="1905" name="Colégio Santa Cruz, Maringá" shortname="Mrga-Santa Cruz,C">
          <ATHLETES>
            <ATHLETE firstname="Gabriel" lastname="Schuch Pimpao" birthdate="2010-05-17" gender="M" nation="BRA" license="355586" swrid="5588908" athleteid="1906" externalid="355586">
              <RESULTS>
                <RESULT eventid="1067" points="351" swimtime="00:01:08.45" resultid="1907" heatid="2086" lane="2" entrytime="00:01:10.45" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="354" swimtime="00:02:34.86" resultid="1908" heatid="2099" lane="7" entrytime="00:02:35.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:13.03" />
                    <SPLIT distance="150" swimtime="00:01:57.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="315" swimtime="00:00:32.47" resultid="1909" heatid="2143" lane="7" entrytime="00:00:34.31" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monique" lastname="Istake" birthdate="2012-04-03" gender="F" nation="BRA" license="372023" swrid="5603857" athleteid="1910" externalid="372023">
              <RESULTS>
                <RESULT eventid="1073" points="335" swimtime="00:00:35.09" resultid="1911" heatid="2096" lane="2" entrytime="00:00:36.43" entrycourse="SCM" />
                <RESULT eventid="1089" points="272" swimtime="00:03:07.98" resultid="1912" heatid="2126" lane="6" entrytime="00:03:08.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.86" />
                    <SPLIT distance="100" swimtime="00:01:27.15" />
                    <SPLIT distance="150" swimtime="00:02:24.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="250" swimtime="00:01:25.70" resultid="1913" heatid="2131" lane="2" entrytime="00:01:25.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18830" nation="BRA" region="PR" clubid="1709" name="Colégio Estadual Prof. Jaime Rodrigues, Guaíra" shortname="Guai-Jaime Rodri.,Ce">
          <ATHLETES>
            <ATHLETE firstname="Ana" lastname="Julia Andreolla" birthdate="2011-12-19" gender="F" nation="BRA" license="V413887" athleteid="1710" externalid="V413887">
              <RESULTS>
                <RESULT eventid="1065" points="175" swimtime="00:00:40.96" resultid="1711" heatid="2077" lane="3" />
                <RESULT eventid="1085" points="145" swimtime="00:01:35.56" resultid="1712" heatid="2113" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="100" swimtime="00:00:54.27" resultid="1713" heatid="2135" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="889" nation="BRA" region="PR" clubid="1284" name="Colégio Estadual Do Paraná, Curitiba" shortname="Ctba-Cep,Ce">
          <ATHLETES>
            <ATHLETE firstname="Geovana" lastname="Dos Santos" birthdate="2011-01-20" gender="F" nation="BRA" license="367254" swrid="5602533" athleteid="1285" externalid="367254">
              <RESULTS>
                <RESULT eventid="1069" points="260" swimtime="00:01:25.90" resultid="1286" heatid="2088" lane="4" entrytime="00:01:33.77" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="310" swimtime="00:00:33.85" resultid="1287" heatid="2082" lane="1" entrytime="00:00:34.14" entrycourse="SCM" />
                <RESULT eventid="1085" points="288" swimtime="00:01:16.02" resultid="1288" heatid="2115" lane="2" entrytime="00:01:16.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Galdino Silva" birthdate="2012-06-08" gender="F" nation="BRA" license="V413861" athleteid="1289" externalid="V413861">
              <RESULTS>
                <RESULT eventid="1065" points="135" swimtime="00:00:44.64" resultid="1290" heatid="2079" lane="3" />
                <RESULT eventid="1085" points="130" swimtime="00:01:39.12" resultid="1291" heatid="2112" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="105" swimtime="00:00:53.46" resultid="1292" heatid="2135" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Oliveira Dprospero" birthdate="2012-12-06" gender="F" nation="BRA" license="V413862" athleteid="1293" externalid="V413862">
              <RESULTS>
                <RESULT eventid="1065" points="136" swimtime="00:00:44.51" resultid="1294" heatid="2079" lane="2" />
                <RESULT eventid="1085" points="108" swimtime="00:01:45.43" resultid="1295" heatid="2114" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" status="DSQ" swimtime="00:01:05.65" resultid="1296" heatid="2104" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Sufredini Machado" birthdate="2012-09-21" gender="M" nation="BRA" license="V413934" athleteid="1297" externalid="V413934">
              <RESULTS>
                <RESULT eventid="1063" points="103" swimtime="00:00:42.94" resultid="1298" heatid="2070" lane="5" />
                <RESULT eventid="1087" points="92" swimtime="00:01:39.07" resultid="1299" heatid="2120" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="90" swimtime="00:07:52.60" resultid="1300" heatid="2102" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.60" />
                    <SPLIT distance="100" swimtime="00:01:39.00" />
                    <SPLIT distance="150" swimtime="00:02:40.62" />
                    <SPLIT distance="200" swimtime="00:03:42.40" />
                    <SPLIT distance="250" swimtime="00:04:46.23" />
                    <SPLIT distance="300" swimtime="00:05:45.56" />
                    <SPLIT distance="350" swimtime="00:06:50.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cesar" lastname="Danilo Da Silva Andruzinski" birthdate="2011-03-27" gender="M" nation="BRA" license="V413935" athleteid="1301" externalid="V413935">
              <RESULTS>
                <RESULT eventid="1071" status="WDR" swimtime="00:00:00.00" resultid="1302" />
                <RESULT eventid="1063" status="WDR" swimtime="00:00:00.00" resultid="1303" />
                <RESULT eventid="1087" status="WDR" swimtime="00:00:00.00" resultid="1304" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ehab" lastname="Moayad Abdallah" birthdate="2012-04-23" gender="M" nation="BRA" license="V413936" athleteid="1305" externalid="V413936">
              <RESULTS>
                <RESULT eventid="1063" points="143" swimtime="00:00:38.55" resultid="1306" heatid="2070" lane="2" />
                <RESULT eventid="1087" points="122" swimtime="00:01:30.26" resultid="1307" heatid="2121" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" status="DNS" swimtime="00:00:00.00" resultid="1308" heatid="2140" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Gabriel Schloegel Zacarias" birthdate="2012-09-05" gender="M" nation="BRA" license="V413937" athleteid="1309" externalid="V413937">
              <RESULTS>
                <RESULT eventid="1063" points="184" swimtime="00:00:35.42" resultid="1310" heatid="2069" lane="3" />
                <RESULT eventid="1087" points="163" swimtime="00:01:22.07" resultid="1311" heatid="2121" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="146" swimtime="00:06:42.39" resultid="1312" heatid="2102" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.88" />
                    <SPLIT distance="100" swimtime="00:01:33.63" />
                    <SPLIT distance="150" swimtime="00:02:24.43" />
                    <SPLIT distance="200" swimtime="00:03:16.57" />
                    <SPLIT distance="250" swimtime="00:04:09.32" />
                    <SPLIT distance="300" swimtime="00:05:01.53" />
                    <SPLIT distance="350" swimtime="00:05:51.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CTBA-CEP,CE &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1091" status="WDR" swimtime="00:00:00.00" resultid="1313" />
                <RESULT eventid="1109" status="WDR" swimtime="00:00:00.00" resultid="1314" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="CTBA-CEP,CE &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1077" points="105" swimtime="00:03:21.14" resultid="1315" heatid="2100" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.83" />
                    <SPLIT distance="100" swimtime="00:01:51.07" />
                    <SPLIT distance="150" swimtime="00:02:42.85" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1285" number="1" />
                    <RELAYPOSITION athleteid="1293" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1309" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1305" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="13506" nation="BRA" region="PR" clubid="1413" name="Colégio Marista Anjo Da Guarda, Curitiba" shortname="Ctba-Marista Anjo.,C">
          <ATHLETES>
            <ATHLETE firstname="Lorena" lastname="Mascarenhas" birthdate="2011-08-31" gender="F" nation="BRA" license="370581" swrid="5602558" athleteid="1414" externalid="370581">
              <RESULTS>
                <RESULT eventid="1069" points="372" swimtime="00:01:16.26" resultid="1415" heatid="2089" lane="5" entrytime="00:01:19.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="352" swimtime="00:00:40.17" resultid="1416" heatid="2104" lane="3" />
                <RESULT eventid="1099" points="345" swimtime="00:00:35.97" resultid="1417" heatid="2134" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Galvao" birthdate="2011-03-11" gender="M" nation="BRA" license="381989" swrid="5602541" athleteid="1418" externalid="381989">
              <RESULTS>
                <RESULT eventid="1063" status="DNS" swimtime="00:00:00.00" resultid="1419" heatid="2070" lane="7" entrytime="00:00:31.14" entrycourse="SCM" />
                <RESULT eventid="1087" status="DNS" swimtime="00:00:00.00" resultid="1420" heatid="2123" lane="6" entrytime="00:01:09.39" entrycourse="SCM" />
                <RESULT eventid="1101" status="DNS" swimtime="00:00:00.00" resultid="1421" heatid="2139" lane="4" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3725" nation="BRA" region="PR" clubid="1748" name="Colégio Sagrada Família, Mandaguari" shortname="Mdri-Sagrada Fami.,C">
          <ATHLETES>
            <ATHLETE firstname="Mariana" lastname="Vitoria Henriques" birthdate="2011-03-26" gender="F" nation="BRA" license="V413890" athleteid="1749" externalid="V413890">
              <RESULTS>
                <RESULT eventid="1065" points="57" swimtime="00:00:59.44" resultid="1750" heatid="2079" lane="7" />
                <RESULT eventid="1099" points="68" swimtime="00:01:01.71" resultid="1751" heatid="2135" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18816" nation="BRA" region="PR" clubid="1690" name="Colégio Bom Pastor Lancaster, Foz Do Iguaçu" shortname="Fozi-Lancaster,C">
          <ATHLETES>
            <ATHLETE firstname="Mayumi" lastname="Napole" birthdate="2010-02-01" gender="F" nation="BRA" license="376446" swrid="5596918" athleteid="1691" externalid="376446" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1065" points="398" swimtime="00:00:31.15" resultid="1692" heatid="2083" lane="7" entrytime="00:00:31.09" entrycourse="SCM" />
                <RESULT eventid="1085" points="366" swimtime="00:01:10.22" resultid="1693" heatid="2116" lane="4" entrytime="00:01:08.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="284" swimtime="00:01:34.82" resultid="1694" heatid="2147" lane="8" entrytime="00:01:28.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18853" nation="BRA" region="PR" clubid="1539" name="Escola Trilhas, Curitiba" shortname="Ctba-Trilhas,E">
          <ATHLETES>
            <ATHLETE firstname="Joaquim" lastname="Pellanda" birthdate="2010-11-12" gender="M" nation="BRA" license="356352" swrid="5600233" athleteid="1540" externalid="356352">
              <RESULTS>
                <RESULT eventid="1075" points="416" swimtime="00:02:26.79" resultid="1541" heatid="2099" lane="3" entrytime="00:02:28.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                    <SPLIT distance="100" swimtime="00:01:10.26" />
                    <SPLIT distance="150" swimtime="00:01:54.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="460" swimtime="00:00:58.07" resultid="1542" heatid="2119" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="541" swimtime="00:04:20.48" resultid="1543" heatid="2103" lane="4" entrytime="00:04:21.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                    <SPLIT distance="100" swimtime="00:01:03.39" />
                    <SPLIT distance="150" swimtime="00:01:37.10" />
                    <SPLIT distance="200" swimtime="00:02:10.75" />
                    <SPLIT distance="250" swimtime="00:02:43.98" />
                    <SPLIT distance="300" swimtime="00:03:17.17" />
                    <SPLIT distance="350" swimtime="00:03:50.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11552" nation="BRA" region="PR" clubid="1570" name="Colégio Fag, Cascavel" shortname="Cvel-Fag,C">
          <ATHLETES>
            <ATHLETE firstname="Bernardo" lastname="Dillenburg Benetti" birthdate="2011-03-10" gender="M" nation="BRA" license="368119" swrid="5588656" athleteid="1575" externalid="368119">
              <RESULTS>
                <RESULT eventid="1067" points="287" swimtime="00:01:13.20" resultid="1576" heatid="2086" lane="7" entrytime="00:01:10.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="258" swimtime="00:01:26.77" resultid="1577" heatid="2149" lane="4" entrytime="00:01:28.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="282" swimtime="00:00:33.68" resultid="1578" heatid="2143" lane="6" entrytime="00:00:34.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Vitoria Gugel" birthdate="2011-12-08" gender="F" nation="BRA" license="365490" swrid="5588960" athleteid="1583" externalid="365490">
              <RESULTS>
                <RESULT eventid="1073" points="286" swimtime="00:00:36.97" resultid="1584" heatid="2094" lane="4" />
                <RESULT eventid="1089" points="333" swimtime="00:02:55.70" resultid="1585" heatid="2127" lane="8" entrytime="00:02:55.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.05" />
                    <SPLIT distance="100" swimtime="00:01:24.56" />
                    <SPLIT distance="150" swimtime="00:02:14.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="263" swimtime="00:01:24.35" resultid="1586" heatid="2130" lane="4" entrytime="00:01:31.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Stein Duarte" birthdate="2010-10-03" gender="F" nation="BRA" license="351635" swrid="5588923" athleteid="1571" externalid="351635">
              <RESULTS>
                <RESULT eventid="1069" points="465" swimtime="00:01:10.84" resultid="1572" heatid="2090" lane="5" entrytime="00:01:14.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1089" points="459" swimtime="00:02:37.87" resultid="1573" heatid="2127" lane="3" entrytime="00:02:42.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.38" />
                    <SPLIT distance="100" swimtime="00:01:13.44" />
                    <SPLIT distance="150" swimtime="00:02:00.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="428" swimtime="00:00:33.48" resultid="1574" heatid="2135" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emanuel" lastname="Ranieri" birthdate="2011-01-24" gender="M" nation="BRA" license="390838" swrid="5596930" athleteid="1579" externalid="390838">
              <RESULTS>
                <RESULT eventid="1067" status="DNS" swimtime="00:00:00.00" resultid="1580" heatid="2085" lane="7" entrytime="00:01:17.41" entrycourse="SCM" />
                <RESULT eventid="1087" status="DSQ" swimtime="00:01:16.60" resultid="1581" heatid="2123" lane="4" entrytime="00:01:05.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="231" swimtime="00:00:36.02" resultid="1582" heatid="2142" lane="3" entrytime="00:00:39.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="CVEL-FAG,C &quot;A&apos;" number="1">
              <RESULTS>
                <RESULT eventid="1077" points="311" swimtime="00:02:20.43" resultid="1587" heatid="2100" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:13.74" />
                    <SPLIT distance="150" swimtime="00:01:50.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1571" number="1" />
                    <RELAYPOSITION athleteid="1575" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1583" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1579" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="12478" nation="BRA" region="PR" clubid="1886" name="Colégio Paraná, Maringá" shortname="Mrga-Paraná,C">
          <ATHLETES>
            <ATHLETE firstname="Sarah" lastname="Chaim" birthdate="2011-05-29" gender="F" nation="BRA" license="370662" swrid="5409721" athleteid="1887" externalid="370662">
              <RESULTS>
                <RESULT eventid="1069" points="217" swimtime="00:01:31.25" resultid="1888" heatid="2089" lane="8" entrytime="00:01:33.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="296" swimtime="00:01:15.32" resultid="1889" heatid="2115" lane="6" entrytime="00:01:15.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="227" swimtime="00:00:41.38" resultid="1890" heatid="2137" lane="3" entrytime="00:00:43.17" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="8201" nation="BRA" region="PR" clubid="1675" name="Colégio Cooperativa Educacional, Foz Do Iguaçu" shortname="Fozi-Cooperativa,C">
          <ATHLETES>
            <ATHLETE firstname="Luisa" lastname="Franco" birthdate="2010-06-09" gender="F" nation="BRA" license="383849" swrid="5596896" athleteid="1676" externalid="383849">
              <RESULTS>
                <RESULT eventid="1061" points="342" swimtime="00:05:30.63" resultid="1677" heatid="2068" lane="6" entrytime="00:05:23.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.74" />
                    <SPLIT distance="100" swimtime="00:01:16.14" />
                    <SPLIT distance="150" swimtime="00:01:57.93" />
                    <SPLIT distance="200" swimtime="00:02:40.38" />
                    <SPLIT distance="250" swimtime="00:03:22.97" />
                    <SPLIT distance="300" swimtime="00:04:06.07" />
                    <SPLIT distance="350" swimtime="00:04:49.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1073" points="285" swimtime="00:00:37.01" resultid="1678" heatid="2096" lane="1" entrytime="00:00:36.82" entrycourse="SCM" />
                <RESULT eventid="1085" points="351" swimtime="00:01:11.21" resultid="1679" heatid="2116" lane="7" entrytime="00:01:12.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11559" nation="BRA" region="PR" clubid="1836" name="Escola Magnus Domini, Maringá" shortname="Mrga-Magnus Domin,E">
          <ATHLETES>
            <ATHLETE firstname="Enzo" lastname="Marques Picolo Vinha" birthdate="2010-07-01" gender="M" nation="BRA" license="366990" swrid="5603869" athleteid="1837" externalid="366990">
              <RESULTS>
                <RESULT eventid="1063" points="338" swimtime="00:00:28.94" resultid="1838" heatid="2076" lane="1" entrytime="00:00:29.23" entrycourse="SCM" />
                <RESULT eventid="1079" points="330" swimtime="00:05:07.02" resultid="1839" heatid="2101" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:09.73" />
                    <SPLIT distance="150" swimtime="00:01:47.80" />
                    <SPLIT distance="200" swimtime="00:02:27.74" />
                    <SPLIT distance="250" swimtime="00:03:08.11" />
                    <SPLIT distance="300" swimtime="00:03:48.77" />
                    <SPLIT distance="350" swimtime="00:04:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="262" swimtime="00:00:34.54" resultid="1840" heatid="2141" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Tonet Arruda Botelho" birthdate="2010-04-16" gender="M" nation="BRA" license="V413928" athleteid="1841" externalid="V413928">
              <RESULTS>
                <RESULT eventid="1063" points="239" swimtime="00:00:32.47" resultid="1842" heatid="2071" lane="7" />
                <RESULT eventid="1087" points="216" swimtime="00:01:14.66" resultid="1843" heatid="2118" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="188" swimtime="00:00:38.57" resultid="1844" heatid="2141" lane="8" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4210" nation="BRA" region="PR" clubid="2034" name="Colégio Estadual Francisco Galdin De Lima, Toledo" shortname="Tole-Ver. Franci.,Ce">
          <ATHLETES>
            <ATHLETE firstname="Isadora" lastname="Marafon" birthdate="2011-03-23" gender="F" nation="BRA" license="380287" swrid="5652623" athleteid="2035" externalid="380287">
              <RESULTS>
                <RESULT eventid="1065" points="407" swimtime="00:00:30.93" resultid="2036" heatid="2082" lane="4" entrytime="00:00:31.68" entrycourse="SCM" />
                <RESULT eventid="1081" points="397" swimtime="00:00:38.58" resultid="2037" heatid="2107" lane="2" entrytime="00:00:39.49" entrycourse="SCM" />
                <RESULT eventid="1103" points="356" swimtime="00:01:27.94" resultid="2038" heatid="2147" lane="7" entrytime="00:01:24.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6485" nation="BRA" region="PR" clubid="1137" name="Colégio Integrado, Campo Mourão" shortname="Cmou-Integrado,C">
          <ATHLETES>
            <ATHLETE firstname="Samuel" lastname="Massuda Santos" birthdate="2012-06-09" gender="M" nation="BRA" license="392189" swrid="5603872" athleteid="1138" externalid="392189">
              <RESULTS>
                <RESULT eventid="1063" points="215" swimtime="00:00:33.62" resultid="1139" heatid="2071" lane="4" />
                <RESULT eventid="1087" points="182" swimtime="00:01:19.05" resultid="1140" heatid="2120" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="168" swimtime="00:00:45.14" resultid="1141" heatid="2108" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Porto Schork Filho" birthdate="2012-12-28" gender="M" nation="BRA" license="V413906" athleteid="1142" externalid="V413906">
              <RESULTS>
                <RESULT eventid="1063" points="94" swimtime="00:00:44.28" resultid="1143" heatid="2071" lane="3" />
                <RESULT eventid="1087" points="79" swimtime="00:01:44.23" resultid="1144" heatid="2121" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="71" swimtime="00:01:00.14" resultid="1145" heatid="2109" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henry" lastname="Sadao Kague Da Silva" birthdate="2012-10-02" gender="M" nation="BRA" license="V413907" athleteid="1146" externalid="V413907">
              <RESULTS>
                <RESULT eventid="1063" points="79" swimtime="00:00:46.84" resultid="1147" heatid="2069" lane="6" />
                <RESULT eventid="1087" points="62" swimtime="00:01:53.12" resultid="1148" heatid="2121" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18831" nation="BRA" region="PR" clubid="1120" name="Colégio Estadual Profª. Elenir Linke, Cantagalo" shortname="Cant-Elenir Linke,Ce">
          <ATHLETES>
            <ATHLETE firstname="Yasmin" lastname="Daros" birthdate="2011-10-31" gender="F" nation="BRA" license="V413863" athleteid="1121" externalid="V413863">
              <RESULTS>
                <RESULT eventid="1065" status="DNS" swimtime="00:00:00.00" resultid="1122" heatid="2078" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Antonio Dalacort Gomes" birthdate="2012-08-17" gender="M" nation="BRA" license="V413939" athleteid="1125" externalid="V413939">
              <RESULTS>
                <RESULT eventid="1063" status="DNS" swimtime="00:00:00.00" resultid="1126" heatid="2069" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Vinicius Zapanovski De Oliveira" birthdate="2011-06-04" gender="M" nation="BRA" license="V413938" athleteid="1123" externalid="V413938">
              <RESULTS>
                <RESULT eventid="1063" status="DNS" swimtime="00:00:00.00" resultid="1124" heatid="2069" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11566" nation="BRA" region="PR" clubid="1487" name="Colégio Positivo Júnior, Curitiba" shortname="Ctba-Posi. Júnior,C">
          <ATHLETES>
            <ATHLETE firstname="Caua" lastname="Coelho" birthdate="2011-11-11" gender="M" nation="BRA" license="366889" swrid="5602527" athleteid="1488" externalid="366889">
              <RESULTS>
                <RESULT eventid="1075" points="295" swimtime="00:02:44.50" resultid="1489" heatid="2098" lane="5" entrytime="00:02:58.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:18.62" />
                    <SPLIT distance="150" swimtime="00:02:09.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="311" swimtime="00:01:06.17" resultid="1490" heatid="2124" lane="1" entrytime="00:01:04.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="265" swimtime="00:01:14.33" resultid="1491" heatid="2133" lane="8" entrytime="00:01:16.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gael" lastname="Gluck" birthdate="2011-01-28" gender="M" nation="BRA" license="366891" swrid="5588726" athleteid="1492" externalid="366891">
              <RESULTS>
                <RESULT eventid="1075" points="341" swimtime="00:02:36.83" resultid="1493" heatid="2099" lane="8" entrytime="00:02:53.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.29" />
                    <SPLIT distance="100" swimtime="00:01:16.36" />
                    <SPLIT distance="150" swimtime="00:02:00.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="312" swimtime="00:00:36.77" resultid="1494" heatid="2111" lane="2" entrytime="00:00:40.32" entrycourse="SCM" />
                <RESULT eventid="1105" points="330" swimtime="00:01:19.92" resultid="1495" heatid="2150" lane="2" entrytime="00:01:22.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="De Almeida Dias" birthdate="2012-02-18" gender="F" nation="BRA" license="369262" swrid="5588638" athleteid="1496" externalid="369262">
              <RESULTS>
                <RESULT eventid="1069" points="382" swimtime="00:01:15.59" resultid="1497" heatid="2089" lane="4" entrytime="00:01:18.41" entrycourse="SCM" />
                <RESULT eventid="1085" points="423" swimtime="00:01:06.90" resultid="1498" heatid="2117" lane="6" entrytime="00:01:05.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="345" swimtime="00:01:28.84" resultid="1499" heatid="2147" lane="1" entrytime="00:01:28.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="10585" nation="BRA" region="PR" clubid="1534" name="Colégio Estadual Santa Cândida, Curitiba" shortname="Ctba-Stª. Candida,Ce">
          <ATHLETES>
            <ATHLETE firstname="Heloisa" lastname="Daniele Silva" birthdate="2010-07-06" gender="F" nation="BRA" license="359593" swrid="5588628" athleteid="1535" externalid="359593" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1065" points="493" swimtime="00:00:29.01" resultid="1536" heatid="2083" lane="6" entrytime="00:00:30.08" entrycourse="SCM" />
                <RESULT eventid="1085" points="489" swimtime="00:01:03.76" resultid="1537" heatid="2117" lane="2" entrytime="00:01:05.94" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="388" swimtime="00:00:34.61" resultid="1538" heatid="2136" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13383" nation="BRA" region="PR" clubid="1183" name="Colégio Bom Jesus Água Verde, Curitiba" shortname="Ctba-Bj Água Verde,C">
          <ATHLETES>
            <ATHLETE firstname="Sarah" lastname="Emili Da Silva Gomes Xavier" birthdate="2010-09-08" gender="F" nation="BRA" license="372519" swrid="5717260" athleteid="1192" externalid="372519">
              <RESULTS>
                <RESULT eventid="1069" points="345" swimtime="00:01:18.23" resultid="1193" heatid="2089" lane="7" entrytime="00:01:23.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="409" swimtime="00:00:38.19" resultid="1194" heatid="2107" lane="7" entrytime="00:00:39.96" entrycourse="SCM" />
                <RESULT eventid="1099" points="341" swimtime="00:00:36.12" resultid="1195" heatid="2138" lane="6" entrytime="00:00:36.76" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Brandt De Macedo" birthdate="2010-01-13" gender="M" nation="BRA" license="338925" swrid="5588565" athleteid="1184" externalid="338925">
              <RESULTS>
                <RESULT eventid="1071" points="303" swimtime="00:00:32.36" resultid="1185" heatid="2091" lane="6" />
                <RESULT eventid="1087" points="400" swimtime="00:01:00.81" resultid="1186" heatid="2118" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="479" swimtime="00:04:31.20" resultid="1187" heatid="2102" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                    <SPLIT distance="100" swimtime="00:01:05.01" />
                    <SPLIT distance="150" swimtime="00:01:39.57" />
                    <SPLIT distance="200" swimtime="00:02:14.60" />
                    <SPLIT distance="250" swimtime="00:02:48.43" />
                    <SPLIT distance="300" swimtime="00:03:23.24" />
                    <SPLIT distance="350" swimtime="00:03:57.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Martynychen" birthdate="2011-12-19" gender="M" nation="BRA" license="366893" swrid="5602557" athleteid="1188" externalid="366893">
              <RESULTS>
                <RESULT eventid="1067" points="243" swimtime="00:01:17.36" resultid="1189" heatid="2084" lane="4" entrytime="00:01:22.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="279" swimtime="00:01:08.61" resultid="1190" heatid="2123" lane="1" entrytime="00:01:10.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="206" swimtime="00:00:37.42" resultid="1191" heatid="2142" lane="6" entrytime="00:00:39.99" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="14743" nation="BRA" region="PR" clubid="1914" name="Colégio Santo Inácio, Maringá" shortname="Mrga-Santo Inácio,C">
          <ATHLETES>
            <ATHLETE firstname="Lara" lastname="Constantino" birthdate="2012-06-02" gender="F" nation="BRA" license="382208" swrid="5420069" athleteid="1915" externalid="382208">
              <RESULTS>
                <RESULT eventid="1065" points="326" swimtime="00:00:33.31" resultid="1916" heatid="2081" lane="4" entrytime="00:00:35.62" entrycourse="SCM" />
                <RESULT eventid="1085" points="253" swimtime="00:01:19.36" resultid="1917" heatid="2114" lane="6" entrytime="00:01:28.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="322" swimtime="00:00:41.36" resultid="1918" heatid="2107" lane="8" entrytime="00:00:41.26" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17661" nation="BRA" region="PR" clubid="1992" name="Escola Literal, Pinhais" shortname="Pinh-Literal,E">
          <ATHLETES>
            <ATHLETE firstname="Lucca" lastname="Maceno Araujo" birthdate="2010-09-29" gender="M" nation="BRA" license="367056" swrid="5588788" athleteid="1993" externalid="367056">
              <RESULTS>
                <RESULT eventid="1071" points="345" swimtime="00:00:31.01" resultid="1994" heatid="2093" lane="2" entrytime="00:00:33.30" entrycourse="SCM" />
                <RESULT eventid="1087" points="373" swimtime="00:01:02.28" resultid="1995" heatid="2124" lane="8" entrytime="00:01:05.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="309" swimtime="00:01:10.63" resultid="1996" heatid="2133" lane="6" entrytime="00:01:13.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marjori" lastname="Leticia Oliveira" birthdate="2011-05-23" gender="F" nation="BRA" license="406869" swrid="5717279" athleteid="1997" externalid="406869">
              <RESULTS>
                <RESULT eventid="1065" points="275" swimtime="00:00:35.24" resultid="1998" heatid="2080" lane="4" entrytime="00:00:38.80" entrycourse="SCM" />
                <RESULT eventid="1085" status="DNS" swimtime="00:00:00.00" resultid="1999" heatid="2112" lane="5" />
                <RESULT eventid="1099" points="211" swimtime="00:00:42.41" resultid="2000" heatid="2137" lane="6" entrytime="00:00:44.10" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6486" nation="BRA" region="PR" clubid="1316" name="Colégio Da Polícia Militar, Curitiba" shortname="Ctba-Cpmpr,C">
          <ATHLETES>
            <ATHLETE firstname="Bruno" lastname="Gabriel Sarmento Buski" birthdate="2010-04-05" gender="M" nation="BRA" license="399533" swrid="5717264" athleteid="1317" externalid="399533">
              <RESULTS>
                <RESULT eventid="1079" points="364" swimtime="00:04:57.08" resultid="1318" heatid="2102" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                    <SPLIT distance="100" swimtime="00:01:07.48" />
                    <SPLIT distance="150" swimtime="00:01:45.56" />
                    <SPLIT distance="200" swimtime="00:02:23.97" />
                    <SPLIT distance="250" swimtime="00:03:02.80" />
                    <SPLIT distance="300" swimtime="00:03:41.39" />
                    <SPLIT distance="350" swimtime="00:04:20.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="264" swimtime="00:00:38.88" resultid="1319" heatid="2109" lane="7" />
                <RESULT eventid="1105" points="275" swimtime="00:01:24.91" resultid="1320" heatid="2149" lane="3" entrytime="00:01:30.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Rosa Silva" birthdate="2011-03-25" gender="F" nation="BRA" license="392120" swrid="5602579" athleteid="2054" externalid="392120">
              <RESULTS>
                <RESULT eventid="1081" points="186" swimtime="00:00:49.67" resultid="2056" heatid="2105" lane="5" entrytime="00:00:51.51" entrycourse="SCM" />
                <RESULT eventid="1085" status="RJC" swimtime="00:00:00.00" resultid="2057" entrytime="00:01:26.70" entrycourse="SCM" />
                <RESULT eventid="1089" status="RJC" swimtime="00:00:00.00" resultid="2058" />
                <RESULT eventid="1103" points="179" swimtime="00:01:50.64" resultid="2059" heatid="2145" lane="7" entrytime="00:01:48.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="226" swimtime="00:00:37.64" resultid="2060" heatid="2081" lane="8" entrytime="00:00:38.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Portella Da Silva" birthdate="2010-07-19" gender="M" nation="BRA" license="399534" swrid="5717288" athleteid="1321" externalid="399534">
              <RESULTS>
                <RESULT eventid="1063" points="196" swimtime="00:00:34.66" resultid="1322" heatid="2073" lane="2" entrytime="00:00:40.74" entrycourse="SCM" />
                <RESULT eventid="1083" points="201" swimtime="00:00:42.56" resultid="1323" heatid="2108" lane="6" />
                <RESULT eventid="1105" points="183" swimtime="00:01:37.35" resultid="1324" heatid="2148" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Yoshie Kimura" birthdate="2010-07-08" gender="F" nation="BRA" license="391142" swrid="5600277" athleteid="1325" externalid="391142">
              <RESULTS>
                <RESULT eventid="1089" points="347" swimtime="00:02:53.29" resultid="1326" heatid="2125" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.61" />
                    <SPLIT distance="100" swimtime="00:01:26.85" />
                    <SPLIT distance="150" swimtime="00:02:13.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1081" points="418" swimtime="00:00:37.92" resultid="1327" heatid="2107" lane="3" entrytime="00:00:38.22" entrycourse="SCM" />
                <RESULT eventid="1103" points="431" swimtime="00:01:22.50" resultid="1328" heatid="2147" lane="2" entrytime="00:01:24.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauan" lastname="De Lima Dos Reis" birthdate="2010-04-18" gender="M" nation="BRA" license="V413923" athleteid="1352" externalid="V413923">
              <RESULTS>
                <RESULT eventid="1063" points="247" swimtime="00:00:32.09" resultid="1353" heatid="2071" lane="8" />
                <RESULT eventid="1083" points="150" swimtime="00:00:46.87" resultid="1354" heatid="2108" lane="2" />
                <RESULT eventid="1105" points="165" swimtime="00:01:40.60" resultid="1355" heatid="2148" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Eduardo Santana" birthdate="2010-05-02" gender="M" nation="BRA" license="V413924" athleteid="1356" externalid="V413924">
              <RESULTS>
                <RESULT eventid="1087" points="194" swimtime="00:01:17.39" resultid="1357" heatid="2119" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1083" points="173" swimtime="00:00:44.71" resultid="1358" heatid="2108" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Micaella" lastname="Precybilovicz" birthdate="2010-10-06" gender="F" nation="BRA" license="V339343" athleteid="1329" externalid="V339343">
              <RESULTS>
                <RESULT eventid="1069" points="229" swimtime="00:01:29.63" resultid="1330" heatid="2088" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="272" swimtime="00:01:17.52" resultid="1331" heatid="2113" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="223" swimtime="00:00:41.58" resultid="1332" heatid="2137" lane="5" entrytime="00:00:42.08" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Bernardi Iurk" birthdate="2012-04-14" gender="M" nation="BRA" license="408687" swrid="5725984" athleteid="1333" externalid="408687">
              <RESULTS>
                <RESULT eventid="1087" points="148" swimtime="00:01:24.67" resultid="1334" heatid="2122" lane="2" entrytime="00:01:22.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1105" points="102" swimtime="00:01:57.99" resultid="1335" heatid="2148" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="107" swimtime="00:00:46.55" resultid="1336" heatid="2139" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Machado Oliveira" birthdate="2010-02-08" gender="F" nation="BRA" license="V413857" athleteid="1337" externalid="V413857">
              <RESULTS>
                <RESULT eventid="1065" points="162" swimtime="00:00:42.02" resultid="1338" heatid="2078" lane="1" />
                <RESULT eventid="1081" points="128" swimtime="00:00:56.23" resultid="1339" heatid="2105" lane="2" />
                <RESULT eventid="1103" status="DSQ" swimtime="00:02:03.66" resultid="1340" heatid="2144" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabio" lastname="Chiquito Do Brasil" birthdate="2011-05-11" gender="M" nation="BRA" license="V413921" athleteid="1345" externalid="V413921">
              <RESULTS>
                <RESULT eventid="1071" points="230" swimtime="00:00:35.46" resultid="1346" heatid="2091" lane="2" />
                <RESULT eventid="1063" points="301" swimtime="00:00:30.05" resultid="1347" heatid="2069" lane="7" />
                <RESULT eventid="1079" points="232" swimtime="00:05:45.18" resultid="1348" heatid="2101" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.12" />
                    <SPLIT distance="100" swimtime="00:01:21.55" />
                    <SPLIT distance="150" swimtime="00:02:04.60" />
                    <SPLIT distance="200" swimtime="00:02:48.44" />
                    <SPLIT distance="250" swimtime="00:03:32.62" />
                    <SPLIT distance="300" swimtime="00:04:16.95" />
                    <SPLIT distance="350" swimtime="00:05:01.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Zanatta Flizikowski" birthdate="2010-02-01" gender="F" nation="BRA" license="V413858" swrid="5588969" athleteid="1341" externalid="V413858">
              <RESULTS>
                <RESULT eventid="1073" points="344" swimtime="00:00:34.79" resultid="1342" heatid="2095" lane="8" />
                <RESULT eventid="1065" points="379" swimtime="00:00:31.68" resultid="1343" heatid="2078" lane="7" />
                <RESULT eventid="1085" points="391" swimtime="00:01:08.70" resultid="1344" heatid="2112" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Goncalves Plocharski" birthdate="2011-08-01" gender="M" nation="BRA" license="V413922" athleteid="1349" externalid="V413922">
              <RESULTS>
                <RESULT eventid="1063" points="157" swimtime="00:00:37.36" resultid="1350" heatid="2072" lane="6" />
                <RESULT eventid="1087" points="110" swimtime="00:01:33.44" resultid="1351" heatid="2119" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="M" name="CTBA-POL. MILITAR,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1091" points="258" swimtime="00:02:08.33" resultid="1361" heatid="2128" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.36" />
                    <SPLIT distance="100" swimtime="00:01:08.30" />
                    <SPLIT distance="150" swimtime="00:01:38.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1321" number="1" />
                    <RELAYPOSITION athleteid="1352" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1317" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1345" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1109" points="228" swimtime="00:02:26.70" resultid="1362" heatid="2152" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.05" />
                    <SPLIT distance="100" swimtime="00:01:17.93" />
                    <SPLIT distance="150" swimtime="00:01:53.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1321" number="1" />
                    <RELAYPOSITION athleteid="1317" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1345" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1352" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="CTBA-POL. MILITAR,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1093" points="292" swimtime="00:02:19.29" resultid="1359" heatid="2129" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.51" />
                    <SPLIT distance="100" swimtime="00:01:16.61" />
                    <SPLIT distance="150" swimtime="00:01:47.99" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1337" number="1" />
                    <RELAYPOSITION athleteid="1329" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1325" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1341" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1107" points="277" swimtime="00:02:36.88" resultid="1360" heatid="2151" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.55" />
                    <SPLIT distance="100" swimtime="00:01:19.94" />
                    <SPLIT distance="150" swimtime="00:01:55.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1329" number="1" />
                    <RELAYPOSITION athleteid="1325" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1341" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1337" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="CTBA-POL. MILITAR,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1077" points="258" swimtime="00:02:29.33" resultid="1363" heatid="2100" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.01" />
                    <SPLIT distance="100" swimtime="00:01:19.43" />
                    <SPLIT distance="150" swimtime="00:01:55.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1329" number="1" />
                    <RELAYPOSITION athleteid="1325" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1317" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1321" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="13978" nation="BRA" region="PR" clubid="1464" name="Colégio Modelo Do Paraná, Curitiba" shortname="Ctba-Modelo,C">
          <ATHLETES>
            <ATHLETE firstname="Bernardo" lastname="Lopes Rempel" birthdate="2010-09-25" gender="M" nation="BRA" license="399739" swrid="5653294" athleteid="1465" externalid="399739">
              <RESULTS>
                <RESULT eventid="1067" points="190" swimtime="00:01:24.05" resultid="1466" heatid="2084" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="250" swimtime="00:00:31.96" resultid="1467" heatid="2071" lane="6" />
                <RESULT eventid="1101" points="212" swimtime="00:00:37.06" resultid="1468" heatid="2141" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="9870" nation="BRA" region="PR" clubid="1780" name="Colégio Anglo, Maringá" shortname="Mrga-Anglo,C">
          <ATHLETES>
            <ATHLETE firstname="Caua" lastname="Pazinato" birthdate="2011-01-05" gender="M" nation="BRA" license="368149" swrid="5603889" athleteid="1781" externalid="368149">
              <RESULTS>
                <RESULT eventid="1067" points="234" swimtime="00:01:18.38" resultid="1782" heatid="2085" lane="1" entrytime="00:01:18.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="311" swimtime="00:00:29.74" resultid="1783" heatid="2075" lane="6" entrytime="00:00:30.40" entrycourse="SCM" />
                <RESULT eventid="1087" points="300" swimtime="00:01:06.91" resultid="1784" heatid="2123" lane="5" entrytime="00:01:06.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11380" nation="BRA" region="PR" clubid="1544" name="Colégio Nossa Srª. Auxiliadora, Cascavel" shortname="Cvel-Auxiliadora,C">
          <ATHLETES>
            <ATHLETE firstname="João" lastname="Pedro Serafini" birthdate="2012-05-15" gender="M" nation="BRA" license="365488" swrid="5596924" athleteid="1549" externalid="365488">
              <RESULTS>
                <RESULT eventid="1075" points="170" swimtime="00:03:17.77" resultid="1550" heatid="2097" lane="4" entrytime="00:03:19.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.07" />
                    <SPLIT distance="100" swimtime="00:01:36.39" />
                    <SPLIT distance="150" swimtime="00:02:36.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="207" swimtime="00:05:58.70" resultid="1551" heatid="2153" lane="4" entrytime="00:06:08.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                    <SPLIT distance="100" swimtime="00:01:24.68" />
                    <SPLIT distance="150" swimtime="00:02:11.43" />
                    <SPLIT distance="200" swimtime="00:02:58.23" />
                    <SPLIT distance="250" swimtime="00:03:45.42" />
                    <SPLIT distance="300" swimtime="00:04:30.60" />
                    <SPLIT distance="350" swimtime="00:05:16.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="114" swimtime="00:01:38.28" resultid="1552" heatid="2132" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laisa" lastname="Bernardini" birthdate="2012-06-25" gender="F" nation="BRA" license="390843" swrid="5596872" athleteid="1553" externalid="390843">
              <RESULTS>
                <RESULT eventid="1073" points="160" swimtime="00:00:44.84" resultid="1554" heatid="2095" lane="2" entrytime="00:00:47.34" entrycourse="SCM" />
                <RESULT eventid="1089" points="229" swimtime="00:03:19.01" resultid="1555" heatid="2126" lane="7" entrytime="00:03:28.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.28" />
                    <SPLIT distance="100" swimtime="00:01:36.19" />
                    <SPLIT distance="150" swimtime="00:02:33.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="198" swimtime="00:01:46.95" resultid="1556" heatid="2145" lane="2" entrytime="00:01:47.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raul" lastname="Bonamigo" birthdate="2010-12-01" gender="M" nation="BRA" license="344397" swrid="5588559" athleteid="1545" externalid="344397">
              <RESULTS>
                <RESULT eventid="1067" points="368" swimtime="00:01:07.42" resultid="1546" heatid="2086" lane="1" entrytime="00:01:10.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="400" swimtime="00:02:28.73" resultid="1547" heatid="2099" lane="6" entrytime="00:02:32.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="100" swimtime="00:01:09.57" />
                    <SPLIT distance="150" swimtime="00:01:54.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="393" swimtime="00:01:01.17" resultid="1548" heatid="2120" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2670" nation="BRA" region="PR" clubid="1422" name="Colégio Marista Paranaense, Curitiba" shortname="Ctba-Marista Pr,C">
          <ATHLETES>
            <ATHLETE firstname="Mariana" lastname="Stoberl" birthdate="2010-07-09" gender="F" nation="BRA" license="356250" swrid="5600265" athleteid="1423" externalid="356250">
              <RESULTS>
                <RESULT eventid="1065" points="473" swimtime="00:00:29.41" resultid="1424" heatid="2083" lane="5" entrytime="00:00:29.79" entrycourse="SCM" />
                <RESULT eventid="1085" points="503" swimtime="00:01:03.17" resultid="1425" heatid="2117" lane="4" entrytime="00:01:04.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="384" swimtime="00:00:34.71" resultid="1426" heatid="2138" lane="3" entrytime="00:00:35.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Cabrini Vieira" birthdate="2012-02-11" gender="F" nation="BRA" license="376961" swrid="5588571" athleteid="1443" externalid="376961">
              <RESULTS>
                <RESULT eventid="1069" points="334" swimtime="00:01:19.09" resultid="1444" heatid="2090" lane="2" entrytime="00:01:15.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="415" swimtime="00:00:30.74" resultid="1445" heatid="2082" lane="5" entrytime="00:00:31.88" entrycourse="SCM" />
                <RESULT eventid="1085" points="389" swimtime="00:01:08.82" resultid="1446" heatid="2117" lane="8" entrytime="00:01:06.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Salomao" birthdate="2012-05-07" gender="M" nation="BRA" license="369261" swrid="5602581" athleteid="1431" externalid="369261">
              <RESULTS>
                <RESULT eventid="1071" points="194" swimtime="00:00:37.55" resultid="1432" heatid="2092" lane="3" entrytime="00:00:37.94" entrycourse="SCM" />
                <RESULT eventid="1063" points="233" swimtime="00:00:32.74" resultid="1433" heatid="2074" lane="5" entrytime="00:00:32.07" entrycourse="SCM" />
                <RESULT eventid="1087" points="253" swimtime="00:01:10.84" resultid="1434" heatid="2123" lane="2" entrytime="00:01:09.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Karam Barbosa Lima" birthdate="2012-12-11" gender="F" nation="BRA" license="376956" swrid="5588758" athleteid="1439" externalid="376956">
              <RESULTS>
                <RESULT eventid="1069" points="260" swimtime="00:01:25.91" resultid="1440" heatid="2089" lane="1" entrytime="00:01:23.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1061" points="295" swimtime="00:05:47.35" resultid="1441" heatid="2068" lane="1" entrytime="00:05:37.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.54" />
                    <SPLIT distance="100" swimtime="00:01:19.49" />
                    <SPLIT distance="150" swimtime="00:02:04.04" />
                    <SPLIT distance="200" swimtime="00:02:48.94" />
                    <SPLIT distance="250" swimtime="00:03:33.95" />
                    <SPLIT distance="300" swimtime="00:04:18.99" />
                    <SPLIT distance="350" swimtime="00:05:03.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="267" swimtime="00:01:17.96" resultid="1442" heatid="2116" lane="1" entrytime="00:01:12.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Clivatti" birthdate="2010-05-24" gender="M" nation="BRA" license="368007" swrid="5600139" athleteid="1427" externalid="368007">
              <RESULTS>
                <RESULT eventid="1063" points="407" swimtime="00:00:27.20" resultid="1428" heatid="2076" lane="3" entrytime="00:00:27.48" entrycourse="SCM" />
                <RESULT eventid="1087" points="460" swimtime="00:00:58.07" resultid="1429" heatid="2124" lane="5" entrytime="00:00:59.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1079" points="512" swimtime="00:04:25.22" resultid="1430" heatid="2103" lane="3" entrytime="00:04:34.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                    <SPLIT distance="100" swimtime="00:01:03.29" />
                    <SPLIT distance="150" swimtime="00:01:37.09" />
                    <SPLIT distance="200" swimtime="00:02:10.95" />
                    <SPLIT distance="250" swimtime="00:02:45.01" />
                    <SPLIT distance="300" swimtime="00:03:18.61" />
                    <SPLIT distance="350" swimtime="00:03:52.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Tallao Benke" birthdate="2012-01-02" gender="F" nation="BRA" license="376984" swrid="5588931" athleteid="1447" externalid="376984">
              <RESULTS>
                <RESULT eventid="1069" points="436" swimtime="00:01:12.35" resultid="1448" heatid="2090" lane="3" entrytime="00:01:14.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1061" points="513" swimtime="00:04:48.93" resultid="1449" heatid="2068" lane="4" entrytime="00:04:48.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                    <SPLIT distance="100" swimtime="00:01:07.61" />
                    <SPLIT distance="150" swimtime="00:01:44.58" />
                    <SPLIT distance="200" swimtime="00:02:21.33" />
                    <SPLIT distance="250" swimtime="00:02:58.12" />
                    <SPLIT distance="300" swimtime="00:03:35.39" />
                    <SPLIT distance="350" swimtime="00:04:12.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1095" points="439" swimtime="00:01:11.07" resultid="1450" heatid="2131" lane="5" entrytime="00:01:10.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Szpak De Vasconcelos" birthdate="2012-06-29" gender="M" nation="BRA" license="369271" swrid="5588928" athleteid="1435" externalid="369271">
              <RESULTS>
                <RESULT eventid="1063" points="289" swimtime="00:00:30.49" resultid="1436" heatid="2075" lane="3" entrytime="00:00:29.99" entrycourse="SCM" />
                <RESULT eventid="1083" points="273" swimtime="00:00:38.45" resultid="1437" heatid="2111" lane="6" entrytime="00:00:38.19" entrycourse="SCM" />
                <RESULT eventid="1105" points="256" swimtime="00:01:27.04" resultid="1438" heatid="2150" lane="7" entrytime="00:01:23.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F">
              <RESULTS>
                <RESULT eventid="1107" status="DNS" swimtime="00:00:00.00" resultid="2154" heatid="2151" lane="5" late="yes">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1443" number="1" />
                    <RELAYPOSITION athleteid="1439" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1447" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1423" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="F" name="CTBA-MARISTA PR,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1093" status="DSQ" swimtime="00:02:03.98" resultid="1451" heatid="2129" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                    <SPLIT distance="100" swimtime="00:01:03.24" />
                    <SPLIT distance="150" swimtime="00:01:34.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1447" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="1439" number="2" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1443" number="3" reactiontime="0" status="DSQ" />
                    <RELAYPOSITION athleteid="1423" number="4" reactiontime="0" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="-1" agetotalmax="-1" agetotalmin="-1" gender="X" name="CTBA-MARISTA PR,C &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1077" points="355" swimtime="00:02:14.37" resultid="1453" heatid="2100" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                    <SPLIT distance="100" swimtime="00:01:15.37" />
                    <SPLIT distance="150" swimtime="00:01:46.26" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="1443" number="1" />
                    <RELAYPOSITION athleteid="1435" number="2" reactiontime="0" />
                    <RELAYPOSITION athleteid="1447" number="3" reactiontime="0" />
                    <RELAYPOSITION athleteid="1427" number="4" reactiontime="0" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="18818" nation="BRA" region="PR" clubid="2039" name="Colégio Vila Militar (CVM), Toledo" shortname="Tole-Vila Militar,C">
          <ATHLETES>
            <ATHLETE firstname="Eduardo" lastname="Murilo Fernandes Apolinario" birthdate="2011-05-13" gender="M" nation="BRA" license="V413931" athleteid="2040" externalid="V413931">
              <RESULTS>
                <RESULT eventid="1063" points="32" swimtime="00:01:03.05" resultid="2041" heatid="2070" lane="1" />
                <RESULT eventid="1101" status="DSQ" swimtime="00:01:17.33" resultid="2042" heatid="2140" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17649" nation="BRA" region="PR" clubid="1802" name="Colégio Criarte, Maringá" shortname="Mrga-Criarte,C">
          <ATHLETES>
            <ATHLETE firstname="Pietro" lastname="Nabas De Assis" birthdate="2011-07-09" gender="M" nation="BRA" license="366968" swrid="5603878" athleteid="1803" externalid="366968">
              <RESULTS>
                <RESULT eventid="1083" points="363" swimtime="00:00:34.95" resultid="1804" heatid="2111" lane="5" entrytime="00:00:37.30" entrycourse="SCM" />
                <RESULT eventid="1105" points="347" swimtime="00:01:18.60" resultid="1805" heatid="2150" lane="3" entrytime="00:01:19.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.42" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="4222" nation="BRA" region="PR" clubid="1660" name="Colégio Bertoni Internacional, Foz Do Iguaçu" shortname="Fozi-Bertoni Int.,C">
          <ATHLETES>
            <ATHLETE firstname="Edward" lastname="Mikael De Lima" birthdate="2012-03-11" gender="M" nation="BRA" license="376445" swrid="5588816" athleteid="1661" externalid="376445" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1063" status="DSQ" swimtime="00:00:27.97" resultid="1662" heatid="2076" lane="5" entrytime="00:00:27.35" entrycourse="SCM" />
                <RESULT eventid="1079" points="364" swimtime="00:04:57.00" resultid="1663" heatid="2103" lane="2" entrytime="00:04:58.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:08.67" />
                    <SPLIT distance="150" swimtime="00:01:46.44" />
                    <SPLIT distance="200" swimtime="00:02:25.03" />
                    <SPLIT distance="250" swimtime="00:03:03.44" />
                    <SPLIT distance="300" swimtime="00:03:42.65" />
                    <SPLIT distance="350" swimtime="00:04:20.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1097" points="253" swimtime="00:01:15.47" resultid="1664" heatid="2132" lane="5" entrytime="00:01:18.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13450" nation="BRA" region="PR" clubid="1730" name="Colégio Anglo Londrinense, Londrina" shortname="Ldna-Anglo.Londri.,C">
          <ATHLETES>
            <ATHLETE firstname="Luisa" lastname="Genvigir" birthdate="2011-04-02" gender="F" nation="BRA" license="V413856" athleteid="1739" externalid="V413856">
              <RESULTS>
                <RESULT eventid="1065" points="178" swimtime="00:00:40.76" resultid="1740" heatid="2079" lane="6" />
                <RESULT eventid="1085" points="158" swimtime="00:01:32.95" resultid="1741" heatid="2113" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" status="DNS" swimtime="00:00:00.00" resultid="1742" heatid="2135" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Takemura Couto" birthdate="2010-02-08" gender="F" nation="BRA" license="376950" swrid="5603919" athleteid="1735" externalid="376950">
              <RESULTS>
                <RESULT eventid="1065" points="487" swimtime="00:00:29.14" resultid="1736" heatid="2083" lane="4" entrytime="00:00:29.49" entrycourse="SCM" />
                <RESULT eventid="1085" points="466" swimtime="00:01:04.79" resultid="1737" heatid="2117" lane="5" entrytime="00:01:05.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="303" swimtime="00:01:32.77" resultid="1738" heatid="2146" lane="2" entrytime="00:01:35.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Poletti Veiga" birthdate="2010-10-01" gender="F" nation="BRA" license="376951" swrid="5603895" athleteid="1731" externalid="376951">
              <RESULTS>
                <RESULT eventid="1069" points="367" swimtime="00:01:16.66" resultid="1732" heatid="2090" lane="7" entrytime="00:01:16.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="408" swimtime="00:01:07.73" resultid="1733" heatid="2117" lane="7" entrytime="00:01:05.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="381" swimtime="00:00:34.82" resultid="1734" heatid="2134" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13980" nation="BRA" region="PR" clubid="1680" name="CCM Presidente Costa E Silva, Foz Do Iguaçu" shortname="Fozi-Costa Silva,CCM">
          <ATHLETES>
            <ATHLETE firstname="Faisal" lastname="Basem Ghotme" birthdate="2010-12-18" gender="M" nation="BRA" license="390809" swrid="5596871" athleteid="1681" externalid="390809" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1063" points="439" swimtime="00:00:26.52" resultid="1682" heatid="2076" lane="6" entrytime="00:00:27.65" entrycourse="SCM" />
                <RESULT eventid="1087" points="396" swimtime="00:01:01.05" resultid="1683" heatid="2124" lane="3" entrytime="00:01:01.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1101" points="378" swimtime="00:00:30.57" resultid="1684" heatid="2141" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16472" nation="BRA" region="PR" clubid="1919" name="Colegio Est Prof Agostinho Pereira, Pato Branco Pr" shortname="Pbco-Agostinho F.,Ce">
          <ATHLETES>
            <ATHLETE firstname="Otavio" lastname="Augusto Bergamaschi" birthdate="2010-11-08" gender="M" nation="BRA" license="V399600" athleteid="1920" externalid="V399600">
              <RESULTS>
                <RESULT eventid="1063" points="257" swimtime="00:00:31.68" resultid="1921" heatid="2073" lane="4" entrytime="00:00:35.26" entrycourse="SCM" />
                <RESULT eventid="1083" points="212" swimtime="00:00:41.80" resultid="1922" heatid="2110" lane="3" entrytime="00:00:43.50" entrycourse="SCM" />
                <RESULT eventid="1101" points="208" swimtime="00:00:37.26" resultid="1923" heatid="2142" lane="2" entrytime="00:00:41.05" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Orliczek Couto" birthdate="2011-05-13" gender="M" nation="BRA" license="V413940" athleteid="1924" externalid="V413940">
              <RESULTS>
                <RESULT eventid="1063" status="WDR" swimtime="00:00:00.00" resultid="1925" />
                <RESULT eventid="1101" status="WDR" swimtime="00:00:00.00" resultid="1926" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2654" nation="BRA" region="PR" clubid="1891" name="Colégio Platão, Maringá" shortname="Mrga-Platão,C">
          <ATHLETES>
            <ATHLETE firstname="Rafael" lastname="Britto" birthdate="2012-10-04" gender="M" nation="BRA" license="378350" swrid="5588566" athleteid="1896" externalid="378350">
              <RESULTS>
                <RESULT eventid="1067" status="DNS" swimtime="00:00:00.00" resultid="1897" heatid="2085" lane="6" entrytime="00:01:15.63" entrycourse="SCM" />
                <RESULT eventid="1075" status="DNS" swimtime="00:00:00.00" resultid="1898" heatid="2098" lane="6" entrytime="00:03:01.68" entrycourse="SCM" />
                <RESULT eventid="1101" points="255" swimtime="00:00:34.84" resultid="1899" heatid="2143" lane="1" entrytime="00:00:36.08" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benicio" lastname="Garcia" birthdate="2011-09-09" gender="M" nation="BRA" license="378347" swrid="5603842" athleteid="1892" externalid="378347">
              <RESULTS>
                <RESULT eventid="1067" points="224" swimtime="00:01:19.51" resultid="1893" heatid="2085" lane="2" entrytime="00:01:17.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1075" points="222" swimtime="00:03:00.93" resultid="1894" heatid="2098" lane="7" entrytime="00:03:13.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.22" />
                    <SPLIT distance="100" swimtime="00:01:22.33" />
                    <SPLIT distance="150" swimtime="00:01:52.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1087" points="254" swimtime="00:01:10.76" resultid="1895" heatid="2123" lane="7" entrytime="00:01:10.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="17657" nation="BRA" region="PR" clubid="1743" name="Colégio Luterano Rui Barbosa, M. Cândido Rondon" shortname="Mcro-Luterano Rui.,C">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Fernanda Ribeiro Do Prado" birthdate="2011-03-18" gender="F" nation="BRA" license="V399531" athleteid="1744" externalid="V399531">
              <RESULTS>
                <RESULT eventid="1065" points="168" swimtime="00:00:41.52" resultid="1745" heatid="2078" lane="4" />
                <RESULT eventid="1085" points="136" swimtime="00:01:37.63" resultid="1746" heatid="2113" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" status="DSQ" swimtime="00:00:51.68" resultid="1747" heatid="2135" lane="7" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13438" nation="BRA" region="PR" clubid="1519" name="Colégio Santo Anjo, Curitiba" shortname="Ctba-Santo Anjo,C">
          <ATHLETES>
            <ATHLETE firstname="Laura" lastname="Lazzarotti Matias" birthdate="2012-03-19" gender="F" nation="BRA" license="391026" swrid="5602552" athleteid="1520" externalid="391026">
              <RESULTS>
                <RESULT eventid="1069" points="296" swimtime="00:01:22.31" resultid="1521" heatid="2090" lane="8" entrytime="00:01:17.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1103" points="256" swimtime="00:01:38.09" resultid="1522" heatid="2146" lane="7" entrytime="00:01:35.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1099" points="351" swimtime="00:00:35.77" resultid="1523" heatid="2138" lane="5" entrytime="00:00:34.84" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="18824" nation="BRA" region="PR" clubid="1927" name="Escola Crescer, Pato Branco" shortname="Pbco-Crescer,E">
          <ATHLETES>
            <ATHLETE firstname="Sofia" lastname="Barreto" birthdate="2011-05-11" gender="F" nation="BRA" license="V413867" athleteid="1928" externalid="V413867">
              <RESULTS>
                <RESULT eventid="1065" points="185" swimtime="00:00:40.18" resultid="1929" heatid="2077" lane="4" />
                <RESULT eventid="1099" points="143" swimtime="00:00:48.23" resultid="1930" heatid="2134" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="14735" nation="BRA" region="PR" clubid="1726" name="2º Colégio Da Polícia Militar, Londrina" shortname="Ldna-2ºcpmpr,C">
          <ATHLETES>
            <ATHLETE firstname="Brenda" lastname="Paulino Rodrigues Reina" birthdate="2012-06-05" gender="F" nation="BRA" license="V413891" athleteid="1727" externalid="V413891">
              <RESULTS>
                <RESULT eventid="1065" points="227" swimtime="00:00:37.55" resultid="1728" heatid="2082" lane="2" />
                <RESULT eventid="1099" points="224" swimtime="00:00:41.52" resultid="1729" heatid="2134" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="6473" nation="BRA" region="PR" clubid="1665" name="Colégio Caesp, Foz Do Iguaçu" shortname="Fozi-Caesp,C">
          <ATHLETES>
            <ATHLETE firstname="Ysadora" lastname="Bertoldo" birthdate="2010-04-09" gender="F" nation="BRA" license="376444" swrid="5588553" athleteid="1666" externalid="376444" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1061" points="450" swimtime="00:05:01.80" resultid="1667" heatid="2068" lane="2" entrytime="00:05:25.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.64" />
                    <SPLIT distance="100" swimtime="00:01:13.92" />
                    <SPLIT distance="150" swimtime="00:01:52.52" />
                    <SPLIT distance="200" swimtime="00:02:30.86" />
                    <SPLIT distance="250" swimtime="00:03:08.83" />
                    <SPLIT distance="300" swimtime="00:03:47.05" />
                    <SPLIT distance="350" swimtime="00:04:25.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1065" points="349" swimtime="00:00:32.55" resultid="1668" heatid="2082" lane="8" entrytime="00:00:34.24" entrycourse="SCM" />
                <RESULT eventid="1085" points="377" swimtime="00:01:09.54" resultid="1669" heatid="2116" lane="8" entrytime="00:01:12.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="8446" nation="BRA" region="PR" clubid="1806" name="Colégio Cristão Integrado, Maringá" shortname="Mrga-Cristao Integ,C">
          <ATHLETES>
            <ATHLETE firstname="Felype" lastname="Gongora Zago" birthdate="2011-09-14" gender="M" nation="BRA" license="392099" swrid="5603848" athleteid="1807" externalid="392099">
              <RESULTS>
                <RESULT eventid="1071" points="221" swimtime="00:00:35.97" resultid="1808" heatid="2091" lane="3" />
                <RESULT eventid="1063" points="225" swimtime="00:00:33.10" resultid="1809" heatid="2074" lane="7" entrytime="00:00:33.30" entrycourse="SCM" />
                <RESULT eventid="1087" points="204" swimtime="00:01:16.06" resultid="1810" heatid="2122" lane="3" entrytime="00:01:16.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13444" nation="BRA" region="PR" clubid="1943" name="Escola Estadual Medalha Milagrosa, Ponta Grossa" shortname="Pgro-Medalha MIL.,Ee">
          <ATHLETES>
            <ATHLETE firstname="Joao" lastname="Vyctor Cadene Brantes" birthdate="2011-03-04" gender="M" nation="BRA" license="V413927" athleteid="1944" externalid="V413927">
              <RESULTS>
                <RESULT eventid="1063" points="203" swimtime="00:00:34.30" resultid="1945" heatid="2069" lane="2" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="8871" nation="BRA" region="PR" clubid="1454" name="Colégio Marista Santa Maria, Curitiba" shortname="Ctba-Marista St.Mª,C">
          <ATHLETES>
            <ATHLETE firstname="Isadora" lastname="Albuquerque" birthdate="2012-08-17" gender="F" nation="BRA" license="369275" swrid="5602507" athleteid="1455" externalid="369275">
              <RESULTS>
                <RESULT eventid="1073" status="DNS" swimtime="00:00:00.00" resultid="1456" heatid="2096" lane="7" entrytime="00:00:36.53" entrycourse="SCM" />
                <RESULT eventid="1081" status="DNS" swimtime="00:00:00.00" resultid="1457" heatid="2107" lane="4" entrytime="00:00:37.52" entrycourse="SCM" />
                <RESULT eventid="1103" status="DNS" swimtime="00:00:00.00" resultid="1458" heatid="2147" lane="3" entrytime="00:01:22.87" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2273" nation="BRA" region="PR" clubid="1845" name="Colégio Marista, Maringá" shortname="Mrga-Marista,C">
          <ATHLETES>
            <ATHLETE firstname="Bruna" lastname="Scalise Drapzichinski" birthdate="2012-03-07" gender="F" nation="BRA" license="378349" swrid="5603909" athleteid="1846" externalid="378349">
              <RESULTS>
                <RESULT eventid="1073" points="334" swimtime="00:00:35.11" resultid="1847" heatid="2096" lane="6" entrytime="00:00:35.33" entrycourse="SCM" />
                <RESULT eventid="1081" points="424" swimtime="00:00:37.74" resultid="1848" heatid="2107" lane="6" entrytime="00:00:38.38" entrycourse="SCM" />
                <RESULT eventid="1103" points="393" swimtime="00:01:25.11" resultid="1849" heatid="2146" lane="6" entrytime="00:01:35.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Traci Rodrigues" birthdate="2011-03-06" gender="M" nation="BRA" license="406927" swrid="5718893" athleteid="1850" externalid="406927">
              <RESULTS>
                <RESULT eventid="1063" status="SICK" swimtime="00:00:00.00" resultid="1851" entrytime="00:00:37.34" entrycourse="SCM" />
                <RESULT eventid="1087" status="SICK" swimtime="00:00:00.00" resultid="1852" />
                <RESULT eventid="1083" status="SICK" swimtime="00:00:00.00" resultid="1853" />
                <RESULT eventid="1105" status="SICK" swimtime="00:00:00.00" resultid="1854" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
