<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.79293">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Curitiba" name="Torneio Regional da 1ª Região (Pré-Mirim/Petiz)" course="SCM" deadline="2024-03-31" entrystartdate="2024-03-26" entrytype="INVITATION" hostclub="Clube Curitibano" hostclub.url="https://clubecuritibano.com.br/" number="38305" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/evento/natacao/38305" startmethod="1" timing="AUTOMATIC" masters="F" withdrawuntil="2024-04-02" state="PR" nation="BRA">
      <AGEDATE value="2024-04-06" type="YEAR" />
      <POOL name="Parque Aquático do Clube Curitibano" lanemin="1" lanemax="8" />
      <FACILITY city="Curitiba" name="Parque Aquático do Clube Curitibano" nation="BRA" state="PR" street="Avenida Presidente Getúlio Vargas, 2857" street2="Água Verde" zip="80240-040" />
      <POINTTABLE pointtableid="3016" name="FINA Point Scoring" version="2023" />
      <QUALIFY from="2023-04-06" until="2024-04-05" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-04-06" daytime="09:10" endtime="12:01" number="1" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1060" daytime="09:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1062" daytime="09:10" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1063" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1064" daytime="09:10" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1065" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1872" />
                    <RANKING order="2" place="2" resultid="1659" />
                    <RANKING order="3" place="3" resultid="1881" />
                    <RANKING order="4" place="4" resultid="1699" />
                    <RANKING order="5" place="5" resultid="1640" />
                    <RANKING order="6" place="6" resultid="2065" />
                    <RANKING order="7" place="7" resultid="1751" />
                    <RANKING order="8" place="8" resultid="1694" />
                    <RANKING order="9" place="9" resultid="1635" />
                    <RANKING order="10" place="10" resultid="1674" />
                    <RANKING order="11" place="11" resultid="1796" />
                    <RANKING order="12" place="-1" resultid="1704" />
                    <RANKING order="13" place="-1" resultid="1724" />
                    <RANKING order="14" place="-1" resultid="1766" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1066" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1913" />
                    <RANKING order="2" place="2" resultid="1515" />
                    <RANKING order="3" place="3" resultid="2004" />
                    <RANKING order="4" place="4" resultid="2060" />
                    <RANKING order="5" place="5" resultid="1595" />
                    <RANKING order="6" place="6" resultid="1575" />
                    <RANKING order="7" place="7" resultid="1610" />
                    <RANKING order="8" place="8" resultid="1620" />
                    <RANKING order="9" place="9" resultid="1664" />
                    <RANKING order="10" place="10" resultid="1520" />
                    <RANKING order="11" place="11" resultid="1157" />
                    <RANKING order="12" place="12" resultid="2009" />
                    <RANKING order="13" place="13" resultid="1555" />
                    <RANKING order="14" place="14" resultid="1709" />
                    <RANKING order="15" place="15" resultid="1580" />
                    <RANKING order="16" place="16" resultid="1243" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2072" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2073" daytime="09:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2074" daytime="09:22" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2075" daytime="09:28" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1067" daytime="09:32" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1068" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1645" />
                    <RANKING order="2" place="2" resultid="1991" />
                    <RANKING order="3" place="3" resultid="1630" />
                    <RANKING order="4" place="4" resultid="1689" />
                    <RANKING order="5" place="5" resultid="1756" />
                    <RANKING order="6" place="6" resultid="1719" />
                    <RANKING order="7" place="7" resultid="1741" />
                    <RANKING order="8" place="8" resultid="1761" />
                    <RANKING order="9" place="9" resultid="1776" />
                    <RANKING order="10" place="10" resultid="1781" />
                    <RANKING order="11" place="-1" resultid="1729" />
                    <RANKING order="12" place="-1" resultid="1805" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1505" />
                    <RANKING order="2" place="2" resultid="1590" />
                    <RANKING order="3" place="3" resultid="1714" />
                    <RANKING order="4" place="4" resultid="1535" />
                    <RANKING order="5" place="5" resultid="1525" />
                    <RANKING order="6" place="6" resultid="1952" />
                    <RANKING order="7" place="7" resultid="1530" />
                    <RANKING order="8" place="8" resultid="1585" />
                    <RANKING order="9" place="9" resultid="2022" />
                    <RANKING order="10" place="10" resultid="1182" />
                    <RANKING order="11" place="11" resultid="1943" />
                    <RANKING order="12" place="12" resultid="1565" />
                    <RANKING order="13" place="13" resultid="2014" />
                    <RANKING order="14" place="14" resultid="1968" />
                    <RANKING order="15" place="15" resultid="2027" />
                    <RANKING order="16" place="16" resultid="1545" />
                    <RANKING order="17" place="17" resultid="2036" />
                    <RANKING order="18" place="18" resultid="1550" />
                    <RANKING order="19" place="-1" resultid="1570" />
                    <RANKING order="20" place="-1" resultid="1654" />
                    <RANKING order="21" place="-1" resultid="1669" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2076" daytime="09:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2077" daytime="09:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2078" daytime="09:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2079" daytime="09:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2080" daytime="09:54" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1070" daytime="10:00" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1071" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1384" />
                    <RANKING order="2" place="2" resultid="1827" />
                    <RANKING order="3" place="3" resultid="1938" />
                    <RANKING order="4" place="4" resultid="1491" />
                    <RANKING order="5" place="5" resultid="1786" />
                    <RANKING order="6" place="6" resultid="1918" />
                    <RANKING order="7" place="7" resultid="1438" />
                    <RANKING order="8" place="8" resultid="1510" />
                    <RANKING order="9" place="9" resultid="1560" />
                    <RANKING order="10" place="-1" resultid="1423" />
                    <RANKING order="11" place="-1" resultid="1605" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1462" />
                    <RANKING order="2" place="2" resultid="1306" />
                    <RANKING order="3" place="3" resultid="1301" />
                    <RANKING order="4" place="4" resultid="1341" />
                    <RANKING order="5" place="5" resultid="1361" />
                    <RANKING order="6" place="6" resultid="1600" />
                    <RANKING order="7" place="7" resultid="1389" />
                    <RANKING order="8" place="8" resultid="1336" />
                    <RANKING order="9" place="9" resultid="1933" />
                    <RANKING order="10" place="-1" resultid="2032" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2081" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2082" daytime="10:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2083" daytime="10:10" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1073" daytime="10:16" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1074" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1224" />
                    <RANKING order="2" place="2" resultid="1453" />
                    <RANKING order="3" place="3" resultid="1986" />
                    <RANKING order="4" place="4" resultid="1443" />
                    <RANKING order="5" place="5" resultid="1615" />
                    <RANKING order="6" place="6" resultid="1923" />
                    <RANKING order="7" place="7" resultid="1418" />
                    <RANKING order="8" place="-1" resultid="1467" />
                    <RANKING order="9" place="-1" resultid="1404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1075" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1326" />
                    <RANKING order="2" place="2" resultid="1286" />
                    <RANKING order="3" place="3" resultid="1903" />
                    <RANKING order="4" place="4" resultid="1351" />
                    <RANKING order="5" place="5" resultid="1356" />
                    <RANKING order="6" place="6" resultid="1496" />
                    <RANKING order="7" place="7" resultid="1311" />
                    <RANKING order="8" place="8" resultid="1862" />
                    <RANKING order="9" place="9" resultid="1928" />
                    <RANKING order="10" place="-1" resultid="1996" />
                    <RANKING order="11" place="-1" resultid="1321" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2084" daytime="10:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2085" daytime="10:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2086" daytime="10:26" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1076" daytime="10:30" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1077" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1238" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2087" daytime="10:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1078" daytime="10:34" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1079" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1247" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2088" daytime="10:34" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1080" daytime="10:36" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1081" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1684" />
                    <RANKING order="2" place="2" resultid="1673" />
                    <RANKING order="3" place="3" resultid="1639" />
                    <RANKING order="4" place="4" resultid="1177" />
                    <RANKING order="5" place="5" resultid="1703" />
                    <RANKING order="6" place="6" resultid="1698" />
                    <RANKING order="7" place="7" resultid="1634" />
                    <RANKING order="8" place="8" resultid="2064" />
                    <RANKING order="9" place="9" resultid="1649" />
                    <RANKING order="10" place="10" resultid="1795" />
                    <RANKING order="11" place="-1" resultid="1733" />
                    <RANKING order="12" place="-1" resultid="1765" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1082" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1912" />
                    <RANKING order="2" place="2" resultid="1619" />
                    <RANKING order="3" place="3" resultid="2059" />
                    <RANKING order="4" place="4" resultid="1609" />
                    <RANKING order="5" place="5" resultid="1594" />
                    <RANKING order="6" place="6" resultid="1166" />
                    <RANKING order="7" place="7" resultid="1258" />
                    <RANKING order="8" place="8" resultid="1242" />
                    <RANKING order="9" place="9" resultid="2008" />
                    <RANKING order="10" place="10" resultid="1890" />
                    <RANKING order="11" place="11" resultid="1579" />
                    <RANKING order="12" place="12" resultid="1810" />
                    <RANKING order="13" place="13" resultid="2051" />
                    <RANKING order="14" place="14" resultid="1885" />
                    <RANKING order="15" place="-1" resultid="1625" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2089" daytime="10:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2090" daytime="10:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2091" daytime="10:40" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2092" daytime="10:42" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1083" daytime="10:46" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1084" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1629" />
                    <RANKING order="2" place="2" resultid="1760" />
                    <RANKING order="3" place="3" resultid="1679" />
                    <RANKING order="4" place="4" resultid="1267" />
                    <RANKING order="5" place="5" resultid="1718" />
                    <RANKING order="6" place="6" resultid="1775" />
                    <RANKING order="7" place="7" resultid="1800" />
                    <RANKING order="8" place="8" resultid="1740" />
                    <RANKING order="9" place="9" resultid="1755" />
                    <RANKING order="10" place="10" resultid="1853" />
                    <RANKING order="11" place="11" resultid="1780" />
                    <RANKING order="12" place="12" resultid="1791" />
                    <RANKING order="13" place="-1" resultid="1728" />
                    <RANKING order="14" place="-1" resultid="1804" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1085" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1589" />
                    <RANKING order="2" place="2" resultid="1951" />
                    <RANKING order="3" place="3" resultid="1564" />
                    <RANKING order="4" place="4" resultid="2021" />
                    <RANKING order="5" place="5" resultid="1524" />
                    <RANKING order="6" place="6" resultid="1529" />
                    <RANKING order="7" place="7" resultid="1181" />
                    <RANKING order="8" place="8" resultid="2026" />
                    <RANKING order="9" place="9" resultid="1549" />
                    <RANKING order="10" place="10" resultid="1942" />
                    <RANKING order="11" place="11" resultid="2013" />
                    <RANKING order="12" place="12" resultid="1967" />
                    <RANKING order="13" place="13" resultid="1199" />
                    <RANKING order="14" place="14" resultid="1746" />
                    <RANKING order="15" place="15" resultid="1544" />
                    <RANKING order="16" place="-1" resultid="1569" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2093" daytime="10:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2094" daytime="10:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2095" daytime="10:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2096" daytime="10:52" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1086" daytime="10:56" gender="F" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1087" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1379" />
                    <RANKING order="2" place="2" resultid="1937" />
                    <RANKING order="3" place="3" resultid="1216" />
                    <RANKING order="4" place="4" resultid="1428" />
                    <RANKING order="5" place="5" resultid="1826" />
                    <RANKING order="6" place="6" resultid="1490" />
                    <RANKING order="7" place="7" resultid="1273" />
                    <RANKING order="8" place="8" resultid="1917" />
                    <RANKING order="9" place="9" resultid="1253" />
                    <RANKING order="10" place="10" resultid="1193" />
                    <RANKING order="11" place="11" resultid="1437" />
                    <RANKING order="12" place="12" resultid="1978" />
                    <RANKING order="13" place="13" resultid="1174" />
                    <RANKING order="14" place="14" resultid="1540" />
                    <RANKING order="15" place="15" resultid="1604" />
                    <RANKING order="16" place="16" resultid="1866" />
                    <RANKING order="17" place="17" resultid="1190" />
                    <RANKING order="18" place="18" resultid="1960" />
                    <RANKING order="19" place="19" resultid="1842" />
                    <RANKING order="20" place="20" resultid="1834" />
                    <RANKING order="21" place="21" resultid="1413" />
                    <RANKING order="22" place="22" resultid="2069" />
                    <RANKING order="23" place="23" resultid="2000" />
                    <RANKING order="24" place="-1" resultid="1394" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1088" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1461" />
                    <RANKING order="2" place="2" resultid="1399" />
                    <RANKING order="3" place="3" resultid="1300" />
                    <RANKING order="4" place="4" resultid="1346" />
                    <RANKING order="5" place="5" resultid="1599" />
                    <RANKING order="6" place="6" resultid="1932" />
                    <RANKING order="7" place="7" resultid="1388" />
                    <RANKING order="8" place="8" resultid="1771" />
                    <RANKING order="9" place="9" resultid="1228" />
                    <RANKING order="10" place="10" resultid="1263" />
                    <RANKING order="11" place="11" resultid="1188" />
                    <RANKING order="12" place="12" resultid="1816" />
                    <RANKING order="13" place="13" resultid="2031" />
                    <RANKING order="14" place="14" resultid="1448" />
                    <RANKING order="15" place="15" resultid="1161" />
                    <RANKING order="16" place="16" resultid="1895" />
                    <RANKING order="17" place="17" resultid="1500" />
                    <RANKING order="18" place="18" resultid="1202" />
                    <RANKING order="19" place="19" resultid="1235" />
                    <RANKING order="20" place="20" resultid="2043" />
                    <RANKING order="21" place="-1" resultid="1908" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2097" daytime="10:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2098" daytime="10:58" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2099" daytime="11:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2100" daytime="11:04" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2101" daytime="11:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2102" daytime="11:10" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1089" daytime="11:12" gender="M" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1090" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1152" />
                    <RANKING order="2" place="2" resultid="1376" />
                    <RANKING order="3" place="3" resultid="1472" />
                    <RANKING order="4" place="4" resultid="1985" />
                    <RANKING order="5" place="5" resultid="1481" />
                    <RANKING order="6" place="6" resultid="1442" />
                    <RANKING order="7" place="7" resultid="1922" />
                    <RANKING order="8" place="8" resultid="1614" />
                    <RANKING order="9" place="9" resultid="1973" />
                    <RANKING order="10" place="10" resultid="1848" />
                    <RANKING order="11" place="11" resultid="1433" />
                    <RANKING order="12" place="12" resultid="1417" />
                    <RANKING order="13" place="13" resultid="1486" />
                    <RANKING order="14" place="14" resultid="1963" />
                    <RANKING order="15" place="15" resultid="1981" />
                    <RANKING order="16" place="16" resultid="2040" />
                    <RANKING order="17" place="17" resultid="1948" />
                    <RANKING order="18" place="18" resultid="1838" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1325" />
                    <RANKING order="2" place="2" resultid="1316" />
                    <RANKING order="3" place="3" resultid="1232" />
                    <RANKING order="4" place="3" resultid="1902" />
                    <RANKING order="5" place="5" resultid="1331" />
                    <RANKING order="6" place="6" resultid="1291" />
                    <RANKING order="7" place="7" resultid="1296" />
                    <RANKING order="8" place="8" resultid="1310" />
                    <RANKING order="9" place="9" resultid="1350" />
                    <RANKING order="10" place="10" resultid="1220" />
                    <RANKING order="11" place="11" resultid="1196" />
                    <RANKING order="12" place="12" resultid="1476" />
                    <RANKING order="13" place="13" resultid="1371" />
                    <RANKING order="14" place="14" resultid="2055" />
                    <RANKING order="15" place="15" resultid="1408" />
                    <RANKING order="16" place="16" resultid="2018" />
                    <RANKING order="17" place="17" resultid="1956" />
                    <RANKING order="18" place="18" resultid="1208" />
                    <RANKING order="19" place="19" resultid="1277" />
                    <RANKING order="20" place="20" resultid="1211" />
                    <RANKING order="21" place="21" resultid="2046" />
                    <RANKING order="22" place="22" resultid="1457" />
                    <RANKING order="23" place="-1" resultid="1320" />
                    <RANKING order="24" place="-1" resultid="1366" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2103" daytime="11:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2104" daytime="11:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2105" daytime="11:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2106" daytime="11:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2107" daytime="11:24" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="2108" daytime="11:26" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1092" daytime="11:30" gender="F" number="13" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1093" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1871" />
                    <RANKING order="2" place="2" resultid="1880" />
                    <RANKING order="3" place="3" resultid="1658" />
                    <RANKING order="4" place="4" resultid="1683" />
                    <RANKING order="5" place="5" resultid="1750" />
                    <RANKING order="6" place="6" resultid="1693" />
                    <RANKING order="7" place="-1" resultid="1723" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1094" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1514" />
                    <RANKING order="2" place="2" resultid="1574" />
                    <RANKING order="3" place="3" resultid="1708" />
                    <RANKING order="4" place="4" resultid="1519" />
                    <RANKING order="5" place="5" resultid="2003" />
                    <RANKING order="6" place="6" resultid="1257" />
                    <RANKING order="7" place="7" resultid="1156" />
                    <RANKING order="8" place="8" resultid="1165" />
                    <RANKING order="9" place="9" resultid="1663" />
                    <RANKING order="10" place="10" resultid="1876" />
                    <RANKING order="11" place="11" resultid="1554" />
                    <RANKING order="12" place="12" resultid="2050" />
                    <RANKING order="13" place="13" resultid="1889" />
                    <RANKING order="14" place="14" resultid="1809" />
                    <RANKING order="15" place="-1" resultid="1624" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2109" daytime="11:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2110" daytime="11:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2111" daytime="11:34" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1095" daytime="11:36" gender="M" number="14" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1096" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1644" />
                    <RANKING order="2" place="2" resultid="1990" />
                    <RANKING order="3" place="3" resultid="1280" />
                    <RANKING order="4" place="4" resultid="1688" />
                    <RANKING order="5" place="5" resultid="1266" />
                    <RANKING order="6" place="6" resultid="1678" />
                    <RANKING order="7" place="7" resultid="1790" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1097" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1504" />
                    <RANKING order="2" place="2" resultid="1534" />
                    <RANKING order="3" place="3" resultid="1584" />
                    <RANKING order="4" place="4" resultid="1713" />
                    <RANKING order="5" place="5" resultid="1745" />
                    <RANKING order="6" place="-1" resultid="1653" />
                    <RANKING order="7" place="-1" resultid="1668" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2112" daytime="11:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2113" daytime="11:38" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1098" daytime="11:42" gender="F" number="15" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1099" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1383" />
                    <RANKING order="2" place="2" resultid="1785" />
                    <RANKING order="3" place="3" resultid="1378" />
                    <RANKING order="4" place="4" resultid="1422" />
                    <RANKING order="5" place="5" resultid="1845" />
                    <RANKING order="6" place="6" resultid="1427" />
                    <RANKING order="7" place="7" resultid="1559" />
                    <RANKING order="8" place="8" resultid="1215" />
                    <RANKING order="9" place="9" resultid="1272" />
                    <RANKING order="10" place="10" resultid="1173" />
                    <RANKING order="11" place="11" resultid="1509" />
                    <RANKING order="12" place="12" resultid="1977" />
                    <RANKING order="13" place="13" resultid="1539" />
                    <RANKING order="14" place="14" resultid="1412" />
                    <RANKING order="15" place="-1" resultid="1252" />
                    <RANKING order="16" place="-1" resultid="1393" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1100" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1345" />
                    <RANKING order="2" place="2" resultid="1305" />
                    <RANKING order="3" place="3" resultid="1340" />
                    <RANKING order="4" place="4" resultid="1398" />
                    <RANKING order="5" place="5" resultid="1335" />
                    <RANKING order="6" place="6" resultid="1227" />
                    <RANKING order="7" place="7" resultid="1360" />
                    <RANKING order="8" place="8" resultid="1907" />
                    <RANKING order="9" place="9" resultid="1770" />
                    <RANKING order="10" place="10" resultid="1262" />
                    <RANKING order="11" place="11" resultid="1187" />
                    <RANKING order="12" place="12" resultid="1815" />
                    <RANKING order="13" place="13" resultid="1737" />
                    <RANKING order="14" place="14" resultid="1894" />
                    <RANKING order="15" place="15" resultid="1447" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2114" daytime="11:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2115" daytime="11:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2116" daytime="11:46" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2117" daytime="11:48" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1101" daytime="11:50" gender="M" number="16" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1102" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1151" />
                    <RANKING order="2" place="2" resultid="1223" />
                    <RANKING order="3" place="3" resultid="1466" />
                    <RANKING order="4" place="4" resultid="1375" />
                    <RANKING order="5" place="5" resultid="1471" />
                    <RANKING order="6" place="6" resultid="1403" />
                    <RANKING order="7" place="7" resultid="1452" />
                    <RANKING order="8" place="8" resultid="1480" />
                    <RANKING order="9" place="9" resultid="1485" />
                    <RANKING order="10" place="10" resultid="1432" />
                    <RANKING order="11" place="11" resultid="1972" />
                    <RANKING order="12" place="12" resultid="1947" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1103" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1285" />
                    <RANKING order="2" place="2" resultid="1355" />
                    <RANKING order="3" place="3" resultid="1231" />
                    <RANKING order="4" place="4" resultid="1315" />
                    <RANKING order="5" place="5" resultid="1330" />
                    <RANKING order="6" place="6" resultid="1495" />
                    <RANKING order="7" place="7" resultid="1219" />
                    <RANKING order="8" place="8" resultid="1290" />
                    <RANKING order="9" place="9" resultid="1295" />
                    <RANKING order="10" place="10" resultid="1861" />
                    <RANKING order="11" place="11" resultid="1927" />
                    <RANKING order="12" place="12" resultid="1370" />
                    <RANKING order="13" place="13" resultid="1276" />
                    <RANKING order="14" place="-1" resultid="1995" />
                    <RANKING order="15" place="-1" resultid="1365" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2118" daytime="11:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2119" daytime="11:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2120" daytime="11:54" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2121" daytime="11:56" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-04-06" daytime="15:40" endtime="19:00" number="2" officialmeeting="15:00" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1107" daytime="15:40" gender="F" number="17" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1108" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1240" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2126" daytime="15:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1109" daytime="15:42" gender="M" number="18" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1110" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1249" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2127" daytime="15:42" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1111" daytime="15:44" gender="F" number="19" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1112" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1874" />
                    <RANKING order="2" place="2" resultid="1661" />
                    <RANKING order="3" place="3" resultid="1883" />
                    <RANKING order="4" place="4" resultid="1686" />
                    <RANKING order="5" place="5" resultid="1642" />
                    <RANKING order="6" place="6" resultid="1753" />
                    <RANKING order="7" place="7" resultid="1701" />
                    <RANKING order="8" place="8" resultid="1696" />
                    <RANKING order="9" place="9" resultid="1637" />
                    <RANKING order="10" place="10" resultid="1726" />
                    <RANKING order="11" place="11" resultid="1676" />
                    <RANKING order="12" place="12" resultid="1798" />
                    <RANKING order="13" place="-1" resultid="1706" />
                    <RANKING order="14" place="-1" resultid="1768" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1915" />
                    <RANKING order="2" place="2" resultid="1517" />
                    <RANKING order="3" place="3" resultid="2006" />
                    <RANKING order="4" place="4" resultid="1577" />
                    <RANKING order="5" place="5" resultid="1612" />
                    <RANKING order="6" place="6" resultid="1522" />
                    <RANKING order="7" place="7" resultid="1711" />
                    <RANKING order="8" place="8" resultid="1597" />
                    <RANKING order="9" place="9" resultid="1622" />
                    <RANKING order="10" place="10" resultid="1666" />
                    <RANKING order="11" place="11" resultid="1260" />
                    <RANKING order="12" place="12" resultid="1878" />
                    <RANKING order="13" place="13" resultid="1887" />
                    <RANKING order="14" place="14" resultid="1557" />
                    <RANKING order="15" place="15" resultid="2053" />
                    <RANKING order="16" place="-1" resultid="1582" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2128" daytime="15:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2129" daytime="15:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2130" daytime="15:52" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2131" daytime="15:56" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1114" daytime="16:00" gender="M" number="20" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1115" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1647" />
                    <RANKING order="2" place="2" resultid="1993" />
                    <RANKING order="3" place="3" resultid="1632" />
                    <RANKING order="4" place="4" resultid="1691" />
                    <RANKING order="5" place="5" resultid="1681" />
                    <RANKING order="6" place="6" resultid="1763" />
                    <RANKING order="7" place="7" resultid="1721" />
                    <RANKING order="8" place="8" resultid="1778" />
                    <RANKING order="9" place="9" resultid="1758" />
                    <RANKING order="10" place="10" resultid="1793" />
                    <RANKING order="11" place="-1" resultid="1731" />
                    <RANKING order="12" place="-1" resultid="1807" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1507" />
                    <RANKING order="2" place="2" resultid="1537" />
                    <RANKING order="3" place="3" resultid="1171" />
                    <RANKING order="4" place="4" resultid="1592" />
                    <RANKING order="5" place="5" resultid="1184" />
                    <RANKING order="6" place="6" resultid="1527" />
                    <RANKING order="7" place="7" resultid="1567" />
                    <RANKING order="8" place="8" resultid="1716" />
                    <RANKING order="9" place="9" resultid="2024" />
                    <RANKING order="10" place="10" resultid="1532" />
                    <RANKING order="11" place="11" resultid="1945" />
                    <RANKING order="12" place="12" resultid="1587" />
                    <RANKING order="13" place="13" resultid="2016" />
                    <RANKING order="14" place="14" resultid="1552" />
                    <RANKING order="15" place="15" resultid="1748" />
                    <RANKING order="16" place="-1" resultid="1547" />
                    <RANKING order="17" place="-1" resultid="1572" />
                    <RANKING order="18" place="-1" resultid="1656" />
                    <RANKING order="19" place="-1" resultid="1671" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2132" daytime="16:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2133" daytime="16:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2134" daytime="16:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2135" daytime="16:10" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1104" daytime="16:14" gender="F" number="21" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1105" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1939" />
                    <RANKING order="2" place="2" resultid="1828" />
                    <RANKING order="3" place="3" resultid="1787" />
                    <RANKING order="4" place="4" resultid="1380" />
                    <RANKING order="5" place="5" resultid="1385" />
                    <RANKING order="6" place="6" resultid="1492" />
                    <RANKING order="7" place="7" resultid="1429" />
                    <RANKING order="8" place="8" resultid="1424" />
                    <RANKING order="9" place="9" resultid="1511" />
                    <RANKING order="10" place="10" resultid="1439" />
                    <RANKING order="11" place="11" resultid="1561" />
                    <RANKING order="12" place="12" resultid="1606" />
                    <RANKING order="13" place="13" resultid="1541" />
                    <RANKING order="14" place="14" resultid="1414" />
                    <RANKING order="15" place="-1" resultid="1898" />
                    <RANKING order="16" place="-1" resultid="1395" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1463" />
                    <RANKING order="2" place="2" resultid="1307" />
                    <RANKING order="3" place="3" resultid="1302" />
                    <RANKING order="4" place="4" resultid="1400" />
                    <RANKING order="5" place="5" resultid="1342" />
                    <RANKING order="6" place="6" resultid="1347" />
                    <RANKING order="7" place="7" resultid="1362" />
                    <RANKING order="8" place="8" resultid="1390" />
                    <RANKING order="9" place="9" resultid="1772" />
                    <RANKING order="10" place="10" resultid="1934" />
                    <RANKING order="11" place="11" resultid="1229" />
                    <RANKING order="12" place="12" resultid="1337" />
                    <RANKING order="13" place="13" resultid="1449" />
                    <RANKING order="14" place="14" resultid="1162" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2122" daytime="16:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2123" daytime="16:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2124" daytime="16:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2125" daytime="16:38" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2176" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1117" daytime="16:48" gender="M" number="22" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1118" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1154" />
                    <RANKING order="2" place="2" resultid="1988" />
                    <RANKING order="3" place="3" resultid="1474" />
                    <RANKING order="4" place="4" resultid="1445" />
                    <RANKING order="5" place="5" resultid="1483" />
                    <RANKING order="6" place="6" resultid="1617" />
                    <RANKING order="7" place="7" resultid="1469" />
                    <RANKING order="8" place="8" resultid="1455" />
                    <RANKING order="9" place="9" resultid="1435" />
                    <RANKING order="10" place="10" resultid="1406" />
                    <RANKING order="11" place="11" resultid="1488" />
                    <RANKING order="12" place="12" resultid="1420" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1119" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1328" />
                    <RANKING order="2" place="2" resultid="1288" />
                    <RANKING order="3" place="3" resultid="1905" />
                    <RANKING order="4" place="4" resultid="1333" />
                    <RANKING order="5" place="5" resultid="1318" />
                    <RANKING order="6" place="6" resultid="1298" />
                    <RANKING order="7" place="7" resultid="1293" />
                    <RANKING order="8" place="8" resultid="1368" />
                    <RANKING order="9" place="9" resultid="1313" />
                    <RANKING order="10" place="10" resultid="1358" />
                    <RANKING order="11" place="11" resultid="1221" />
                    <RANKING order="12" place="12" resultid="1998" />
                    <RANKING order="13" place="13" resultid="1373" />
                    <RANKING order="14" place="-1" resultid="1498" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2136" daytime="16:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2137" daytime="16:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2138" daytime="17:02" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2139" daytime="17:10" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1120" daytime="17:18" gender="F" number="23" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1121" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1239" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2140" daytime="17:18" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1122" daytime="17:20" gender="M" number="24" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1123" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1248" />
                    <RANKING order="2" place="2" resultid="1823" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2141" daytime="17:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1124" daytime="17:22" gender="F" number="25" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1125" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1873" />
                    <RANKING order="2" place="2" resultid="1641" />
                    <RANKING order="3" place="3" resultid="1660" />
                    <RANKING order="4" place="4" resultid="1179" />
                    <RANKING order="5" place="5" resultid="1725" />
                    <RANKING order="6" place="6" resultid="1206" />
                    <RANKING order="7" place="7" resultid="2067" />
                    <RANKING order="8" place="8" resultid="1636" />
                    <RANKING order="9" place="9" resultid="1695" />
                    <RANKING order="10" place="10" resultid="1651" />
                    <RANKING order="11" place="11" resultid="1675" />
                    <RANKING order="12" place="12" resultid="1797" />
                    <RANKING order="13" place="-1" resultid="1735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1126" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2005" />
                    <RANKING order="2" place="2" resultid="1159" />
                    <RANKING order="3" place="3" resultid="1665" />
                    <RANKING order="4" place="4" resultid="2062" />
                    <RANKING order="5" place="5" resultid="2011" />
                    <RANKING order="6" place="6" resultid="1611" />
                    <RANKING order="7" place="7" resultid="1621" />
                    <RANKING order="8" place="8" resultid="1521" />
                    <RANKING order="9" place="9" resultid="1168" />
                    <RANKING order="10" place="10" resultid="1858" />
                    <RANKING order="11" place="11" resultid="1245" />
                    <RANKING order="12" place="12" resultid="1892" />
                    <RANKING order="13" place="13" resultid="1812" />
                    <RANKING order="14" place="14" resultid="1877" />
                    <RANKING order="15" place="15" resultid="1819" />
                    <RANKING order="16" place="-1" resultid="1581" />
                    <RANKING order="17" place="-1" resultid="1627" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2142" daytime="17:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2143" daytime="17:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2144" daytime="17:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2145" daytime="17:30" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1127" daytime="17:34" gender="M" number="26" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1128" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1282" />
                    <RANKING order="2" place="2" resultid="1680" />
                    <RANKING order="3" place="3" resultid="1690" />
                    <RANKING order="4" place="4" resultid="1269" />
                    <RANKING order="5" place="5" resultid="1743" />
                    <RANKING order="6" place="6" resultid="1855" />
                    <RANKING order="7" place="7" resultid="1832" />
                    <RANKING order="8" place="8" resultid="1757" />
                    <RANKING order="9" place="9" resultid="1762" />
                    <RANKING order="10" place="10" resultid="1783" />
                    <RANKING order="11" place="11" resultid="1802" />
                    <RANKING order="12" place="12" resultid="1720" />
                    <RANKING order="13" place="13" resultid="1792" />
                    <RANKING order="14" place="-1" resultid="1730" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1129" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1506" />
                    <RANKING order="2" place="2" resultid="1715" />
                    <RANKING order="3" place="3" resultid="1954" />
                    <RANKING order="4" place="4" resultid="2029" />
                    <RANKING order="5" place="5" resultid="1970" />
                    <RANKING order="6" place="6" resultid="2038" />
                    <RANKING order="7" place="-1" resultid="1655" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2146" daytime="17:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2147" daytime="17:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2148" daytime="17:40" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1130" daytime="17:42" gender="F" number="27" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1131" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1381" />
                    <RANKING order="2" place="2" resultid="1430" />
                    <RANKING order="3" place="3" resultid="1425" />
                    <RANKING order="4" place="4" resultid="1217" />
                    <RANKING order="5" place="4" resultid="1940" />
                    <RANKING order="6" place="6" resultid="1920" />
                    <RANKING order="7" place="7" resultid="1440" />
                    <RANKING order="8" place="8" resultid="1512" />
                    <RANKING order="9" place="9" resultid="1255" />
                    <RANKING order="10" place="10" resultid="1194" />
                    <RANKING order="11" place="11" resultid="1979" />
                    <RANKING order="12" place="12" resultid="1843" />
                    <RANKING order="13" place="13" resultid="1836" />
                    <RANKING order="14" place="14" resultid="2071" />
                    <RANKING order="15" place="-1" resultid="1821" />
                    <RANKING order="16" place="-1" resultid="1899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1132" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1464" />
                    <RANKING order="2" place="2" resultid="1303" />
                    <RANKING order="3" place="3" resultid="1401" />
                    <RANKING order="4" place="4" resultid="1308" />
                    <RANKING order="5" place="5" resultid="1602" />
                    <RANKING order="6" place="6" resultid="1391" />
                    <RANKING order="7" place="7" resultid="1935" />
                    <RANKING order="8" place="8" resultid="1910" />
                    <RANKING order="9" place="9" resultid="2034" />
                    <RANKING order="10" place="10" resultid="1163" />
                    <RANKING order="11" place="11" resultid="1502" />
                    <RANKING order="12" place="12" resultid="1236" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2149" daytime="17:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2150" daytime="17:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2151" daytime="17:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2152" daytime="17:52" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1133" daytime="17:56" gender="M" number="28" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1134" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1153" />
                    <RANKING order="2" place="2" resultid="1473" />
                    <RANKING order="3" place="3" resultid="1616" />
                    <RANKING order="4" place="4" resultid="1925" />
                    <RANKING order="5" place="5" resultid="1482" />
                    <RANKING order="6" place="6" resultid="1975" />
                    <RANKING order="7" place="7" resultid="1487" />
                    <RANKING order="8" place="8" resultid="1419" />
                    <RANKING order="9" place="9" resultid="1850" />
                    <RANKING order="10" place="10" resultid="1965" />
                    <RANKING order="11" place="11" resultid="1949" />
                    <RANKING order="12" place="-1" resultid="1983" />
                    <RANKING order="13" place="-1" resultid="1840" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1287" />
                    <RANKING order="2" place="2" resultid="1864" />
                    <RANKING order="3" place="3" resultid="1317" />
                    <RANKING order="4" place="4" resultid="1332" />
                    <RANKING order="5" place="5" resultid="1292" />
                    <RANKING order="6" place="6" resultid="1312" />
                    <RANKING order="7" place="7" resultid="1353" />
                    <RANKING order="8" place="8" resultid="1297" />
                    <RANKING order="9" place="9" resultid="1930" />
                    <RANKING order="10" place="10" resultid="1197" />
                    <RANKING order="11" place="11" resultid="1478" />
                    <RANKING order="12" place="12" resultid="2019" />
                    <RANKING order="13" place="13" resultid="1372" />
                    <RANKING order="14" place="14" resultid="2057" />
                    <RANKING order="15" place="15" resultid="1410" />
                    <RANKING order="16" place="16" resultid="2048" />
                    <RANKING order="17" place="17" resultid="1209" />
                    <RANKING order="18" place="18" resultid="1958" />
                    <RANKING order="19" place="19" resultid="1459" />
                    <RANKING order="20" place="-1" resultid="1278" />
                    <RANKING order="21" place="-1" resultid="1323" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2153" daytime="17:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2154" daytime="18:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2155" daytime="18:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2156" daytime="18:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2157" daytime="18:12" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1136" daytime="18:14" gender="F" number="29" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1137" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1882" />
                    <RANKING order="2" place="2" resultid="1700" />
                    <RANKING order="3" place="3" resultid="1685" />
                    <RANKING order="4" place="4" resultid="1752" />
                    <RANKING order="5" place="5" resultid="1178" />
                    <RANKING order="6" place="6" resultid="1205" />
                    <RANKING order="7" place="7" resultid="2066" />
                    <RANKING order="8" place="8" resultid="1650" />
                    <RANKING order="9" place="-1" resultid="1705" />
                    <RANKING order="10" place="-1" resultid="1734" />
                    <RANKING order="11" place="-1" resultid="1767" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1914" />
                    <RANKING order="2" place="2" resultid="1516" />
                    <RANKING order="3" place="3" resultid="1158" />
                    <RANKING order="4" place="4" resultid="1710" />
                    <RANKING order="5" place="5" resultid="2010" />
                    <RANKING order="6" place="6" resultid="1576" />
                    <RANKING order="7" place="7" resultid="2061" />
                    <RANKING order="8" place="8" resultid="1167" />
                    <RANKING order="9" place="9" resultid="1596" />
                    <RANKING order="10" place="10" resultid="1556" />
                    <RANKING order="11" place="11" resultid="1259" />
                    <RANKING order="12" place="12" resultid="1857" />
                    <RANKING order="13" place="13" resultid="1886" />
                    <RANKING order="14" place="14" resultid="2052" />
                    <RANKING order="15" place="15" resultid="1244" />
                    <RANKING order="16" place="16" resultid="1891" />
                    <RANKING order="17" place="17" resultid="1811" />
                    <RANKING order="18" place="18" resultid="1818" />
                    <RANKING order="19" place="-1" resultid="1626" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2158" daytime="18:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2159" daytime="18:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2160" daytime="18:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2161" daytime="18:20" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1139" daytime="18:24" gender="M" number="30" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1140" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1646" />
                    <RANKING order="2" place="2" resultid="1992" />
                    <RANKING order="3" place="3" resultid="1281" />
                    <RANKING order="4" place="4" resultid="1268" />
                    <RANKING order="5" place="5" resultid="1631" />
                    <RANKING order="6" place="6" resultid="1831" />
                    <RANKING order="7" place="7" resultid="1742" />
                    <RANKING order="8" place="8" resultid="1854" />
                    <RANKING order="9" place="9" resultid="1801" />
                    <RANKING order="10" place="10" resultid="1777" />
                    <RANKING order="11" place="11" resultid="1782" />
                    <RANKING order="12" place="-1" resultid="1806" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1141" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1591" />
                    <RANKING order="2" place="2" resultid="1536" />
                    <RANKING order="3" place="3" resultid="1170" />
                    <RANKING order="4" place="4" resultid="1953" />
                    <RANKING order="5" place="5" resultid="1531" />
                    <RANKING order="6" place="6" resultid="1526" />
                    <RANKING order="7" place="7" resultid="1944" />
                    <RANKING order="8" place="8" resultid="1183" />
                    <RANKING order="9" place="9" resultid="1869" />
                    <RANKING order="10" place="10" resultid="1200" />
                    <RANKING order="11" place="11" resultid="1586" />
                    <RANKING order="12" place="12" resultid="1566" />
                    <RANKING order="13" place="13" resultid="2023" />
                    <RANKING order="14" place="14" resultid="2015" />
                    <RANKING order="15" place="15" resultid="1551" />
                    <RANKING order="16" place="16" resultid="1969" />
                    <RANKING order="17" place="17" resultid="1747" />
                    <RANKING order="18" place="18" resultid="2028" />
                    <RANKING order="19" place="19" resultid="1546" />
                    <RANKING order="20" place="-1" resultid="1571" />
                    <RANKING order="21" place="-1" resultid="1670" />
                    <RANKING order="22" place="-1" resultid="2037" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2162" daytime="18:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2163" daytime="18:26" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2164" daytime="18:28" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2165" daytime="18:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2166" daytime="18:32" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1142" daytime="18:34" gender="F" number="31" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1143" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1788" />
                    <RANKING order="2" place="2" resultid="1386" />
                    <RANKING order="3" place="3" resultid="1274" />
                    <RANKING order="4" place="4" resultid="1175" />
                    <RANKING order="5" place="5" resultid="1493" />
                    <RANKING order="6" place="6" resultid="1829" />
                    <RANKING order="7" place="7" resultid="1542" />
                    <RANKING order="8" place="8" resultid="1846" />
                    <RANKING order="9" place="9" resultid="1919" />
                    <RANKING order="10" place="10" resultid="1415" />
                    <RANKING order="11" place="11" resultid="1254" />
                    <RANKING order="12" place="12" resultid="1961" />
                    <RANKING order="13" place="13" resultid="1562" />
                    <RANKING order="14" place="14" resultid="2001" />
                    <RANKING order="15" place="15" resultid="1191" />
                    <RANKING order="16" place="16" resultid="1867" />
                    <RANKING order="17" place="17" resultid="2070" />
                    <RANKING order="18" place="-1" resultid="1835" />
                    <RANKING order="19" place="-1" resultid="1607" />
                    <RANKING order="20" place="-1" resultid="1396" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1144" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1338" />
                    <RANKING order="2" place="2" resultid="1363" />
                    <RANKING order="3" place="3" resultid="1348" />
                    <RANKING order="4" place="4" resultid="1773" />
                    <RANKING order="5" place="5" resultid="1601" />
                    <RANKING order="6" place="6" resultid="1909" />
                    <RANKING order="7" place="7" resultid="1343" />
                    <RANKING order="8" place="8" resultid="1264" />
                    <RANKING order="9" place="9" resultid="1501" />
                    <RANKING order="10" place="10" resultid="1450" />
                    <RANKING order="11" place="11" resultid="1203" />
                    <RANKING order="12" place="12" resultid="1738" />
                    <RANKING order="13" place="13" resultid="1896" />
                    <RANKING order="14" place="14" resultid="2044" />
                    <RANKING order="15" place="-1" resultid="2033" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2167" daytime="18:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2168" daytime="18:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2169" daytime="18:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2170" daytime="18:40" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="2171" daytime="18:42" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1145" daytime="18:44" gender="M" number="32" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1146" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1454" />
                    <RANKING order="2" place="2" resultid="1405" />
                    <RANKING order="3" place="3" resultid="1444" />
                    <RANKING order="4" place="4" resultid="1987" />
                    <RANKING order="5" place="5" resultid="1468" />
                    <RANKING order="6" place="6" resultid="1974" />
                    <RANKING order="7" place="7" resultid="1982" />
                    <RANKING order="8" place="8" resultid="1924" />
                    <RANKING order="9" place="9" resultid="1434" />
                    <RANKING order="10" place="10" resultid="2041" />
                    <RANKING order="11" place="11" resultid="1849" />
                    <RANKING order="12" place="12" resultid="1839" />
                    <RANKING order="13" place="-1" resultid="1225" />
                    <RANKING order="14" place="-1" resultid="1964" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1147" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1327" />
                    <RANKING order="2" place="2" resultid="1904" />
                    <RANKING order="3" place="3" resultid="1352" />
                    <RANKING order="4" place="4" resultid="1367" />
                    <RANKING order="5" place="5" resultid="1497" />
                    <RANKING order="6" place="6" resultid="1357" />
                    <RANKING order="7" place="7" resultid="1233" />
                    <RANKING order="8" place="8" resultid="1997" />
                    <RANKING order="9" place="9" resultid="1409" />
                    <RANKING order="10" place="10" resultid="1212" />
                    <RANKING order="11" place="11" resultid="1863" />
                    <RANKING order="12" place="12" resultid="1477" />
                    <RANKING order="13" place="13" resultid="1929" />
                    <RANKING order="14" place="14" resultid="1957" />
                    <RANKING order="15" place="15" resultid="1458" />
                    <RANKING order="16" place="16" resultid="2047" />
                    <RANKING order="17" place="-1" resultid="1322" />
                    <RANKING order="18" place="-1" resultid="2056" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="2172" daytime="18:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="2173" daytime="18:48" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="2174" daytime="18:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="2175" daytime="18:52" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="18151" nation="BRA" region="PR" clubid="1270" swrid="95180" name="Clube Uniao Recreativo Palmense" shortname="Clube União">
          <ATHLETES>
            <ATHLETE firstname="Pedro" lastname="Durli Giusti" birthdate="2012-11-06" gender="M" nation="BRA" license="408512" athleteid="1275" externalid="408512">
              <RESULTS>
                <RESULT eventid="1101" points="64" swimtime="00:00:54.32" resultid="1276" heatid="2118" lane="5" />
                <RESULT eventid="1089" points="107" swimtime="00:01:34.21" resultid="1277" heatid="2103" lane="4" />
                <RESULT eventid="1133" status="DSQ" swimtime="00:01:41.37" resultid="1278" heatid="2154" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Langaro Spaniol" birthdate="2013-06-18" gender="F" nation="BRA" license="406600" swrid="5074027" athleteid="1271" externalid="406600">
              <RESULTS>
                <RESULT eventid="1098" points="138" swimtime="00:00:47.12" resultid="1272" heatid="2115" lane="1" />
                <RESULT eventid="1086" points="230" swimtime="00:01:21.96" resultid="1273" heatid="2097" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="264" swimtime="00:00:44.17" resultid="1274" heatid="2169" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Durli Giusti" birthdate="2015-07-05" gender="M" nation="BRA" license="408516" athleteid="1279" externalid="408516">
              <RESULTS>
                <RESULT eventid="1095" points="64" swimtime="00:00:54.37" resultid="1280" heatid="2112" lane="7" />
                <RESULT eventid="1139" points="114" swimtime="00:00:41.49" resultid="1281" heatid="2163" lane="1" />
                <RESULT eventid="1127" points="93" swimtime="00:00:48.74" resultid="1282" heatid="2146" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2864" nation="BRA" region="PR" clubid="1149" swrid="93756" name="Associacao De Pais E Amigos Da Natacao De Ponta Gr" shortname="Apan Ponta Grossa">
          <ATHLETES>
            <ATHLETE firstname="Mariana" lastname="Brunetti Silva" birthdate="2014-03-24" gender="F" nation="BRA" license="390878" swrid="5602517" athleteid="1164" externalid="390878">
              <RESULTS>
                <RESULT eventid="1092" points="82" swimtime="00:00:55.99" resultid="1165" heatid="2110" lane="6" entrytime="00:01:01.91" entrycourse="SCM" />
                <RESULT eventid="1080" points="127" swimtime="00:00:56.41" resultid="1166" heatid="2092" lane="8" entrytime="00:00:59.75" entrycourse="SCM" />
                <RESULT eventid="1136" points="142" swimtime="00:00:43.86" resultid="1167" heatid="2161" lane="1" entrytime="00:00:44.92" entrycourse="SCM" />
                <RESULT eventid="1124" points="110" swimtime="00:00:52.55" resultid="1168" heatid="2144" lane="4" entrytime="00:00:54.69" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Clara Rigailo" birthdate="2013-04-06" gender="F" nation="BRA" license="396828" swrid="5641758" athleteid="1172" externalid="396828">
              <RESULTS>
                <RESULT eventid="1098" points="125" swimtime="00:00:48.68" resultid="1173" heatid="2115" lane="6" />
                <RESULT eventid="1086" points="169" swimtime="00:01:30.75" resultid="1174" heatid="2098" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="231" swimtime="00:00:46.23" resultid="1175" heatid="2171" lane="8" entrytime="00:00:50.28" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Victoria Borges" birthdate="2014-01-16" gender="F" nation="BRA" license="376737" swrid="5602587" athleteid="1155" externalid="376737">
              <RESULTS>
                <RESULT eventid="1092" points="84" swimtime="00:00:55.47" resultid="1156" heatid="2110" lane="5" entrytime="00:00:58.51" entrycourse="SCM" />
                <RESULT eventid="1064" points="127" swimtime="00:03:38.96" resultid="1157" heatid="2072" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.52" />
                    <SPLIT distance="100" swimtime="00:01:44.24" />
                    <SPLIT distance="150" swimtime="00:02:43.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="177" swimtime="00:00:40.82" resultid="1158" heatid="2161" lane="3" entrytime="00:00:40.10" entrycourse="SCM" />
                <RESULT eventid="1124" points="152" swimtime="00:00:47.29" resultid="1159" heatid="2145" lane="3" entrytime="00:00:47.28" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolly" lastname="Victoria Souza" birthdate="2015-11-15" gender="F" nation="BRA" license="400091" swrid="5652902" athleteid="1176" externalid="400091">
              <RESULTS>
                <RESULT eventid="1080" points="111" swimtime="00:00:58.94" resultid="1177" heatid="2089" lane="5" />
                <RESULT eventid="1136" points="107" swimtime="00:00:48.16" resultid="1178" heatid="2158" lane="3" />
                <RESULT eventid="1124" points="83" swimtime="00:00:57.81" resultid="1179" heatid="2143" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Bischof Rogoski" birthdate="2014-10-03" gender="M" nation="BRA" license="401860" swrid="5661341" athleteid="1180" externalid="401860">
              <RESULTS>
                <RESULT eventid="1083" points="86" swimtime="00:00:56.43" resultid="1181" heatid="2096" lane="7" entrytime="00:00:55.51" entrycourse="SCM" />
                <RESULT eventid="1067" points="114" swimtime="00:03:24.90" resultid="1182" heatid="2077" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.42" />
                    <SPLIT distance="100" swimtime="00:01:34.40" />
                    <SPLIT distance="150" swimtime="00:02:29.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="129" swimtime="00:00:39.83" resultid="1183" heatid="2166" lane="1" entrytime="00:00:39.48" entrycourse="SCM" />
                <RESULT eventid="1114" points="110" swimtime="00:01:42.57" resultid="1184" heatid="2132" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Hilgenberg Lievore" birthdate="2014-04-23" gender="M" nation="BRA" license="391167" swrid="5602546" athleteid="1169" externalid="391167">
              <RESULTS>
                <RESULT eventid="1139" points="160" swimtime="00:00:37.11" resultid="1170" heatid="2166" lane="6" entrytime="00:00:38.36" entrycourse="SCM" />
                <RESULT eventid="1114" points="135" swimtime="00:01:35.93" resultid="1171" heatid="2135" lane="5" entrytime="00:01:48.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Campagnoli" birthdate="2013-03-13" gender="M" nation="BRA" license="370651" swrid="5602519" athleteid="1150" externalid="370651">
              <RESULTS>
                <RESULT eventid="1101" points="244" swimtime="00:00:34.80" resultid="1151" heatid="2121" lane="5" entrytime="00:00:35.27" entrycourse="SCM" />
                <RESULT eventid="1089" points="237" swimtime="00:01:12.42" resultid="1152" heatid="2108" lane="6" entrytime="00:01:11.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="201" swimtime="00:01:22.38" resultid="1153" heatid="2154" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="249" swimtime="00:05:37.36" resultid="1154" heatid="2137" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                    <SPLIT distance="100" swimtime="00:01:17.96" />
                    <SPLIT distance="150" swimtime="00:02:02.01" />
                    <SPLIT distance="200" swimtime="00:02:44.14" />
                    <SPLIT distance="250" swimtime="00:03:26.95" />
                    <SPLIT distance="300" swimtime="00:04:09.93" />
                    <SPLIT distance="350" swimtime="00:04:53.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Clara Domingues" birthdate="2012-01-19" gender="F" nation="BRA" license="377291" swrid="5588599" athleteid="1160" externalid="377291">
              <RESULTS>
                <RESULT eventid="1086" points="212" swimtime="00:01:24.23" resultid="1161" heatid="2100" lane="5" entrytime="00:01:32.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="209" swimtime="00:06:29.16" resultid="1162" heatid="2123" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.48" />
                    <SPLIT distance="100" swimtime="00:01:31.08" />
                    <SPLIT distance="150" swimtime="00:02:21.39" />
                    <SPLIT distance="200" swimtime="00:03:11.69" />
                    <SPLIT distance="250" swimtime="00:04:02.22" />
                    <SPLIT distance="300" swimtime="00:04:52.85" />
                    <SPLIT distance="350" swimtime="00:05:42.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="169" swimtime="00:01:39.16" resultid="1163" heatid="2152" lane="8" entrytime="00:01:47.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11303" nation="BRA" region="PR" clubid="1213" swrid="93760" name="Associação De Talentos Da Natação" shortname="Atn/Curitiba">
          <ATHLETES>
            <ATHLETE firstname="Yohanna" lastname="Vitoria Sousa" birthdate="2012-01-20" gender="F" nation="BRA" license="406710" swrid="5717302" athleteid="1234" externalid="406710">
              <RESULTS>
                <RESULT eventid="1086" points="133" swimtime="00:01:38.43" resultid="1235" heatid="2097" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="100" swimtime="00:01:58.01" resultid="1236" heatid="2150" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maximilian" lastname="Hock" birthdate="2016-11-20" gender="M" nation="DEU" license="408352" athleteid="1246" externalid="408352">
              <RESULTS>
                <RESULT eventid="1078" points="37" swimtime="00:01:06.07" resultid="1247" heatid="2088" lane="4" />
                <RESULT eventid="1122" points="57" swimtime="00:00:52.09" resultid="1248" heatid="2141" lane="4" />
                <RESULT eventid="1109" points="49" swimtime="00:01:07.99" resultid="1249" heatid="2127" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Manuela Souza" birthdate="2016-07-07" gender="F" nation="BRA" license="406759" swrid="5717282" athleteid="1237" externalid="406759">
              <RESULTS>
                <RESULT eventid="1076" points="49" swimtime="00:01:08.54" resultid="1238" heatid="2087" lane="4" />
                <RESULT eventid="1120" points="43" swimtime="00:01:05.10" resultid="1239" heatid="2140" lane="4" />
                <RESULT eventid="1107" points="65" swimtime="00:01:10.38" resultid="1240" heatid="2126" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Leal Kuss" birthdate="2012-10-20" gender="M" nation="BRA" license="385085" swrid="5588768" athleteid="1218" externalid="385085">
              <RESULTS>
                <RESULT eventid="1101" points="175" swimtime="00:00:38.87" resultid="1219" heatid="2121" lane="1" entrytime="00:00:39.42" entrycourse="SCM" />
                <RESULT eventid="1089" points="192" swimtime="00:01:17.65" resultid="1220" heatid="2106" lane="3" entrytime="00:01:25.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="197" swimtime="00:06:04.69" resultid="1221" heatid="2137" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Guedes Braga" birthdate="2013-04-09" gender="F" nation="BRA" license="385009" swrid="5602534" athleteid="1214" externalid="385009">
              <RESULTS>
                <RESULT eventid="1098" points="139" swimtime="00:00:46.97" resultid="1215" heatid="2116" lane="2" entrytime="00:00:47.71" entrycourse="SCM" />
                <RESULT eventid="1086" points="295" swimtime="00:01:15.41" resultid="1216" heatid="2101" lane="5" entrytime="00:01:19.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="196" swimtime="00:01:34.48" resultid="1217" heatid="2150" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Duarte De Almeida" birthdate="2013-12-09" gender="M" nation="BRA" license="385711" swrid="5588666" athleteid="1222" externalid="385711">
              <RESULTS>
                <RESULT eventid="1101" points="204" swimtime="00:00:36.94" resultid="1223" heatid="2121" lane="2" entrytime="00:00:38.20" entrycourse="SCM" />
                <RESULT eventid="1073" points="200" swimtime="00:03:07.25" resultid="1224" heatid="2086" lane="3" entrytime="00:03:14.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.20" />
                    <SPLIT distance="100" swimtime="00:01:32.71" />
                    <SPLIT distance="150" swimtime="00:02:29.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" status="DSQ" swimtime="00:00:44.73" resultid="1225" heatid="2174" lane="4" entrytime="00:00:48.05" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Goncalves Ghion" birthdate="2014-10-15" gender="F" nation="BRA" license="406912" swrid="5717269" athleteid="1241" externalid="406912">
              <RESULTS>
                <RESULT eventid="1080" points="93" swimtime="00:01:02.46" resultid="1242" heatid="2091" lane="6" entrytime="00:01:02.99" entrycourse="SCM" />
                <RESULT eventid="1064" points="91" swimtime="00:04:04.88" resultid="1243" heatid="2073" lane="2" />
                <RESULT eventid="1136" points="92" swimtime="00:00:50.71" resultid="1244" heatid="2160" lane="1" entrytime="00:00:50.77" entrycourse="SCM" />
                <RESULT eventid="1124" points="93" swimtime="00:00:55.64" resultid="1245" heatid="2142" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isis" lastname="De Miranda" birthdate="2012-01-10" gender="F" nation="BRA" license="397278" swrid="5652886" athleteid="1226" externalid="397278">
              <RESULTS>
                <RESULT eventid="1098" points="241" swimtime="00:00:39.13" resultid="1227" heatid="2116" lane="6" entrytime="00:00:45.91" entrycourse="SCM" />
                <RESULT eventid="1086" points="279" swimtime="00:01:16.84" resultid="1228" heatid="2101" lane="1" entrytime="00:01:28.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="275" swimtime="00:05:55.63" resultid="1229" heatid="2125" lane="1" entrytime="00:06:34.72" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                    <SPLIT distance="100" swimtime="00:01:20.90" />
                    <SPLIT distance="150" swimtime="00:02:05.21" />
                    <SPLIT distance="200" swimtime="00:02:50.70" />
                    <SPLIT distance="250" swimtime="00:03:37.34" />
                    <SPLIT distance="300" swimtime="00:04:23.80" />
                    <SPLIT distance="350" swimtime="00:05:10.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Vinicius Zonta" birthdate="2012-11-14" gender="M" nation="BRA" license="399517" swrid="5652903" athleteid="1230" externalid="399517">
              <RESULTS>
                <RESULT eventid="1101" points="209" swimtime="00:00:36.61" resultid="1231" heatid="2119" lane="7" />
                <RESULT eventid="1089" points="283" swimtime="00:01:08.23" resultid="1232" heatid="2104" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="157" swimtime="00:00:46.23" resultid="1233" heatid="2175" lane="8" entrytime="00:00:47.08" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="1007" nation="BRA" region="PR" clubid="1900" swrid="93785" name="Santa Mônica Clube De Campo" shortname="Santa Mônica">
          <ATHLETES>
            <ATHLETE firstname="Joaquim" lastname="Hoffmann Zoschke" birthdate="2015-03-22" gender="M" nation="BRA" license="390917" swrid="5602547" athleteid="1989" externalid="390917">
              <RESULTS>
                <RESULT eventid="1095" points="96" swimtime="00:00:47.46" resultid="1990" heatid="2113" lane="6" entrytime="00:00:46.92" entrycourse="SCM" />
                <RESULT eventid="1067" points="134" swimtime="00:03:13.82" resultid="1991" heatid="2077" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.18" />
                    <SPLIT distance="100" swimtime="00:01:34.53" />
                    <SPLIT distance="150" swimtime="00:02:26.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="133" swimtime="00:00:39.45" resultid="1992" heatid="2165" lane="4" entrytime="00:00:39.88" entrycourse="SCM" />
                <RESULT eventid="1114" points="103" swimtime="00:01:44.83" resultid="1993" heatid="2132" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Prestes Alves Pinto" birthdate="2012-01-19" gender="F" nation="BRA" license="377324" swrid="5588867" athleteid="1931" externalid="377324">
              <RESULTS>
                <RESULT eventid="1086" points="335" swimtime="00:01:12.32" resultid="1932" heatid="2102" lane="3" entrytime="00:01:13.78" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1070" points="249" swimtime="00:03:13.45" resultid="1933" heatid="2081" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.55" />
                    <SPLIT distance="100" swimtime="00:01:32.55" />
                    <SPLIT distance="150" swimtime="00:02:31.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="289" swimtime="00:05:49.49" resultid="1934" heatid="2122" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.82" />
                    <SPLIT distance="100" swimtime="00:01:23.80" />
                    <SPLIT distance="150" swimtime="00:02:08.85" />
                    <SPLIT distance="200" swimtime="00:02:53.61" />
                    <SPLIT distance="250" swimtime="00:03:39.23" />
                    <SPLIT distance="300" swimtime="00:04:25.24" />
                    <SPLIT distance="350" swimtime="00:05:09.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="255" swimtime="00:01:26.46" resultid="1935" heatid="2152" lane="7" entrytime="00:01:30.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Coelho Oliveira" birthdate="2015-03-03" gender="F" nation="BRA" license="406839" swrid="5717252" athleteid="2063" externalid="406839">
              <RESULTS>
                <RESULT eventid="1080" points="63" swimtime="00:01:11.21" resultid="2064" heatid="2091" lane="8" entrytime="00:01:11.91" entrycourse="SCM" />
                <RESULT eventid="1064" points="74" swimtime="00:04:21.75" resultid="2065" heatid="2074" lane="2" />
                <RESULT eventid="1136" points="78" swimtime="00:00:53.44" resultid="2066" heatid="2159" lane="5" entrytime="00:00:55.10" entrycourse="SCM" />
                <RESULT eventid="1124" points="71" swimtime="00:01:00.71" resultid="2067" heatid="2143" lane="4" entrytime="00:01:02.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mathias" lastname="Lopes Batista" birthdate="2012-08-22" gender="M" nation="BRA" license="399740" swrid="5652889" athleteid="2017" externalid="399740">
              <RESULTS>
                <RESULT eventid="1089" points="142" swimtime="00:01:25.88" resultid="2018" heatid="2106" lane="6" entrytime="00:01:27.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="116" swimtime="00:01:39.03" resultid="2019" heatid="2156" lane="3" entrytime="00:01:50.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Celli Schneider" birthdate="2013-02-04" gender="M" nation="BRA" license="377317" swrid="5588588" athleteid="1921" externalid="377317">
              <RESULTS>
                <RESULT eventid="1089" points="156" swimtime="00:01:23.16" resultid="1922" heatid="2106" lane="2" entrytime="00:01:27.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1073" points="140" swimtime="00:03:30.78" resultid="1923" heatid="2085" lane="7" entrytime="00:03:37.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.26" />
                    <SPLIT distance="100" swimtime="00:01:41.94" />
                    <SPLIT distance="150" swimtime="00:02:46.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="96" swimtime="00:00:54.45" resultid="1924" heatid="2172" lane="6" />
                <RESULT eventid="1133" points="131" swimtime="00:01:35.07" resultid="1925" heatid="2155" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tais" lastname="Feltrin Martins" birthdate="2013-01-17" gender="F" nation="BRA" license="406840" swrid="5717262" athleteid="2068" externalid="406840">
              <RESULTS>
                <RESULT eventid="1086" points="78" swimtime="00:01:57.34" resultid="2069" heatid="2097" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="74" swimtime="00:01:07.54" resultid="2070" heatid="2168" lane="8" />
                <RESULT eventid="1130" points="74" swimtime="00:02:10.57" resultid="2071" heatid="2151" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="De Siqueira Machado" birthdate="2012-05-25" gender="F" nation="BRA" license="377312" swrid="5588649" athleteid="1906" externalid="377312">
              <RESULTS>
                <RESULT eventid="1098" points="200" swimtime="00:00:41.65" resultid="1907" heatid="2117" lane="8" entrytime="00:00:40.25" entrycourse="SCM" />
                <RESULT eventid="1086" status="DSQ" swimtime="00:01:14.81" resultid="1908" heatid="2102" lane="6" entrytime="00:01:14.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="251" swimtime="00:00:44.97" resultid="1909" heatid="2169" lane="2" />
                <RESULT eventid="1130" points="238" swimtime="00:01:28.55" resultid="1910" heatid="2152" lane="1" entrytime="00:01:37.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helloisa" lastname="De Bassani" birthdate="2012-09-23" gender="F" nation="BRA" license="403403" swrid="5676296" athleteid="2042" externalid="403403">
              <RESULTS>
                <RESULT eventid="1086" points="108" swimtime="00:01:45.22" resultid="2043" heatid="2098" lane="4" />
                <RESULT eventid="1142" points="86" swimtime="00:01:04.09" resultid="2044" heatid="2168" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauren" lastname="Kurecki" birthdate="2014-03-06" gender="F" nation="BRA" license="377314" swrid="5602549" athleteid="1911" externalid="377314">
              <RESULTS>
                <RESULT eventid="1080" points="218" swimtime="00:00:47.13" resultid="1912" heatid="2092" lane="4" entrytime="00:00:46.45" entrycourse="SCM" />
                <RESULT eventid="1064" points="265" swimtime="00:02:51.72" resultid="1913" heatid="2075" lane="5" entrytime="00:03:10.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.15" />
                    <SPLIT distance="100" swimtime="00:01:19.92" />
                    <SPLIT distance="150" swimtime="00:02:06.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="319" swimtime="00:00:33.54" resultid="1914" heatid="2161" lane="4" entrytime="00:00:34.25" entrycourse="SCM" />
                <RESULT eventid="1111" points="271" swimtime="00:01:27.28" resultid="1915" heatid="2131" lane="4" entrytime="00:01:41.41" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Lucachinski Villatore" birthdate="2013-10-04" gender="M" nation="BRA" license="382248" swrid="5588778" athleteid="1946" externalid="382248">
              <RESULTS>
                <RESULT eventid="1101" points="63" swimtime="00:00:54.56" resultid="1947" heatid="2119" lane="2" entrytime="00:01:07.38" entrycourse="SCM" />
                <RESULT eventid="1089" points="77" swimtime="00:01:44.96" resultid="1948" heatid="2105" lane="2" entrytime="00:01:45.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="75" swimtime="00:01:54.47" resultid="1949" heatid="2154" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Gabriel Broto" birthdate="2014-09-14" gender="M" nation="BRA" license="402171" swrid="5661345" athleteid="2035" externalid="402171">
              <RESULTS>
                <RESULT eventid="1067" points="49" swimtime="00:04:29.93" resultid="2036" heatid="2079" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.63" />
                    <SPLIT distance="100" swimtime="00:02:14.60" />
                    <SPLIT distance="150" swimtime="00:03:25.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" status="DNS" swimtime="00:00:00.00" resultid="2037" heatid="2163" lane="7" />
                <RESULT eventid="1127" points="28" swimtime="00:01:12.33" resultid="2038" heatid="2147" lane="2" entrytime="00:01:11.92" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Prestes" birthdate="2014-01-16" gender="M" nation="BRA" license="382249" swrid="5602574" athleteid="1950" externalid="382249">
              <RESULTS>
                <RESULT eventid="1083" points="117" swimtime="00:00:51.01" resultid="1951" heatid="2096" lane="4" entrytime="00:00:48.48" entrycourse="SCM" />
                <RESULT eventid="1067" points="130" swimtime="00:03:15.67" resultid="1952" heatid="2080" lane="6" entrytime="00:03:22.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.39" />
                    <SPLIT distance="100" swimtime="00:01:30.82" />
                    <SPLIT distance="150" swimtime="00:02:25.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="159" swimtime="00:00:37.16" resultid="1953" heatid="2166" lane="7" entrytime="00:00:39.15" entrycourse="SCM" />
                <RESULT eventid="1127" points="105" swimtime="00:00:46.72" resultid="1954" heatid="2148" lane="3" entrytime="00:00:48.43" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lais" lastname="Manika Broto" birthdate="2013-03-27" gender="F" nation="BRA" license="378054" swrid="5588795" athleteid="1936" externalid="378054">
              <RESULTS>
                <RESULT eventid="1086" points="301" swimtime="00:01:14.98" resultid="1937" heatid="2101" lane="7" entrytime="00:01:24.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1070" points="238" swimtime="00:03:16.37" resultid="1938" heatid="2081" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.06" />
                    <SPLIT distance="100" swimtime="00:01:36.22" />
                    <SPLIT distance="150" swimtime="00:02:35.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="325" swimtime="00:05:36.24" resultid="1939" heatid="2176" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.99" />
                    <SPLIT distance="100" swimtime="00:01:18.60" />
                    <SPLIT distance="150" swimtime="00:02:02.91" />
                    <SPLIT distance="200" swimtime="00:02:46.31" />
                    <SPLIT distance="250" swimtime="00:03:31.42" />
                    <SPLIT distance="300" swimtime="00:04:14.03" />
                    <SPLIT distance="350" swimtime="00:04:57.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="196" swimtime="00:01:34.48" resultid="1940" heatid="2149" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jose" lastname="Vinicius Batistella" birthdate="2012-05-15" gender="M" nation="BRA" license="403785" swrid="5684613" athleteid="2054" externalid="403785">
              <RESULTS>
                <RESULT eventid="1089" points="148" swimtime="00:01:24.66" resultid="2055" heatid="2103" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" status="DNS" swimtime="00:00:00.00" resultid="2056" heatid="2172" lane="8" />
                <RESULT eventid="1133" points="106" swimtime="00:01:42.04" resultid="2057" heatid="2154" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Ryan Rosa" birthdate="2014-01-14" gender="M" nation="BRA" license="400032" swrid="5652898" athleteid="2025" externalid="400032">
              <RESULTS>
                <RESULT eventid="1083" points="79" swimtime="00:00:58.14" resultid="2026" heatid="2095" lane="4" entrytime="00:00:59.34" entrycourse="SCM" />
                <RESULT eventid="1067" points="61" swimtime="00:04:11.44" resultid="2027" heatid="2080" lane="8" entrytime="00:04:23.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.47" />
                    <SPLIT distance="100" swimtime="00:02:01.27" />
                    <SPLIT distance="150" swimtime="00:03:06.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="71" swimtime="00:00:48.67" resultid="2028" heatid="2164" lane="2" entrytime="00:00:50.67" entrycourse="SCM" />
                <RESULT eventid="1127" points="58" swimtime="00:00:56.89" resultid="2029" heatid="2148" lane="1" entrytime="00:01:00.67" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Gouvea" birthdate="2013-04-19" gender="M" nation="BRA" license="387378" swrid="5588729" athleteid="1971" externalid="387378">
              <RESULTS>
                <RESULT eventid="1101" points="85" swimtime="00:00:49.28" resultid="1972" heatid="2119" lane="1" />
                <RESULT eventid="1089" points="152" swimtime="00:01:23.86" resultid="1973" heatid="2105" lane="4" entrytime="00:01:38.86" entrycourse="SCM" />
                <RESULT eventid="1145" points="124" swimtime="00:00:49.94" resultid="1974" heatid="2174" lane="8" entrytime="00:00:58.08" entrycourse="SCM" />
                <RESULT eventid="1133" points="105" swimtime="00:01:42.38" resultid="1975" heatid="2155" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Wenceslau Bitencourt" birthdate="2012-02-11" gender="M" nation="BRA" license="377318" swrid="5602591" athleteid="1926" externalid="377318">
              <RESULTS>
                <RESULT eventid="1101" points="144" swimtime="00:00:41.49" resultid="1927" heatid="2118" lane="4" />
                <RESULT eventid="1073" points="178" swimtime="00:03:14.80" resultid="1928" heatid="2084" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.46" />
                    <SPLIT distance="100" swimtime="00:01:29.37" />
                    <SPLIT distance="150" swimtime="00:02:30.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="110" swimtime="00:00:52.02" resultid="1929" heatid="2173" lane="1" />
                <RESULT eventid="1133" points="148" swimtime="00:01:31.22" resultid="1930" heatid="2156" lane="4" entrytime="00:01:38.08" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Hugo Dos Santos" birthdate="2014-07-25" gender="M" nation="BRA" license="397420" swrid="5641766" athleteid="2012" externalid="397420">
              <RESULTS>
                <RESULT eventid="1083" points="65" swimtime="00:01:02.05" resultid="2013" heatid="2094" lane="4" entrytime="00:01:10.77" entrycourse="SCM" />
                <RESULT eventid="1067" points="105" swimtime="00:03:30.22" resultid="2014" heatid="2077" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.84" />
                    <SPLIT distance="100" swimtime="00:01:37.82" />
                    <SPLIT distance="150" swimtime="00:02:35.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="94" swimtime="00:00:44.21" resultid="2015" heatid="2164" lane="5" entrytime="00:00:44.80" entrycourse="SCM" />
                <RESULT eventid="1114" points="71" swimtime="00:01:58.83" resultid="2016" heatid="2132" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Aparecida Lourenço Alves" birthdate="2013-11-06" gender="F" nation="BRA" license="387374" swrid="5588530" athleteid="1959" externalid="387374">
              <RESULTS>
                <RESULT eventid="1086" points="140" swimtime="00:01:36.64" resultid="1960" heatid="2099" lane="5" entrytime="00:01:43.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="120" swimtime="00:00:57.43" resultid="1961" heatid="2168" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Luiz Cruz" birthdate="2012-10-13" gender="M" nation="BRA" license="393209" swrid="5616447" athleteid="1994" externalid="393209">
              <RESULTS>
                <RESULT eventid="1101" status="DNS" swimtime="00:00:00.00" resultid="1995" heatid="2119" lane="4" entrytime="00:00:45.94" entrycourse="SCM" />
                <RESULT eventid="1073" status="DSQ" swimtime="00:00:00.00" resultid="1996" heatid="2084" lane="6" />
                <RESULT eventid="1145" points="127" swimtime="00:00:49.51" resultid="1997" heatid="2173" lane="6" entrytime="00:01:03.62" entrycourse="SCM" />
                <RESULT eventid="1117" points="169" swimtime="00:06:23.25" resultid="1998" heatid="2137" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="100" swimtime="00:01:25.95" />
                    <SPLIT distance="150" swimtime="00:02:14.99" />
                    <SPLIT distance="200" swimtime="00:03:04.80" />
                    <SPLIT distance="250" swimtime="00:03:54.47" />
                    <SPLIT distance="300" swimtime="00:04:44.15" />
                    <SPLIT distance="350" swimtime="00:05:34.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helenna" lastname="Banzatto Silva" birthdate="2013-07-11" gender="F" nation="BRA" license="393210" swrid="5616439" athleteid="1999" externalid="393210">
              <RESULTS>
                <RESULT eventid="1086" points="58" swimtime="00:02:09.28" resultid="2000" heatid="2098" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="108" swimtime="00:00:59.55" resultid="2001" heatid="2170" lane="8" entrytime="00:01:04.15" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Strapasson" birthdate="2012-03-01" gender="M" nation="BRA" license="371377" swrid="5602585" athleteid="1901" externalid="371377">
              <RESULTS>
                <RESULT eventid="1089" points="283" swimtime="00:01:08.23" resultid="1902" heatid="2108" lane="5" entrytime="00:01:11.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1073" points="234" swimtime="00:02:57.88" resultid="1903" heatid="2084" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.77" />
                    <SPLIT distance="100" swimtime="00:01:29.84" />
                    <SPLIT distance="150" swimtime="00:02:20.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="246" swimtime="00:00:39.81" resultid="1904" heatid="2175" lane="5" entrytime="00:00:41.48" entrycourse="SCM" />
                <RESULT eventid="1117" points="284" swimtime="00:05:22.74" resultid="1905" heatid="2136" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Luiza Rocha Batista" birthdate="2013-11-24" gender="F" nation="BRA" license="387379" swrid="5588784" athleteid="1976" externalid="387379">
              <RESULTS>
                <RESULT eventid="1098" points="107" swimtime="00:00:51.35" resultid="1977" heatid="2115" lane="5" entrytime="00:01:01.35" entrycourse="SCM" />
                <RESULT eventid="1086" points="182" swimtime="00:01:28.56" resultid="1978" heatid="2100" lane="8" entrytime="00:01:42.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="128" swimtime="00:01:48.91" resultid="1979" heatid="2149" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Zanotto De Souza" birthdate="2013-08-24" gender="M" nation="BRA" license="388361" swrid="5588974" athleteid="1984" externalid="388361">
              <RESULTS>
                <RESULT eventid="1089" points="216" swimtime="00:01:14.62" resultid="1985" heatid="2107" lane="5" entrytime="00:01:16.88" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1073" points="171" swimtime="00:03:17.50" resultid="1986" heatid="2085" lane="2" entrytime="00:03:29.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.39" />
                    <SPLIT distance="100" swimtime="00:01:34.60" />
                    <SPLIT distance="150" swimtime="00:02:35.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="129" swimtime="00:00:49.33" resultid="1987" heatid="2172" lane="4" />
                <RESULT eventid="1117" points="221" swimtime="00:05:50.78" resultid="1988" heatid="2137" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:22.04" />
                    <SPLIT distance="150" swimtime="00:02:06.57" />
                    <SPLIT distance="200" swimtime="00:02:51.31" />
                    <SPLIT distance="250" swimtime="00:03:37.66" />
                    <SPLIT distance="300" swimtime="00:04:22.71" />
                    <SPLIT distance="350" swimtime="00:05:07.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Zattar" birthdate="2012-04-19" gender="F" nation="BRA" license="401736" swrid="5661351" athleteid="2030" externalid="401736">
              <RESULTS>
                <RESULT eventid="1086" points="229" swimtime="00:01:22.04" resultid="2031" heatid="2098" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1070" status="DSQ" swimtime="00:03:24.55" resultid="2032" heatid="2081" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.56" />
                    <SPLIT distance="100" swimtime="00:01:39.11" />
                    <SPLIT distance="150" swimtime="00:02:39.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" status="DSQ" swimtime="00:00:49.86" resultid="2033" heatid="2168" lane="3" />
                <RESULT eventid="1130" points="187" swimtime="00:01:35.97" resultid="2034" heatid="2150" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cleverson" lastname="Cardoso" birthdate="2013-07-20" gender="M" nation="BRA" license="387382" swrid="5588577" athleteid="1980" externalid="387382">
              <RESULTS>
                <RESULT eventid="1089" points="111" swimtime="00:01:33.25" resultid="1981" heatid="2105" lane="3" entrytime="00:01:41.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="104" swimtime="00:00:52.92" resultid="1982" heatid="2173" lane="3" entrytime="00:01:02.07" entrycourse="SCM" />
                <RESULT eventid="1133" status="DSQ" swimtime="00:01:48.61" resultid="1983" heatid="2156" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Marini" birthdate="2014-04-09" gender="M" nation="BRA" license="382247" swrid="5684582" athleteid="1941" externalid="382247">
              <RESULTS>
                <RESULT eventid="1083" points="65" swimtime="00:01:01.79" resultid="1942" heatid="2093" lane="4" />
                <RESULT eventid="1067" points="113" swimtime="00:03:25.02" resultid="1943" heatid="2078" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.40" />
                    <SPLIT distance="100" swimtime="00:01:37.11" />
                    <SPLIT distance="150" swimtime="00:02:32.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="130" swimtime="00:00:39.78" resultid="1944" heatid="2165" lane="3" entrytime="00:00:42.17" entrycourse="SCM" />
                <RESULT eventid="1114" points="94" swimtime="00:01:48.02" resultid="1945" heatid="2134" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lis" lastname="Cristini Harmatiuk" birthdate="2014-07-19" gender="F" nation="BRA" license="396830" swrid="5641759" athleteid="2058" externalid="396830">
              <RESULTS>
                <RESULT eventid="1080" points="156" swimtime="00:00:52.59" resultid="2059" heatid="2092" lane="5" entrytime="00:00:52.00" entrycourse="SCM" />
                <RESULT eventid="1064" points="163" swimtime="00:03:21.60" resultid="2060" heatid="2072" lane="4" />
                <RESULT eventid="1136" points="163" swimtime="00:00:41.93" resultid="2061" heatid="2161" lane="2" entrytime="00:00:41.73" entrycourse="SCM" />
                <RESULT eventid="1124" points="142" swimtime="00:00:48.34" resultid="2062" heatid="2145" lane="2" entrytime="00:00:49.22" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Andrade Guarido" birthdate="2014-05-17" gender="M" nation="BRA" license="400031" swrid="5652873" athleteid="2020" externalid="400031">
              <RESULTS>
                <RESULT eventid="1083" points="100" swimtime="00:00:53.59" resultid="2021" heatid="2096" lane="2" entrytime="00:00:55.36" entrycourse="SCM" />
                <RESULT eventid="1067" points="118" swimtime="00:03:22.04" resultid="2022" heatid="2079" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.88" />
                    <SPLIT distance="100" swimtime="00:01:38.66" />
                    <SPLIT distance="150" swimtime="00:02:32.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="112" swimtime="00:00:41.75" resultid="2023" heatid="2165" lane="8" entrytime="00:00:43.55" entrycourse="SCM" />
                <RESULT eventid="1114" points="95" swimtime="00:01:47.65" resultid="2024" heatid="2133" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Rodrigues Bortoluzzi" birthdate="2013-10-07" gender="M" nation="BRA" license="387375" swrid="5652897" athleteid="1962" externalid="387375">
              <RESULTS>
                <RESULT eventid="1089" points="113" swimtime="00:01:32.66" resultid="1963" heatid="2104" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" status="DSQ" swimtime="00:01:02.98" resultid="1964" heatid="2173" lane="7" />
                <RESULT eventid="1133" points="82" swimtime="00:01:50.82" resultid="1965" heatid="2155" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mathias" lastname="Bernardo" birthdate="2014-05-17" gender="M" nation="BRA" license="387376" swrid="5652880" athleteid="1966" externalid="387376">
              <RESULTS>
                <RESULT eventid="1083" points="59" swimtime="00:01:03.75" resultid="1967" heatid="2094" lane="1" />
                <RESULT eventid="1067" points="81" swimtime="00:03:49.47" resultid="1968" heatid="2079" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.73" />
                    <SPLIT distance="100" swimtime="00:01:46.70" />
                    <SPLIT distance="150" swimtime="00:02:49.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="85" swimtime="00:00:45.75" resultid="1969" heatid="2164" lane="6" entrytime="00:00:47.97" entrycourse="SCM" />
                <RESULT eventid="1127" points="55" swimtime="00:00:58.07" resultid="1970" heatid="2147" lane="4" entrytime="00:01:05.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="Cirilo Da Cunha" birthdate="2013-05-26" gender="F" nation="BRA" license="377316" swrid="5588595" athleteid="1916" externalid="377316">
              <RESULTS>
                <RESULT eventid="1086" points="216" swimtime="00:01:23.67" resultid="1917" heatid="2099" lane="4" entrytime="00:01:42.99" entrycourse="SCM" />
                <RESULT eventid="1070" points="207" swimtime="00:03:25.96" resultid="1918" heatid="2082" lane="7" entrytime="00:03:50.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.05" />
                    <SPLIT distance="100" swimtime="00:01:39.06" />
                    <SPLIT distance="150" swimtime="00:02:45.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="131" swimtime="00:00:55.86" resultid="1919" heatid="2168" lane="7" />
                <RESULT eventid="1130" points="180" swimtime="00:01:37.12" resultid="1920" heatid="2150" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Julia Rocha" birthdate="2014-02-10" gender="F" nation="BRA" license="397158" swrid="5641767" athleteid="2002" externalid="397158">
              <RESULTS>
                <RESULT eventid="1092" points="94" swimtime="00:00:53.59" resultid="2003" heatid="2111" lane="7" entrytime="00:00:53.29" entrycourse="SCM" />
                <RESULT eventid="1064" points="165" swimtime="00:03:20.96" resultid="2004" heatid="2075" lane="3" entrytime="00:03:20.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                    <SPLIT distance="100" swimtime="00:01:33.54" />
                    <SPLIT distance="150" swimtime="00:02:28.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="182" swimtime="00:00:44.51" resultid="2005" heatid="2145" lane="5" entrytime="00:00:46.65" entrycourse="SCM" />
                <RESULT eventid="1111" points="156" swimtime="00:01:44.80" resultid="2006" heatid="2129" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Coelho De Oliveira" birthdate="2012-11-11" gender="M" nation="BRA" license="385198" swrid="5588600" athleteid="1955" externalid="385198">
              <RESULTS>
                <RESULT eventid="1089" points="123" swimtime="00:01:29.97" resultid="1956" heatid="2105" lane="6" entrytime="00:01:43.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="92" swimtime="00:00:55.14" resultid="1957" heatid="2172" lane="7" />
                <RESULT eventid="1133" points="70" swimtime="00:01:56.88" resultid="1958" heatid="2156" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Victoria De Medeiros" birthdate="2014-08-14" gender="F" nation="BRA" license="403782" swrid="5684611" athleteid="2049" externalid="403782">
              <RESULTS>
                <RESULT eventid="1092" points="49" swimtime="00:01:06.35" resultid="2050" heatid="2109" lane="5" entrytime="00:01:20.19" entrycourse="SCM" />
                <RESULT eventid="1080" points="66" swimtime="00:01:10.11" resultid="2051" heatid="2090" lane="2" entrytime="00:01:15.69" entrycourse="SCM" />
                <RESULT eventid="1136" points="100" swimtime="00:00:49.31" resultid="2052" heatid="2159" lane="3" entrytime="00:00:55.33" entrycourse="SCM" />
                <RESULT eventid="1111" points="72" swimtime="00:02:15.78" resultid="2053" heatid="2129" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:05.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Camily Moraes" birthdate="2014-07-13" gender="F" nation="BRA" license="397159" swrid="5641755" athleteid="2007" externalid="397159">
              <RESULTS>
                <RESULT eventid="1080" points="90" swimtime="00:01:03.23" resultid="2008" heatid="2089" lane="3" />
                <RESULT eventid="1064" points="121" swimtime="00:03:42.87" resultid="2009" heatid="2074" lane="6" entrytime="00:04:45.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.96" />
                    <SPLIT distance="100" swimtime="00:01:44.54" />
                    <SPLIT distance="150" swimtime="00:02:42.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="169" swimtime="00:00:41.44" resultid="2010" heatid="2160" lane="4" entrytime="00:00:45.29" entrycourse="SCM" />
                <RESULT eventid="1124" points="130" swimtime="00:00:49.78" resultid="2011" heatid="2145" lane="1" entrytime="00:00:52.39" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Fachini Kovalski" birthdate="2012-05-15" gender="M" nation="BRA" license="403404" swrid="5676297" athleteid="2045" externalid="403404">
              <RESULTS>
                <RESULT eventid="1089" points="96" swimtime="00:01:37.88" resultid="2046" heatid="2104" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="67" swimtime="00:01:01.33" resultid="2047" heatid="2172" lane="2" />
                <RESULT eventid="1133" points="85" swimtime="00:01:49.63" resultid="2048" heatid="2154" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Borges Piekarzievicz" birthdate="2013-09-10" gender="M" nation="BRA" license="403142" swrid="5676294" athleteid="2039" externalid="403142">
              <RESULTS>
                <RESULT eventid="1089" points="88" swimtime="00:01:40.73" resultid="2040" heatid="2104" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="77" swimtime="00:00:58.57" resultid="2041" heatid="2172" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13068" nation="BRA" region="PR" clubid="1859" swrid="93787" name="Sociedade Morgenau" shortname="Morgenau">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Luiza Melo" birthdate="2015-02-07" gender="F" nation="BRA" license="406717" swrid="5717280" athleteid="1879" externalid="406717">
              <RESULTS>
                <RESULT eventid="1092" points="87" swimtime="00:00:54.98" resultid="1880" heatid="2110" lane="3" entrytime="00:01:01.54" entrycourse="SCM" />
                <RESULT eventid="1064" points="119" swimtime="00:03:43.84" resultid="1881" heatid="2074" lane="8" />
                <RESULT eventid="1136" points="133" swimtime="00:00:44.83" resultid="1882" heatid="2161" lane="8" entrytime="00:00:44.97" entrycourse="SCM" />
                <RESULT eventid="1111" points="119" swimtime="00:01:54.59" resultid="1883" heatid="2128" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Felipe Kuhn" birthdate="2014-03-22" gender="M" nation="BRA" license="392121" swrid="5602536" athleteid="1868" externalid="392121">
              <RESULTS>
                <RESULT eventid="1139" points="126" swimtime="00:00:40.17" resultid="1869" heatid="2164" lane="4" entrytime="00:00:44.35" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Tomaz Zmievski" birthdate="2012-09-20" gender="F" nation="BRA" license="406725" swrid="5717300" athleteid="1893" externalid="406725">
              <RESULTS>
                <RESULT eventid="1098" points="88" swimtime="00:00:54.70" resultid="1894" heatid="2115" lane="2" />
                <RESULT eventid="1086" points="200" swimtime="00:01:25.90" resultid="1895" heatid="2097" lane="4" />
                <RESULT eventid="1142" points="124" swimtime="00:00:56.75" resultid="1896" heatid="2168" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Lara" birthdate="2014-09-02" gender="F" nation="BRA" license="406686" swrid="5717259" athleteid="1875" externalid="406686">
              <RESULTS>
                <RESULT eventid="1092" points="52" swimtime="00:01:05.04" resultid="1876" heatid="2109" lane="2" />
                <RESULT eventid="1124" points="57" swimtime="00:01:05.39" resultid="1877" heatid="2142" lane="4" />
                <RESULT eventid="1111" points="86" swimtime="00:02:07.88" resultid="1878" heatid="2129" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Fernanda De Lima" birthdate="2013-09-26" gender="F" nation="BRA" license="378290" swrid="5588693" athleteid="1865" externalid="378290">
              <RESULTS>
                <RESULT eventid="1086" points="151" swimtime="00:01:34.30" resultid="1866" heatid="2100" lane="2" entrytime="00:01:35.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="92" swimtime="00:01:02.72" resultid="1867" heatid="2168" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Seiffert Mafra" birthdate="2013-01-11" gender="F" nation="BRA" license="406729" swrid="5717296" athleteid="1897" externalid="406729">
              <RESULTS>
                <RESULT eventid="1104" status="DNS" swimtime="00:00:00.00" resultid="1898" heatid="2124" lane="8" />
                <RESULT eventid="1130" status="DNS" swimtime="00:00:00.00" resultid="1899" heatid="2149" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maryana" lastname="Lemos Carvalho" birthdate="2014-02-10" gender="F" nation="BRA" license="406718" swrid="5717278" athleteid="1884" externalid="406718">
              <RESULTS>
                <RESULT eventid="1080" points="55" swimtime="00:01:14.52" resultid="1885" heatid="2089" lane="4" />
                <RESULT eventid="1136" points="111" swimtime="00:00:47.59" resultid="1886" heatid="2160" lane="2" entrytime="00:00:48.98" entrycourse="SCM" />
                <RESULT eventid="1111" points="84" swimtime="00:02:08.64" resultid="1887" heatid="2130" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Nitz Costa" birthdate="2015-02-09" gender="F" nation="BRA" license="397328" swrid="5641773" athleteid="1870" externalid="397328">
              <RESULTS>
                <RESULT eventid="1092" points="115" swimtime="00:00:50.01" resultid="1871" heatid="2111" lane="5" entrytime="00:00:48.30" entrycourse="SCM" />
                <RESULT eventid="1064" points="156" swimtime="00:03:24.88" resultid="1872" heatid="2073" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.61" />
                    <SPLIT distance="100" swimtime="00:01:36.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="160" swimtime="00:00:46.44" resultid="1873" heatid="2145" lane="4" entrytime="00:00:46.43" entrycourse="SCM" />
                <RESULT eventid="1111" points="145" swimtime="00:01:47.46" resultid="1874" heatid="2131" lane="5" entrytime="00:01:48.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Alves" birthdate="2012-10-12" gender="M" nation="BRA" license="369324" swrid="5588674" athleteid="1860" externalid="369324">
              <RESULTS>
                <RESULT eventid="1101" points="148" swimtime="00:00:41.09" resultid="1861" heatid="2120" lane="7" entrytime="00:00:43.03" entrycourse="SCM" />
                <RESULT eventid="1073" points="184" swimtime="00:03:12.48" resultid="1862" heatid="2085" lane="3" entrytime="00:03:26.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.84" />
                    <SPLIT distance="100" swimtime="00:01:32.80" />
                    <SPLIT distance="150" swimtime="00:02:31.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="111" swimtime="00:00:51.84" resultid="1863" heatid="2172" lane="3" />
                <RESULT eventid="1133" points="219" swimtime="00:01:20.14" resultid="1864" heatid="2157" lane="4" entrytime="00:01:23.65" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cecilia Carstens" birthdate="2014-02-22" gender="F" nation="BRA" license="406721" swrid="5717251" athleteid="1888" externalid="406721">
              <RESULTS>
                <RESULT eventid="1092" points="41" swimtime="00:01:10.67" resultid="1889" heatid="2110" lane="1" entrytime="00:01:07.06" entrycourse="SCM" />
                <RESULT eventid="1080" points="87" swimtime="00:01:03.86" resultid="1890" heatid="2091" lane="4" entrytime="00:01:01.55" entrycourse="SCM" />
                <RESULT eventid="1136" points="82" swimtime="00:00:52.60" resultid="1891" heatid="2159" lane="7" entrytime="00:00:58.38" entrycourse="SCM" />
                <RESULT eventid="1124" points="74" swimtime="00:00:59.98" resultid="1892" heatid="2144" lane="1" entrytime="00:01:01.24" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13038" nation="BRA" region="PR" clubid="1185" swrid="93759" name="Associação De Pais E Atletas De Natação Ws/Crb" shortname="Apan/Ws">
          <ATHLETES>
            <ATHLETE firstname="Julia" lastname="Dos Santos" birthdate="2013-06-26" gender="F" nation="BRA" license="387512" swrid="5588662" athleteid="1192" externalid="387512">
              <RESULTS>
                <RESULT eventid="1086" points="195" swimtime="00:01:26.58" resultid="1193" heatid="2099" lane="2" entrytime="00:01:49.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="148" swimtime="00:01:43.69" resultid="1194" heatid="2151" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leon" lastname="Bernardo Bello" birthdate="2014-11-23" gender="M" nation="BRA" license="400324" swrid="5717246" athleteid="1198" externalid="400324">
              <RESULTS>
                <RESULT eventid="1083" points="57" swimtime="00:01:04.77" resultid="1199" heatid="2093" lane="3" />
                <RESULT eventid="1139" points="119" swimtime="00:00:40.93" resultid="1200" heatid="2165" lane="5" entrytime="00:00:40.80" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Bobko Ganacim" birthdate="2013-08-02" gender="F" nation="BRA" license="397332" swrid="5641754" athleteid="1189" externalid="397332">
              <RESULTS>
                <RESULT eventid="1086" points="149" swimtime="00:01:34.66" resultid="1190" heatid="2099" lane="7" entrytime="00:01:56.18" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="107" swimtime="00:00:59.65" resultid="1191" heatid="2167" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Gramms Dallarosa" birthdate="2015-01-14" gender="F" nation="BRA" license="406868" swrid="5717270" athleteid="1204" externalid="406868">
              <RESULTS>
                <RESULT eventid="1136" points="79" swimtime="00:00:53.37" resultid="1205" heatid="2159" lane="2" entrytime="00:00:56.57" entrycourse="SCM" />
                <RESULT eventid="1124" points="72" swimtime="00:01:00.55" resultid="1206" heatid="2143" lane="5" entrytime="00:01:03.95" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Bernardi Iurk" birthdate="2012-04-14" gender="M" nation="BRA" license="408687" athleteid="1210" externalid="408687">
              <RESULTS>
                <RESULT eventid="1089" points="106" swimtime="00:01:34.59" resultid="1211" heatid="2104" lane="4" />
                <RESULT eventid="1145" points="111" swimtime="00:00:51.80" resultid="1212" heatid="2173" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Bernardi Iurk" birthdate="2012-04-14" gender="M" nation="BRA" license="406940" swrid="5717245" athleteid="1207" externalid="406940">
              <RESULTS>
                <RESULT eventid="1089" points="110" swimtime="00:01:33.56" resultid="1208" heatid="2103" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="84" swimtime="00:01:49.94" resultid="1209" heatid="2155" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.58" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Da Reginalda" birthdate="2012-11-09" gender="M" nation="BRA" license="400275" swrid="5717253" athleteid="1195" externalid="400275">
              <RESULTS>
                <RESULT eventid="1089" points="188" swimtime="00:01:18.22" resultid="1196" heatid="2104" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="138" swimtime="00:01:33.43" resultid="1197" heatid="2153" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Cravcenco Marcondes" birthdate="2012-06-23" gender="F" nation="BRA" license="406866" athleteid="1201" externalid="406866">
              <RESULTS>
                <RESULT eventid="1086" points="155" swimtime="00:01:33.50" resultid="1202" heatid="2098" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="149" swimtime="00:00:53.48" resultid="1203" heatid="2169" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Ferreira" birthdate="2012-12-29" gender="F" nation="BRA" license="382235" swrid="5602538" athleteid="1186" externalid="382235">
              <RESULTS>
                <RESULT eventid="1098" points="154" swimtime="00:00:45.45" resultid="1187" heatid="2116" lane="7" entrytime="00:00:49.33" entrycourse="SCM" />
                <RESULT eventid="1086" points="247" swimtime="00:01:20.08" resultid="1188" heatid="2100" lane="3" entrytime="00:01:33.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="1824" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Theo" lastname="Ribeiro Melo" birthdate="2013-02-25" gender="M" nation="BRA" license="406921" swrid="5717293" athleteid="1847" externalid="406921">
              <RESULTS>
                <RESULT eventid="1089" points="150" swimtime="00:01:24.25" resultid="1848" heatid="2105" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="72" swimtime="00:00:59.90" resultid="1849" heatid="2172" lane="1" />
                <RESULT eventid="1133" points="89" swimtime="00:01:47.90" resultid="1850" heatid="2154" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Schneider Yazbek" birthdate="2013-03-07" gender="F" nation="BRA" license="378329" swrid="5588907" athleteid="1825" externalid="378329">
              <RESULTS>
                <RESULT eventid="1086" points="285" swimtime="00:01:16.29" resultid="1826" heatid="2102" lane="8" entrytime="00:01:17.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1070" points="259" swimtime="00:03:11.08" resultid="1827" heatid="2082" lane="4" entrytime="00:03:21.14" entrycourse="SCM" />
                <RESULT eventid="1104" points="325" swimtime="00:05:36.26" resultid="1828" heatid="2122" lane="5" />
                <RESULT eventid="1142" points="199" swimtime="00:00:48.55" resultid="1829" heatid="2168" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Paes Schemiko" birthdate="2013-02-25" gender="F" nation="BRA" license="406918" athleteid="1844" externalid="406918">
              <RESULTS>
                <RESULT eventid="1098" points="176" swimtime="00:00:43.43" resultid="1845" heatid="2114" lane="2" />
                <RESULT eventid="1142" points="162" swimtime="00:00:51.95" resultid="1846" heatid="2167" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Livia" lastname="Nunes Lingner" birthdate="2013-04-03" gender="F" nation="BRA" license="402280" swrid="5661353" athleteid="1833" externalid="402280">
              <RESULTS>
                <RESULT eventid="1086" points="124" swimtime="00:01:40.70" resultid="1834" heatid="2098" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" status="DSQ" swimtime="00:00:52.50" resultid="1835" heatid="2169" lane="5" />
                <RESULT eventid="1130" points="77" swimtime="00:02:08.78" resultid="1836" heatid="2151" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Henrique Ballatka" birthdate="2013-08-26" gender="M" nation="BRA" license="405839" swrid="5697229" athleteid="1837" externalid="405839">
              <RESULTS>
                <RESULT eventid="1089" points="70" swimtime="00:01:48.64" resultid="1838" heatid="2105" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="33" swimtime="00:01:17.25" resultid="1839" heatid="2173" lane="2" entrytime="00:01:35.13" entrycourse="SCM" />
                <RESULT eventid="1133" status="DSQ" swimtime="00:02:26.35" resultid="1840" heatid="2155" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:10.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Guidin Madureira" birthdate="2015-01-10" gender="M" nation="BRA" license="402116" swrid="5661347" athleteid="1830" externalid="402116">
              <RESULTS>
                <RESULT eventid="1139" points="99" swimtime="00:00:43.45" resultid="1831" heatid="2162" lane="4" />
                <RESULT eventid="1127" points="41" swimtime="00:01:03.68" resultid="1832" heatid="2146" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="De Andrade" birthdate="2015-12-24" gender="M" nation="BRA" license="406922" athleteid="1851" externalid="406922" />
            <ATHLETE firstname="Gabriela" lastname="Borges Duarte" birthdate="2014-02-10" gender="F" nation="BRA" license="408688" athleteid="1856" externalid="408688">
              <RESULTS>
                <RESULT eventid="1136" points="121" swimtime="00:00:46.35" resultid="1857" heatid="2158" lane="4" />
                <RESULT eventid="1124" points="101" swimtime="00:00:54.15" resultid="1858" heatid="2142" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Samuel" lastname="Melo Lima" birthdate="2015-10-30" gender="M" nation="BRA" license="406933" athleteid="1852" externalid="406933">
              <RESULTS>
                <RESULT eventid="1083" points="30" swimtime="00:01:20.27" resultid="1853" heatid="2093" lane="6" />
                <RESULT eventid="1139" points="36" swimtime="00:01:00.93" resultid="1854" heatid="2162" lane="5" />
                <RESULT eventid="1127" points="42" swimtime="00:01:03.49" resultid="1855" heatid="2146" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Zanatta Duda" birthdate="2013-08-28" gender="F" nation="BRA" license="406914" swrid="5717306" athleteid="1841" externalid="406914">
              <RESULTS>
                <RESULT eventid="1086" points="130" swimtime="00:01:39.14" resultid="1842" heatid="2099" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="109" swimtime="00:01:54.70" resultid="1843" heatid="2150" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2539" nation="BRA" region="PR" clubid="1250" swrid="93771" name="Círculo Militar Do Paraná" shortname="Círculo Militar">
          <ATHLETES>
            <ATHLETE firstname="Arya" lastname="Zgoda De Brito Afonso" birthdate="2013-01-03" gender="F" nation="BRA" license="378331" swrid="5588976" athleteid="1251" externalid="378331">
              <RESULTS>
                <RESULT eventid="1098" status="DSQ" swimtime="00:00:53.47" resultid="1252" heatid="2114" lane="1" />
                <RESULT eventid="1086" points="205" swimtime="00:01:25.21" resultid="1253" heatid="2100" lane="4" entrytime="00:01:32.39" entrycourse="SCM" />
                <RESULT eventid="1142" points="127" swimtime="00:00:56.39" resultid="1254" heatid="2170" lane="2" entrytime="00:00:55.39" entrycourse="SCM" />
                <RESULT eventid="1130" points="153" swimtime="00:01:42.48" resultid="1255" heatid="2151" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Cavalcante Pierin" birthdate="2012-10-30" gender="F" nation="BRA" license="406952" swrid="5717250" athleteid="1261" externalid="406952">
              <RESULTS>
                <RESULT eventid="1098" points="162" swimtime="00:00:44.72" resultid="1262" heatid="2114" lane="4" />
                <RESULT eventid="1086" points="277" swimtime="00:01:17.02" resultid="1263" heatid="2098" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="219" swimtime="00:00:47.01" resultid="1264" heatid="2169" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Cavalcante Pierin" birthdate="2015-03-31" gender="M" nation="BRA" license="408082" athleteid="1265" externalid="408082">
              <RESULTS>
                <RESULT eventid="1095" points="43" swimtime="00:01:02.00" resultid="1266" heatid="2112" lane="6" />
                <RESULT eventid="1083" points="67" swimtime="00:01:01.38" resultid="1267" heatid="2094" lane="8" />
                <RESULT eventid="1139" points="104" swimtime="00:00:42.74" resultid="1268" heatid="2162" lane="3" />
                <RESULT eventid="1127" points="68" swimtime="00:00:53.92" resultid="1269" heatid="2146" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Vieira Coelho" birthdate="2014-09-28" gender="F" nation="BRA" license="406951" swrid="5717301" athleteid="1256" externalid="406951">
              <RESULTS>
                <RESULT eventid="1092" points="89" swimtime="00:00:54.59" resultid="1257" heatid="2109" lane="6" />
                <RESULT eventid="1080" points="111" swimtime="00:00:58.86" resultid="1258" heatid="2092" lane="1" entrytime="00:00:58.90" entrycourse="SCM" />
                <RESULT eventid="1136" points="125" swimtime="00:00:45.77" resultid="1259" heatid="2160" lane="7" entrytime="00:00:49.84" entrycourse="SCM" />
                <RESULT eventid="1111" points="118" swimtime="00:01:55.18" resultid="1260" heatid="2129" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="263" nation="BRA" region="PR" clubid="1283" swrid="75436" name="Clube Curitibano" shortname="Curitibano">
          <ATHLETES>
            <ATHLETE firstname="Barbara" lastname="Bittencourt Ribas" birthdate="2013-02-01" gender="F" nation="BRA" license="372682" swrid="5588555" athleteid="1377" externalid="372682">
              <RESULTS>
                <RESULT eventid="1098" points="239" swimtime="00:00:39.28" resultid="1378" heatid="2116" lane="4" entrytime="00:00:40.79" entrycourse="SCM" />
                <RESULT eventid="1086" points="309" swimtime="00:01:14.29" resultid="1379" heatid="2101" lane="3" entrytime="00:01:19.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="302" swimtime="00:05:44.59" resultid="1380" heatid="2123" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                    <SPLIT distance="100" swimtime="00:01:25.48" />
                    <SPLIT distance="150" swimtime="00:02:10.05" />
                    <SPLIT distance="200" swimtime="00:02:54.92" />
                    <SPLIT distance="250" swimtime="00:03:39.81" />
                    <SPLIT distance="300" swimtime="00:04:23.05" />
                    <SPLIT distance="350" swimtime="00:05:05.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="240" swimtime="00:01:28.26" resultid="1381" heatid="2151" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Albuquerque" birthdate="2012-08-17" gender="F" nation="BRA" license="369275" swrid="5602507" athleteid="1334" externalid="369275">
              <RESULTS>
                <RESULT eventid="1098" points="261" swimtime="00:00:38.13" resultid="1335" heatid="2117" lane="2" entrytime="00:00:39.72" entrycourse="SCM" />
                <RESULT eventid="1070" points="273" swimtime="00:03:07.83" resultid="1336" heatid="2083" lane="1" entrytime="00:03:18.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.09" />
                    <SPLIT distance="100" swimtime="00:01:35.26" />
                    <SPLIT distance="150" swimtime="00:02:24.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="252" swimtime="00:06:06.15" resultid="1337" heatid="2124" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.01" />
                    <SPLIT distance="100" swimtime="00:01:26.04" />
                    <SPLIT distance="150" swimtime="00:02:13.01" />
                    <SPLIT distance="200" swimtime="00:03:00.47" />
                    <SPLIT distance="250" swimtime="00:03:47.97" />
                    <SPLIT distance="300" swimtime="00:04:35.20" />
                    <SPLIT distance="350" swimtime="00:05:22.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="391" swimtime="00:00:38.79" resultid="1338" heatid="2171" lane="4" entrytime="00:00:41.62" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="De Lima Cavalcanti" birthdate="2014-10-07" gender="M" nation="BRA" license="385884" swrid="5684550" athleteid="1712" externalid="385884">
              <RESULTS>
                <RESULT eventid="1095" points="48" swimtime="00:00:59.76" resultid="1713" heatid="2113" lane="7" entrytime="00:00:49.23" entrycourse="SCM" />
                <RESULT eventid="1067" points="144" swimtime="00:03:09.19" resultid="1714" heatid="2078" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.23" />
                    <SPLIT distance="100" swimtime="00:01:34.45" />
                    <SPLIT distance="150" swimtime="00:02:23.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="135" swimtime="00:00:43.04" resultid="1715" heatid="2148" lane="5" entrytime="00:00:41.45" entrycourse="SCM" />
                <RESULT eventid="1114" points="96" swimtime="00:01:47.26" resultid="1716" heatid="2134" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcela" lastname="Tallao Benke" birthdate="2014-10-07" gender="F" nation="BRA" license="382075" swrid="5602586" athleteid="1513" externalid="382075">
              <RESULTS>
                <RESULT eventid="1092" points="196" swimtime="00:00:41.92" resultid="1514" heatid="2111" lane="4" entrytime="00:00:40.65" entrycourse="SCM" />
                <RESULT eventid="1064" points="260" swimtime="00:02:52.66" resultid="1515" heatid="2075" lane="4" entrytime="00:03:04.71" entrycourse="SCM" />
                <RESULT eventid="1136" points="234" swimtime="00:00:37.19" resultid="1516" heatid="2161" lane="5" entrytime="00:00:36.93" entrycourse="SCM" />
                <RESULT eventid="1111" points="267" swimtime="00:01:27.67" resultid="1517" heatid="2131" lane="3" entrytime="00:01:52.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Kraemer Geremia" birthdate="2013-08-16" gender="M" nation="BRA" license="377041" swrid="5588762" athleteid="1470" externalid="377041">
              <RESULTS>
                <RESULT eventid="1101" points="152" swimtime="00:00:40.73" resultid="1471" heatid="2120" lane="5" entrytime="00:00:41.30" entrycourse="SCM" />
                <RESULT eventid="1089" points="217" swimtime="00:01:14.51" resultid="1472" heatid="2107" lane="6" entrytime="00:01:17.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="160" swimtime="00:01:28.85" resultid="1473" heatid="2156" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="214" swimtime="00:05:54.45" resultid="1474" heatid="2137" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.93" />
                    <SPLIT distance="100" swimtime="00:01:24.59" />
                    <SPLIT distance="150" swimtime="00:02:10.89" />
                    <SPLIT distance="200" swimtime="00:02:56.29" />
                    <SPLIT distance="250" swimtime="00:03:42.22" />
                    <SPLIT distance="300" swimtime="00:04:27.93" />
                    <SPLIT distance="350" swimtime="00:05:11.78" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Artigas Pinheiro" birthdate="2013-07-31" gender="F" nation="BRA" license="377153" swrid="5588534" athleteid="1508" externalid="377153">
              <RESULTS>
                <RESULT eventid="1098" points="122" swimtime="00:00:49.08" resultid="1509" heatid="2116" lane="1" entrytime="00:00:49.57" entrycourse="SCM" />
                <RESULT eventid="1070" points="177" swimtime="00:03:36.66" resultid="1510" heatid="2082" lane="2" entrytime="00:03:45.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:42.47" />
                    <SPLIT distance="150" swimtime="00:02:51.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="214" swimtime="00:06:26.20" resultid="1511" heatid="2122" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.95" />
                    <SPLIT distance="100" swimtime="00:01:32.00" />
                    <SPLIT distance="150" swimtime="00:02:21.99" />
                    <SPLIT distance="200" swimtime="00:03:12.11" />
                    <SPLIT distance="250" swimtime="00:04:02.04" />
                    <SPLIT distance="300" swimtime="00:04:52.48" />
                    <SPLIT distance="350" swimtime="00:05:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="178" swimtime="00:01:37.52" resultid="1512" heatid="2149" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Stramandinoli Zanicotti" birthdate="2013-06-18" gender="F" nation="BRA" license="376967" swrid="5588924" athleteid="1411" externalid="376967">
              <RESULTS>
                <RESULT eventid="1098" points="57" swimtime="00:01:03.32" resultid="1412" heatid="2115" lane="7" />
                <RESULT eventid="1086" points="102" swimtime="00:01:47.41" resultid="1413" heatid="2099" lane="1" entrytime="00:02:07.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="106" swimtime="00:08:08.51" resultid="1414" heatid="2122" lane="4" />
                <RESULT eventid="1142" points="127" swimtime="00:00:56.34" resultid="1415" heatid="2170" lane="1" entrytime="00:01:03.44" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alan" lastname="Batista Grise" birthdate="2014-03-27" gender="M" nation="BRA" license="391007" swrid="5602513" athleteid="1543" externalid="391007">
              <RESULTS>
                <RESULT eventid="1083" points="55" swimtime="00:01:05.53" resultid="1544" heatid="2095" lane="6" entrytime="00:01:04.24" entrycourse="SCM" />
                <RESULT eventid="1067" points="50" swimtime="00:04:28.58" resultid="1545" heatid="2079" lane="7">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:02:09.63" />
                    <SPLIT distance="150" swimtime="00:03:23.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="24" swimtime="00:01:09.17" resultid="1546" heatid="2164" lane="7" entrytime="00:00:51.24" entrycourse="SCM" />
                <RESULT eventid="1114" status="DSQ" swimtime="00:00:00.00" resultid="1547" heatid="2134" lane="4" entrytime="00:02:28.92" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olavo" lastname="Valduga Artigas" birthdate="2012-06-26" gender="M" nation="BRA" license="369270" swrid="5588941" athleteid="1319" externalid="369270">
              <RESULTS>
                <RESULT eventid="1089" status="DNS" swimtime="00:00:00.00" resultid="1320" heatid="2106" lane="5" entrytime="00:01:25.05" entrycourse="SCM" />
                <RESULT eventid="1073" status="DNS" swimtime="00:00:00.00" resultid="1321" heatid="2085" lane="4" entrytime="00:03:21.95" entrycourse="SCM" />
                <RESULT eventid="1145" status="DNS" swimtime="00:00:00.00" resultid="1322" heatid="2175" lane="1" entrytime="00:00:46.88" entrycourse="SCM" />
                <RESULT eventid="1133" status="DNS" swimtime="00:00:00.00" resultid="1323" heatid="2156" lane="5" entrytime="00:01:43.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ravi" lastname="Osternack Erbe" birthdate="2013-08-10" gender="M" nation="BRA" license="372681" swrid="5588841" athleteid="1374" externalid="372681">
              <RESULTS>
                <RESULT eventid="1101" points="155" swimtime="00:00:40.45" resultid="1375" heatid="2120" lane="4" entrytime="00:00:40.08" entrycourse="SCM" />
                <RESULT eventid="1089" points="225" swimtime="00:01:13.69" resultid="1376" heatid="2107" lane="1" entrytime="00:01:22.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Vian" birthdate="2014-03-25" gender="F" nation="BRA" license="393919" swrid="5641779" athleteid="1662" externalid="393919">
              <RESULTS>
                <RESULT eventid="1092" points="79" swimtime="00:00:56.77" resultid="1663" heatid="2111" lane="8" entrytime="00:00:55.88" entrycourse="SCM" />
                <RESULT eventid="1064" points="136" swimtime="00:03:34.42" resultid="1664" heatid="2074" lane="4" entrytime="00:04:12.81" entrycourse="SCM" />
                <RESULT eventid="1124" points="145" swimtime="00:00:47.99" resultid="1665" heatid="2145" lane="7" entrytime="00:00:50.47" entrycourse="SCM" />
                <RESULT eventid="1111" points="123" swimtime="00:01:53.56" resultid="1666" heatid="2131" lane="1" entrytime="00:02:11.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Hadad" birthdate="2015-09-09" gender="M" nation="BRA" license="406740" swrid="5717272" athleteid="1717" externalid="406740">
              <RESULTS>
                <RESULT eventid="1083" points="49" swimtime="00:01:08.06" resultid="1718" heatid="2093" lane="7" />
                <RESULT eventid="1067" points="50" swimtime="00:04:29.11" resultid="1719" heatid="2077" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.60" />
                    <SPLIT distance="100" swimtime="00:02:11.91" />
                    <SPLIT distance="150" swimtime="00:03:20.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="33" swimtime="00:01:08.70" resultid="1720" heatid="2147" lane="6" entrytime="00:01:11.14" entrycourse="SCM" />
                <RESULT eventid="1114" points="43" swimtime="00:02:20.30" resultid="1721" heatid="2134" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:11.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Mayer Paludetto" birthdate="2012-10-30" gender="F" nation="BRA" license="369264" swrid="5588811" athleteid="1304" externalid="369264">
              <RESULTS>
                <RESULT eventid="1098" points="315" swimtime="00:00:35.81" resultid="1305" heatid="2117" lane="4" entrytime="00:00:36.12" entrycourse="SCM" />
                <RESULT eventid="1070" points="369" swimtime="00:02:49.82" resultid="1306" heatid="2083" lane="5" entrytime="00:03:00.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                    <SPLIT distance="100" swimtime="00:01:21.19" />
                    <SPLIT distance="150" swimtime="00:02:11.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="424" swimtime="00:05:07.86" resultid="1307" heatid="2123" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:13.26" />
                    <SPLIT distance="150" swimtime="00:01:53.13" />
                    <SPLIT distance="200" swimtime="00:02:32.39" />
                    <SPLIT distance="250" swimtime="00:03:12.04" />
                    <SPLIT distance="300" swimtime="00:03:51.41" />
                    <SPLIT distance="350" swimtime="00:04:30.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="311" swimtime="00:01:20.98" resultid="1308" heatid="2151" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.30" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Carcereri Navarro" birthdate="2013-12-19" gender="M" nation="BRA" license="376962" swrid="5588576" athleteid="1402" externalid="376962">
              <RESULTS>
                <RESULT eventid="1101" points="151" swimtime="00:00:40.82" resultid="1403" heatid="2121" lane="8" entrytime="00:00:39.92" entrycourse="SCM" />
                <RESULT eventid="1073" status="DSQ" swimtime="00:03:25.46" resultid="1404" heatid="2085" lane="5" entrytime="00:03:25.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.85" />
                    <SPLIT distance="100" swimtime="00:01:41.62" />
                    <SPLIT distance="150" swimtime="00:02:41.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="174" swimtime="00:00:44.61" resultid="1405" heatid="2175" lane="2" entrytime="00:00:46.50" entrycourse="SCM" />
                <RESULT eventid="1117" points="158" swimtime="00:06:32.58" resultid="1406" heatid="2137" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.73" />
                    <SPLIT distance="100" swimtime="00:01:31.71" />
                    <SPLIT distance="150" swimtime="00:02:21.85" />
                    <SPLIT distance="200" swimtime="00:03:12.57" />
                    <SPLIT distance="250" swimtime="00:04:03.72" />
                    <SPLIT distance="300" swimtime="00:04:55.91" />
                    <SPLIT distance="350" swimtime="00:05:45.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enrico" lastname="Hallage Bianchini" birthdate="2014-02-27" gender="M" nation="BRA" license="397164" swrid="5661348" athleteid="1667" externalid="397164">
              <RESULTS>
                <RESULT eventid="1095" status="DNS" swimtime="00:00:00.00" resultid="1668" heatid="2113" lane="2" entrytime="00:00:48.69" entrycourse="SCM" />
                <RESULT eventid="1067" status="DNS" swimtime="00:00:00.00" resultid="1669" heatid="2077" lane="7" />
                <RESULT eventid="1139" status="DNS" swimtime="00:00:00.00" resultid="1670" heatid="2166" lane="8" entrytime="00:00:39.66" entrycourse="SCM" />
                <RESULT eventid="1114" status="DNS" swimtime="00:00:00.00" resultid="1671" heatid="2134" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joana" lastname="Asinelli Casagrande" birthdate="2013-10-26" gender="F" nation="BRA" license="376970" swrid="5588536" athleteid="1421" externalid="376970">
              <RESULTS>
                <RESULT eventid="1098" points="206" swimtime="00:00:41.25" resultid="1422" heatid="2116" lane="3" entrytime="00:00:45.63" entrycourse="SCM" />
                <RESULT eventid="1070" status="DSQ" swimtime="00:03:20.06" resultid="1423" heatid="2082" lane="6" entrytime="00:03:39.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.59" />
                    <SPLIT distance="100" swimtime="00:01:38.12" />
                    <SPLIT distance="150" swimtime="00:02:36.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="220" swimtime="00:06:22.66" resultid="1424" heatid="2123" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.15" />
                    <SPLIT distance="100" swimtime="00:01:33.55" />
                    <SPLIT distance="150" swimtime="00:02:21.44" />
                    <SPLIT distance="200" swimtime="00:03:11.17" />
                    <SPLIT distance="250" swimtime="00:04:00.81" />
                    <SPLIT distance="300" swimtime="00:04:50.60" />
                    <SPLIT distance="350" swimtime="00:05:38.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="211" swimtime="00:01:32.07" resultid="1425" heatid="2151" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Guimaraes Mesquita" birthdate="2015-10-05" gender="F" nation="BRA" license="393263" swrid="5616444" athleteid="1648" externalid="393263">
              <RESULTS>
                <RESULT eventid="1080" points="55" swimtime="00:01:14.46" resultid="1649" heatid="2090" lane="8" />
                <RESULT eventid="1136" points="40" swimtime="00:01:07.03" resultid="1650" heatid="2159" lane="8" entrytime="00:01:15.20" entrycourse="SCM" />
                <RESULT eventid="1124" points="56" swimtime="00:01:05.90" resultid="1651" heatid="2143" lane="3" entrytime="00:01:06.79" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Albuquerque" birthdate="2012-11-16" gender="F" nation="BRA" license="369281" swrid="5602506" athleteid="1359" externalid="369281">
              <RESULTS>
                <RESULT eventid="1098" points="241" swimtime="00:00:39.17" resultid="1360" heatid="2114" lane="5" />
                <RESULT eventid="1070" points="312" swimtime="00:02:59.53" resultid="1361" heatid="2083" lane="7" entrytime="00:03:14.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.82" />
                    <SPLIT distance="100" swimtime="00:01:27.38" />
                    <SPLIT distance="150" swimtime="00:02:20.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="336" swimtime="00:05:32.44" resultid="1362" heatid="2125" lane="7" entrytime="00:05:58.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:19.61" />
                    <SPLIT distance="150" swimtime="00:02:01.83" />
                    <SPLIT distance="200" swimtime="00:02:44.88" />
                    <SPLIT distance="250" swimtime="00:03:27.22" />
                    <SPLIT distance="300" swimtime="00:04:10.24" />
                    <SPLIT distance="350" swimtime="00:04:52.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="285" swimtime="00:00:43.09" resultid="1363" heatid="2171" lane="6" entrytime="00:00:46.76" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Alice Silva Gomes Xavier" birthdate="2013-02-25" gender="F" nation="BRA" license="371040" swrid="5717241" athleteid="1784" externalid="371040">
              <RESULTS>
                <RESULT eventid="1098" points="241" swimtime="00:00:39.17" resultid="1785" heatid="2117" lane="1" entrytime="00:00:40.03" entrycourse="SCM" />
                <RESULT eventid="1070" points="229" swimtime="00:03:19.05" resultid="1786" heatid="2081" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.62" />
                    <SPLIT distance="100" swimtime="00:01:38.91" />
                    <SPLIT distance="150" swimtime="00:02:36.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="305" swimtime="00:05:43.51" resultid="1787" heatid="2122" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.56" />
                    <SPLIT distance="100" swimtime="00:01:23.53" />
                    <SPLIT distance="150" swimtime="00:02:07.84" />
                    <SPLIT distance="200" swimtime="00:02:51.45" />
                    <SPLIT distance="250" swimtime="00:03:35.52" />
                    <SPLIT distance="300" swimtime="00:04:19.52" />
                    <SPLIT distance="350" swimtime="00:05:02.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="278" swimtime="00:00:43.45" resultid="1788" heatid="2171" lane="3" entrytime="00:00:46.60" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Pisani Ferreira" birthdate="2014-01-26" gender="M" nation="BRA" license="391017" swrid="5602570" athleteid="1563" externalid="391017">
              <RESULTS>
                <RESULT eventid="1083" points="115" swimtime="00:00:51.28" resultid="1564" heatid="2096" lane="1" entrytime="00:00:55.62" entrycourse="SCM" />
                <RESULT eventid="1067" points="108" swimtime="00:03:28.57" resultid="1565" heatid="2078" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.44" />
                    <SPLIT distance="100" swimtime="00:01:38.13" />
                    <SPLIT distance="150" swimtime="00:02:33.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="112" swimtime="00:00:41.72" resultid="1566" heatid="2165" lane="7" entrytime="00:00:42.99" entrycourse="SCM" />
                <RESULT eventid="1114" points="99" swimtime="00:01:46.18" resultid="1567" heatid="2135" lane="7" entrytime="00:02:04.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luisa" lastname="Della Villa Yang" birthdate="2012-10-08" gender="F" nation="BRA" license="369276" swrid="5588653" athleteid="1339" externalid="369276">
              <RESULTS>
                <RESULT eventid="1098" points="276" swimtime="00:00:37.44" resultid="1340" heatid="2117" lane="6" entrytime="00:00:39.42" entrycourse="SCM" />
                <RESULT eventid="1070" points="344" swimtime="00:02:53.77" resultid="1341" heatid="2083" lane="2" entrytime="00:03:13.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                    <SPLIT distance="100" swimtime="00:01:23.17" />
                    <SPLIT distance="150" swimtime="00:02:17.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="409" swimtime="00:05:11.41" resultid="1342" heatid="2125" lane="5" entrytime="00:05:22.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.10" />
                    <SPLIT distance="100" swimtime="00:01:15.78" />
                    <SPLIT distance="150" swimtime="00:01:55.91" />
                    <SPLIT distance="200" swimtime="00:02:35.87" />
                    <SPLIT distance="250" swimtime="00:03:15.66" />
                    <SPLIT distance="300" swimtime="00:03:54.33" />
                    <SPLIT distance="350" swimtime="00:04:33.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="234" swimtime="00:00:45.98" resultid="1343" heatid="2167" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia" lastname="Ziliotto Mehl" birthdate="2015-10-09" gender="F" nation="BRA" license="400122" swrid="5652905" athleteid="1702" externalid="400122">
              <RESULTS>
                <RESULT eventid="1080" points="107" swimtime="00:00:59.63" resultid="1703" heatid="2091" lane="2" entrytime="00:01:03.12" entrycourse="SCM" />
                <RESULT eventid="1064" status="DNS" swimtime="00:00:00.00" resultid="1704" heatid="2073" lane="4" />
                <RESULT eventid="1136" status="DNS" swimtime="00:00:00.00" resultid="1705" heatid="2160" lane="8" entrytime="00:00:51.36" entrycourse="SCM" />
                <RESULT eventid="1111" status="DNS" swimtime="00:00:00.00" resultid="1706" heatid="2130" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Afonso Fowler" birthdate="2014-01-22" gender="M" nation="BRA" license="393264" swrid="5661338" athleteid="1652" externalid="393264">
              <RESULTS>
                <RESULT eventid="1095" status="DNS" swimtime="00:00:00.00" resultid="1653" heatid="2112" lane="5" entrytime="00:01:02.85" entrycourse="SCM" />
                <RESULT eventid="1067" status="DNS" swimtime="00:00:00.00" resultid="1654" heatid="2079" lane="2" />
                <RESULT eventid="1127" status="DNS" swimtime="00:00:00.00" resultid="1655" heatid="2148" lane="6" entrytime="00:00:53.27" entrycourse="SCM" />
                <RESULT eventid="1114" status="DNS" swimtime="00:00:00.00" resultid="1656" heatid="2133" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Wolf Macedo" birthdate="2012-01-27" gender="F" nation="BRA" license="369277" swrid="5602592" athleteid="1344" externalid="369277">
              <RESULTS>
                <RESULT eventid="1098" points="360" swimtime="00:00:34.24" resultid="1345" heatid="2117" lane="5" entrytime="00:00:36.22" entrycourse="SCM" />
                <RESULT eventid="1086" points="373" swimtime="00:01:09.77" resultid="1346" heatid="2102" lane="2" entrytime="00:01:14.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="361" swimtime="00:05:24.59" resultid="1347" heatid="2125" lane="3" entrytime="00:05:31.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:15.49" />
                    <SPLIT distance="150" swimtime="00:01:56.44" />
                    <SPLIT distance="200" swimtime="00:02:37.86" />
                    <SPLIT distance="250" swimtime="00:03:19.33" />
                    <SPLIT distance="300" swimtime="00:04:02.04" />
                    <SPLIT distance="350" swimtime="00:04:44.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="277" swimtime="00:00:43.49" resultid="1348" heatid="2169" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Lazzarotti Matias" birthdate="2012-03-19" gender="F" nation="BRA" license="391026" swrid="5602552" athleteid="1598" externalid="391026">
              <RESULTS>
                <RESULT eventid="1086" points="336" swimtime="00:01:12.24" resultid="1599" heatid="2102" lane="1" entrytime="00:01:17.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1070" points="311" swimtime="00:02:59.73" resultid="1600" heatid="2082" lane="5" entrytime="00:03:21.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                    <SPLIT distance="100" swimtime="00:01:27.68" />
                    <SPLIT distance="150" swimtime="00:02:22.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="257" swimtime="00:00:44.61" resultid="1601" heatid="2171" lane="1" entrytime="00:00:50.13" entrycourse="SCM" />
                <RESULT eventid="1130" points="293" swimtime="00:01:22.62" resultid="1602" heatid="2152" lane="6" entrytime="00:01:26.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Rossi Mattioli" birthdate="2013-05-08" gender="F" nation="BRA" license="376988" swrid="5588892" athleteid="1489" externalid="376988">
              <RESULTS>
                <RESULT eventid="1086" points="273" swimtime="00:01:17.43" resultid="1490" heatid="2101" lane="4" entrytime="00:01:19.37" entrycourse="SCM" />
                <RESULT eventid="1070" points="237" swimtime="00:03:16.65" resultid="1491" heatid="2083" lane="8" entrytime="00:03:18.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.01" />
                    <SPLIT distance="100" swimtime="00:01:34.44" />
                    <SPLIT distance="150" swimtime="00:02:32.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="253" swimtime="00:06:05.42" resultid="1492" heatid="2124" lane="4" />
                <RESULT eventid="1142" points="215" swimtime="00:00:47.29" resultid="1493" heatid="2171" lane="7" entrytime="00:00:48.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Pacheco" birthdate="2012-10-13" gender="F" nation="BRA" license="376981" swrid="5602566" athleteid="1446" externalid="376981">
              <RESULTS>
                <RESULT eventid="1098" points="86" swimtime="00:00:55.16" resultid="1447" heatid="2115" lane="3" entrytime="00:01:06.51" entrycourse="SCM" />
                <RESULT eventid="1086" points="219" swimtime="00:01:23.30" resultid="1448" heatid="2100" lane="6" entrytime="00:01:34.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="211" swimtime="00:06:28.40" resultid="1449" heatid="2125" lane="8" entrytime="00:07:22.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.19" />
                    <SPLIT distance="100" swimtime="00:01:32.45" />
                    <SPLIT distance="150" swimtime="00:02:23.77" />
                    <SPLIT distance="200" swimtime="00:03:14.81" />
                    <SPLIT distance="250" swimtime="00:04:05.19" />
                    <SPLIT distance="300" swimtime="00:04:53.94" />
                    <SPLIT distance="350" swimtime="00:05:43.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="174" swimtime="00:00:50.76" resultid="1450" heatid="2170" lane="6" entrytime="00:00:54.22" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Nishimura Ramina" birthdate="2013-11-25" gender="M" nation="BRA" license="376989" swrid="5588831" athleteid="1484" externalid="376989">
              <RESULTS>
                <RESULT eventid="1101" points="102" swimtime="00:00:46.55" resultid="1485" heatid="2119" lane="6" entrytime="00:00:51.88" entrycourse="SCM" />
                <RESULT eventid="1089" points="118" swimtime="00:01:31.31" resultid="1486" heatid="2105" lane="5" entrytime="00:01:39.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="103" swimtime="00:01:42.98" resultid="1487" heatid="2154" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="152" swimtime="00:06:37.32" resultid="1488" heatid="2137" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.60" />
                    <SPLIT distance="100" swimtime="00:01:31.84" />
                    <SPLIT distance="150" swimtime="00:02:21.62" />
                    <SPLIT distance="200" swimtime="00:03:13.29" />
                    <SPLIT distance="250" swimtime="00:04:03.66" />
                    <SPLIT distance="300" swimtime="00:04:56.14" />
                    <SPLIT distance="350" swimtime="00:05:46.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gael" lastname="Stramandinoli Zanicotti" birthdate="2015-03-21" gender="M" nation="BRA" license="406954" swrid="5717298" athleteid="1789" externalid="406954">
              <RESULTS>
                <RESULT eventid="1095" points="6" swimtime="00:01:54.14" resultid="1790" heatid="2112" lane="3" entrytime="00:01:31.38" entrycourse="SCM" />
                <RESULT eventid="1083" points="19" swimtime="00:01:32.93" resultid="1791" heatid="2094" lane="7" />
                <RESULT eventid="1127" points="25" swimtime="00:01:14.77" resultid="1792" heatid="2147" lane="5" entrytime="00:01:07.50" entrycourse="SCM" />
                <RESULT eventid="1114" points="22" swimtime="00:02:55.06" resultid="1793" heatid="2133" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:26.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Guimaraes Mesquita" birthdate="2013-12-30" gender="F" nation="BRA" license="391027" swrid="5602544" athleteid="1603" externalid="391027">
              <RESULTS>
                <RESULT eventid="1086" points="152" swimtime="00:01:33.99" resultid="1604" heatid="2100" lane="1" entrytime="00:01:40.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1070" status="DSQ" swimtime="00:03:48.08" resultid="1605" heatid="2082" lane="1" entrytime="00:04:07.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.81" />
                    <SPLIT distance="100" swimtime="00:01:57.43" />
                    <SPLIT distance="150" swimtime="00:03:00.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="158" swimtime="00:07:07.55" resultid="1606" heatid="2124" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.72" />
                    <SPLIT distance="100" swimtime="00:01:43.01" />
                    <SPLIT distance="150" swimtime="00:02:38.45" />
                    <SPLIT distance="200" swimtime="00:03:34.64" />
                    <SPLIT distance="250" swimtime="00:04:29.97" />
                    <SPLIT distance="300" swimtime="00:05:24.69" />
                    <SPLIT distance="350" swimtime="00:06:17.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" status="DSQ" swimtime="00:00:55.27" resultid="1607" heatid="2170" lane="7" entrytime="00:00:58.22" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Francia Soares" birthdate="2014-06-01" gender="F" nation="BRA" license="391011" swrid="5602540" athleteid="1553" externalid="391011">
              <RESULTS>
                <RESULT eventid="1092" points="49" swimtime="00:01:06.21" resultid="1554" heatid="2109" lane="7" />
                <RESULT eventid="1064" points="117" swimtime="00:03:45.37" resultid="1555" heatid="2074" lane="5" entrytime="00:04:17.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.27" />
                    <SPLIT distance="100" swimtime="00:01:52.38" />
                    <SPLIT distance="150" swimtime="00:02:53.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="138" swimtime="00:00:44.34" resultid="1556" heatid="2159" lane="4" entrytime="00:00:54.66" entrycourse="SCM" />
                <RESULT eventid="1111" points="81" swimtime="00:02:10.44" resultid="1557" heatid="2130" lane="5" entrytime="00:02:35.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="De Macedo Martynychen" birthdate="2015-06-12" gender="F" nation="BRA" license="399681" swrid="5652885" athleteid="1692" externalid="399681">
              <RESULTS>
                <RESULT eventid="1092" points="59" swimtime="00:01:02.44" resultid="1693" heatid="2110" lane="2" entrytime="00:01:06.67" entrycourse="SCM" />
                <RESULT eventid="1064" points="71" swimtime="00:04:25.59" resultid="1694" heatid="2072" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.52" />
                    <SPLIT distance="100" swimtime="00:02:07.76" />
                    <SPLIT distance="150" swimtime="00:03:18.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="59" swimtime="00:01:04.80" resultid="1695" heatid="2143" lane="6" entrytime="00:01:08.54" entrycourse="SCM" />
                <RESULT eventid="1111" points="76" swimtime="00:02:12.86" resultid="1696" heatid="2129" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:03.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Wolff Contin" birthdate="2015-10-10" gender="M" nation="BRA" license="406745" swrid="5717303" athleteid="1739" externalid="406745">
              <RESULTS>
                <RESULT eventid="1083" points="35" swimtime="00:01:15.58" resultid="1740" heatid="2094" lane="6" entrytime="00:01:28.47" entrycourse="SCM" />
                <RESULT eventid="1067" points="46" swimtime="00:04:36.85" resultid="1741" heatid="2076" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.12" />
                    <SPLIT distance="100" swimtime="00:02:11.24" />
                    <SPLIT distance="150" swimtime="00:03:26.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="60" swimtime="00:00:51.33" resultid="1742" heatid="2164" lane="8" entrytime="00:01:02.31" entrycourse="SCM" />
                <RESULT eventid="1127" points="43" swimtime="00:01:03.08" resultid="1743" heatid="2147" lane="3" entrytime="00:01:07.72" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Garcia" birthdate="2015-10-26" gender="M" nation="BRA" license="406967" swrid="5717271" athleteid="1803" externalid="406967">
              <RESULTS>
                <RESULT eventid="1083" status="DNS" swimtime="00:00:00.00" resultid="1804" heatid="2094" lane="2" entrytime="00:01:34.42" entrycourse="SCM" />
                <RESULT eventid="1067" status="DNS" swimtime="00:00:00.00" resultid="1805" heatid="2078" lane="3" />
                <RESULT eventid="1139" status="DNS" swimtime="00:00:00.00" resultid="1806" heatid="2163" lane="2" entrytime="00:01:16.80" entrycourse="SCM" />
                <RESULT eventid="1114" status="DNS" swimtime="00:00:00.00" resultid="1807" heatid="2132" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Da Cunha Souza" birthdate="2013-09-17" gender="M" nation="BRA" license="376975" swrid="5588618" athleteid="1431" externalid="376975">
              <RESULTS>
                <RESULT eventid="1101" points="100" swimtime="00:00:46.74" resultid="1432" heatid="2119" lane="3" entrytime="00:00:49.38" entrycourse="SCM" />
                <RESULT eventid="1089" points="139" swimtime="00:01:26.40" resultid="1433" heatid="2106" lane="7" entrytime="00:01:31.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="94" swimtime="00:00:54.82" resultid="1434" heatid="2173" lane="5" entrytime="00:01:01.79" entrycourse="SCM" />
                <RESULT eventid="1117" points="166" swimtime="00:06:25.53" resultid="1435" heatid="2136" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                    <SPLIT distance="100" swimtime="00:01:26.95" />
                    <SPLIT distance="150" swimtime="00:02:17.95" />
                    <SPLIT distance="200" swimtime="00:03:09.22" />
                    <SPLIT distance="250" swimtime="00:03:59.30" />
                    <SPLIT distance="300" swimtime="00:04:50.21" />
                    <SPLIT distance="350" swimtime="00:05:37.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Sieczkowski Pacheco" birthdate="2015-11-20" gender="F" nation="BRA" license="393261" swrid="5616450" athleteid="1638" externalid="393261">
              <RESULTS>
                <RESULT eventid="1080" points="128" swimtime="00:00:56.24" resultid="1639" heatid="2092" lane="7" entrytime="00:00:58.63" entrycourse="SCM" />
                <RESULT eventid="1064" points="100" swimtime="00:03:57.22" resultid="1640" heatid="2074" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.98" />
                    <SPLIT distance="100" swimtime="00:01:53.65" />
                    <SPLIT distance="150" swimtime="00:02:56.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="92" swimtime="00:00:55.86" resultid="1641" heatid="2144" lane="6" entrytime="00:00:57.45" entrycourse="SCM" />
                <RESULT eventid="1111" points="100" swimtime="00:02:01.62" resultid="1642" heatid="2129" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="De Moraes" birthdate="2014-09-18" gender="M" nation="BRA" license="391024" swrid="5602529" athleteid="1588" externalid="391024">
              <RESULTS>
                <RESULT eventid="1083" points="122" swimtime="00:00:50.20" resultid="1589" heatid="2096" lane="5" entrytime="00:00:51.67" entrycourse="SCM" />
                <RESULT eventid="1067" points="161" swimtime="00:03:02.41" resultid="1590" heatid="2080" lane="3" entrytime="00:03:13.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.25" />
                    <SPLIT distance="100" swimtime="00:01:29.51" />
                    <SPLIT distance="150" swimtime="00:02:18.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="198" swimtime="00:00:34.56" resultid="1591" heatid="2166" lane="4" entrytime="00:00:35.90" entrycourse="SCM" />
                <RESULT eventid="1114" points="132" swimtime="00:01:36.75" resultid="1592" heatid="2135" lane="6" entrytime="00:01:53.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Almeida Jorge" birthdate="2015-05-27" gender="M" nation="BRA" license="406836" swrid="5717242" athleteid="1774" externalid="406836">
              <RESULTS>
                <RESULT eventid="1083" points="48" swimtime="00:01:08.63" resultid="1775" heatid="2095" lane="8" entrytime="00:01:09.86" entrycourse="SCM" />
                <RESULT eventid="1067" points="38" swimtime="00:04:54.50" resultid="1776" heatid="2078" lane="1" />
                <RESULT eventid="1139" points="31" swimtime="00:01:04.14" resultid="1777" heatid="2163" lane="3" entrytime="00:01:07.06" entrycourse="SCM" />
                <RESULT eventid="1114" points="42" swimtime="00:02:21.20" resultid="1778" heatid="2133" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:08.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Schiavo Vianna" birthdate="2013-04-27" gender="F" nation="BRA" license="391005" swrid="5602582" athleteid="1538" externalid="391005">
              <RESULTS>
                <RESULT eventid="1098" points="82" swimtime="00:00:55.93" resultid="1539" heatid="2114" lane="7" />
                <RESULT eventid="1086" points="155" swimtime="00:01:33.54" resultid="1540" heatid="2099" lane="6" entrytime="00:01:43.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="147" swimtime="00:07:18.05" resultid="1541" heatid="2124" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.98" />
                    <SPLIT distance="100" swimtime="00:01:45.78" />
                    <SPLIT distance="150" swimtime="00:02:42.66" />
                    <SPLIT distance="200" swimtime="00:03:43.55" />
                    <SPLIT distance="250" swimtime="00:04:36.85" />
                    <SPLIT distance="300" swimtime="00:05:33.96" />
                    <SPLIT distance="350" swimtime="00:06:30.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="198" swimtime="00:00:48.64" resultid="1542" heatid="2170" lane="3" entrytime="00:00:53.40" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Henrique Tiboni Araujo" birthdate="2013-06-11" gender="M" nation="BRA" license="376968" swrid="5588747" athleteid="1416" externalid="376968">
              <RESULTS>
                <RESULT eventid="1089" points="130" swimtime="00:01:28.29" resultid="1417" heatid="2106" lane="1" entrytime="00:01:34.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1073" points="118" swimtime="00:03:43.50" resultid="1418" heatid="2085" lane="8" entrytime="00:04:02.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.29" />
                    <SPLIT distance="100" swimtime="00:01:44.95" />
                    <SPLIT distance="150" swimtime="00:02:54.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="99" swimtime="00:01:44.24" resultid="1419" heatid="2156" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="129" swimtime="00:06:59.21" resultid="1420" heatid="2138" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.20" />
                    <SPLIT distance="100" swimtime="00:01:37.20" />
                    <SPLIT distance="150" swimtime="00:02:31.83" />
                    <SPLIT distance="200" swimtime="00:03:25.44" />
                    <SPLIT distance="250" swimtime="00:04:20.84" />
                    <SPLIT distance="300" swimtime="00:05:16.07" />
                    <SPLIT distance="350" swimtime="00:06:09.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Ribas Luz" birthdate="2015-02-05" gender="F" nation="BRA" license="406743" swrid="5717291" athleteid="1732" externalid="406743">
              <RESULTS>
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="1733" heatid="2090" lane="7" entrytime="00:01:30.45" entrycourse="SCM" />
                <RESULT eventid="1136" status="DNS" swimtime="00:00:00.00" resultid="1734" heatid="2159" lane="1" entrytime="00:01:05.73" entrycourse="SCM" />
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="1735" heatid="2143" lane="7" entrytime="00:01:11.89" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Xavier Jardim" birthdate="2012-01-23" gender="M" nation="BRA" license="369259" swrid="5641781" athleteid="1289" externalid="369259">
              <RESULTS>
                <RESULT eventid="1101" points="168" swimtime="00:00:39.40" resultid="1290" heatid="2121" lane="7" entrytime="00:00:38.26" entrycourse="SCM" />
                <RESULT eventid="1089" points="250" swimtime="00:01:11.10" resultid="1291" heatid="2108" lane="3" entrytime="00:01:11.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="178" swimtime="00:01:25.79" resultid="1292" heatid="2157" lane="2" entrytime="00:01:29.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="245" swimtime="00:05:39.13" resultid="1293" heatid="2136" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                    <SPLIT distance="100" swimtime="00:01:20.00" />
                    <SPLIT distance="150" swimtime="00:02:03.50" />
                    <SPLIT distance="200" swimtime="00:02:47.97" />
                    <SPLIT distance="250" swimtime="00:03:31.69" />
                    <SPLIT distance="300" swimtime="00:04:15.07" />
                    <SPLIT distance="350" swimtime="00:04:57.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="De Fortes" birthdate="2015-06-01" gender="M" nation="BRA" license="399680" swrid="5652884" athleteid="1687" externalid="399680">
              <RESULTS>
                <RESULT eventid="1095" points="52" swimtime="00:00:57.94" resultid="1688" heatid="2112" lane="4" entrytime="00:00:57.78" entrycourse="SCM" />
                <RESULT eventid="1067" points="71" swimtime="00:03:59.78" resultid="1689" heatid="2079" lane="4" />
                <RESULT eventid="1127" points="69" swimtime="00:00:53.70" resultid="1690" heatid="2148" lane="2" entrytime="00:00:56.53" entrycourse="SCM" />
                <RESULT eventid="1114" points="61" swimtime="00:02:04.64" resultid="1691" heatid="2134" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Vanzo Assumpcao" birthdate="2012-05-15" gender="M" nation="BRA" license="369258" swrid="5588942" athleteid="1284" externalid="369258">
              <RESULTS>
                <RESULT eventid="1101" points="291" swimtime="00:00:32.82" resultid="1285" heatid="2121" lane="4" entrytime="00:00:33.99" entrycourse="SCM" />
                <RESULT eventid="1073" points="257" swimtime="00:02:52.25" resultid="1286" heatid="2086" lane="5" entrytime="00:02:54.09" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.25" />
                    <SPLIT distance="100" swimtime="00:01:20.86" />
                    <SPLIT distance="150" swimtime="00:02:14.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="227" swimtime="00:01:19.19" resultid="1287" heatid="2157" lane="6" entrytime="00:01:27.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="290" swimtime="00:05:20.58" resultid="1288" heatid="2138" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Toscani Kim" birthdate="2013-02-15" gender="F" nation="BRA" license="372683" swrid="5588939" athleteid="1382" externalid="372683">
              <RESULTS>
                <RESULT eventid="1098" points="243" swimtime="00:00:39.05" resultid="1383" heatid="2117" lane="7" entrytime="00:00:39.90" entrycourse="SCM" />
                <RESULT eventid="1070" points="306" swimtime="00:03:00.65" resultid="1384" heatid="2083" lane="6" entrytime="00:03:08.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:01:27.56" />
                    <SPLIT distance="150" swimtime="00:02:19.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="288" swimtime="00:05:49.86" resultid="1385" heatid="2123" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                    <SPLIT distance="100" swimtime="00:01:23.25" />
                    <SPLIT distance="150" swimtime="00:02:07.93" />
                    <SPLIT distance="200" swimtime="00:02:52.65" />
                    <SPLIT distance="250" swimtime="00:03:37.68" />
                    <SPLIT distance="300" swimtime="00:04:21.35" />
                    <SPLIT distance="350" swimtime="00:05:06.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="277" swimtime="00:00:43.52" resultid="1386" heatid="2171" lane="5" entrytime="00:00:45.06" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Dolberth Alcantara" birthdate="2014-09-26" gender="F" nation="BRA" license="382124" swrid="5602532" athleteid="1518" externalid="382124">
              <RESULTS>
                <RESULT eventid="1092" points="98" swimtime="00:00:52.71" resultid="1519" heatid="2110" lane="4" entrytime="00:00:56.61" entrycourse="SCM" />
                <RESULT eventid="1064" points="131" swimtime="00:03:36.70" resultid="1520" heatid="2075" lane="1" entrytime="00:03:57.65" entrycourse="SCM" />
                <RESULT eventid="1124" points="116" swimtime="00:00:51.72" resultid="1521" heatid="2145" lane="8" entrytime="00:00:54.49" entrycourse="SCM" />
                <RESULT eventid="1111" points="134" swimtime="00:01:50.42" resultid="1522" heatid="2131" lane="6" entrytime="00:02:05.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Szpak Zraik" birthdate="2015-04-10" gender="M" nation="BRA" license="393259" swrid="5616451" athleteid="1628" externalid="393259">
              <RESULTS>
                <RESULT eventid="1083" points="134" swimtime="00:00:48.65" resultid="1629" heatid="2096" lane="3" entrytime="00:00:53.33" entrycourse="SCM" />
                <RESULT eventid="1067" points="85" swimtime="00:03:45.71" resultid="1630" heatid="2078" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.26" />
                    <SPLIT distance="100" swimtime="00:01:42.26" />
                    <SPLIT distance="150" swimtime="00:02:45.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="100" swimtime="00:00:43.41" resultid="1631" heatid="2164" lane="3" entrytime="00:00:45.52" entrycourse="SCM" />
                <RESULT eventid="1114" points="78" swimtime="00:01:55.02" resultid="1632" heatid="2133" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Lauand Lorenci" birthdate="2013-03-06" gender="M" nation="BRA" license="376982" swrid="5588764" athleteid="1451" externalid="376982">
              <RESULTS>
                <RESULT eventid="1101" points="147" swimtime="00:00:41.18" resultid="1452" heatid="2120" lane="8" entrytime="00:00:44.75" entrycourse="SCM" />
                <RESULT eventid="1073" points="180" swimtime="00:03:14.01" resultid="1453" heatid="2085" lane="6" entrytime="00:03:28.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.21" />
                    <SPLIT distance="100" swimtime="00:01:37.52" />
                    <SPLIT distance="150" swimtime="00:02:30.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="196" swimtime="00:00:42.91" resultid="1454" heatid="2175" lane="7" entrytime="00:00:46.59" entrycourse="SCM" />
                <RESULT eventid="1117" points="173" swimtime="00:06:20.26" resultid="1455" heatid="2138" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.28" />
                    <SPLIT distance="100" swimtime="00:01:30.62" />
                    <SPLIT distance="150" swimtime="00:02:19.95" />
                    <SPLIT distance="200" swimtime="00:03:09.70" />
                    <SPLIT distance="250" swimtime="00:03:58.45" />
                    <SPLIT distance="300" swimtime="00:04:47.75" />
                    <SPLIT distance="350" swimtime="00:05:35.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Fernandes Tramujas" birthdate="2015-01-15" gender="F" nation="BRA" license="406750" swrid="5717263" athleteid="1764" externalid="406750">
              <RESULTS>
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="1765" heatid="2090" lane="5" entrytime="00:01:13.59" entrycourse="SCM" />
                <RESULT eventid="1064" status="DNS" swimtime="00:00:00.00" resultid="1766" heatid="2073" lane="3" />
                <RESULT eventid="1136" status="DNS" swimtime="00:00:00.00" resultid="1767" heatid="2158" lane="7" />
                <RESULT eventid="1111" status="DNS" swimtime="00:00:00.00" resultid="1768" heatid="2130" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Magalhaes Dabul" birthdate="2014-01-05" gender="M" nation="BRA" license="391023" swrid="5602555" athleteid="1583" externalid="391023">
              <RESULTS>
                <RESULT eventid="1095" points="97" swimtime="00:00:47.28" resultid="1584" heatid="2113" lane="1" entrytime="00:00:52.71" entrycourse="SCM" />
                <RESULT eventid="1067" points="120" swimtime="00:03:21.24" resultid="1585" heatid="2080" lane="1" entrytime="00:04:18.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.53" />
                    <SPLIT distance="100" swimtime="00:01:36.20" />
                    <SPLIT distance="150" swimtime="00:02:30.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="115" swimtime="00:00:41.45" resultid="1586" heatid="2165" lane="1" entrytime="00:00:43.07" entrycourse="SCM" />
                <RESULT eventid="1114" points="91" swimtime="00:01:49.47" resultid="1587" heatid="2135" lane="1" entrytime="00:02:10.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Trevisan De Paula" birthdate="2014-01-27" gender="M" nation="BRA" license="377152" swrid="5602568" athleteid="1503" externalid="377152">
              <RESULTS>
                <RESULT eventid="1095" points="174" swimtime="00:00:38.93" resultid="1504" heatid="2113" lane="4" entrytime="00:00:38.31" entrycourse="SCM" />
                <RESULT eventid="1067" points="203" swimtime="00:02:48.89" resultid="1505" heatid="2080" lane="4" entrytime="00:03:01.52" entrycourse="SCM" />
                <RESULT eventid="1127" points="146" swimtime="00:00:41.90" resultid="1506" heatid="2148" lane="4" entrytime="00:00:40.67" entrycourse="SCM" />
                <RESULT eventid="1114" points="164" swimtime="00:01:29.95" resultid="1507" heatid="2135" lane="4" entrytime="00:01:36.33" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Viera Correa" birthdate="2012-03-07" gender="M" nation="BRA" license="369269" swrid="5602590" athleteid="1314" externalid="369269">
              <RESULTS>
                <RESULT eventid="1101" points="202" swimtime="00:00:37.05" resultid="1315" heatid="2120" lane="3" entrytime="00:00:41.36" entrycourse="SCM" />
                <RESULT eventid="1089" points="285" swimtime="00:01:08.12" resultid="1316" heatid="2108" lane="7" entrytime="00:01:12.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="211" swimtime="00:01:21.10" resultid="1317" heatid="2157" lane="5" entrytime="00:01:24.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="272" swimtime="00:05:27.58" resultid="1318" heatid="2139" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:17.33" />
                    <SPLIT distance="150" swimtime="00:01:59.88" />
                    <SPLIT distance="200" swimtime="00:02:42.34" />
                    <SPLIT distance="250" swimtime="00:03:23.97" />
                    <SPLIT distance="300" swimtime="00:04:05.99" />
                    <SPLIT distance="350" swimtime="00:04:48.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Simioni Albuquerque" birthdate="2014-12-23" gender="F" nation="BRA" license="401980" swrid="5661355" athleteid="1707" externalid="401980">
              <RESULTS>
                <RESULT eventid="1092" points="113" swimtime="00:00:50.35" resultid="1708" heatid="2111" lane="3" entrytime="00:00:49.56" entrycourse="SCM" />
                <RESULT eventid="1064" points="115" swimtime="00:03:46.80" resultid="1709" heatid="2073" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.69" />
                    <SPLIT distance="100" swimtime="00:01:48.93" />
                    <SPLIT distance="150" swimtime="00:02:51.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="170" swimtime="00:00:41.39" resultid="1710" heatid="2158" lane="2" />
                <RESULT eventid="1111" points="132" swimtime="00:01:50.97" resultid="1711" heatid="2128" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Della Villa Yang" birthdate="2015-02-27" gender="F" nation="BRA" license="393283" swrid="5616442" athleteid="1657" externalid="393283">
              <RESULTS>
                <RESULT eventid="1092" points="80" swimtime="00:00:56.53" resultid="1658" heatid="2111" lane="1" entrytime="00:00:55.39" entrycourse="SCM" />
                <RESULT eventid="1064" points="122" swimtime="00:03:41.88" resultid="1659" heatid="2073" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.50" />
                    <SPLIT distance="100" swimtime="00:01:48.30" />
                    <SPLIT distance="150" swimtime="00:02:47.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="89" swimtime="00:00:56.36" resultid="1660" heatid="2144" lane="8" entrytime="00:01:02.14" entrycourse="SCM" />
                <RESULT eventid="1111" points="127" swimtime="00:01:52.33" resultid="1661" heatid="2128" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Gois Nogueira" birthdate="2014-03-11" gender="F" nation="BRA" license="393258" swrid="5616443" athleteid="1623" externalid="393258">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="1624" heatid="2110" lane="8" entrytime="00:01:07.15" entrycourse="SCM" />
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="1625" heatid="2091" lane="1" entrytime="00:01:04.50" entrycourse="SCM" />
                <RESULT eventid="1136" status="DNS" swimtime="00:00:00.00" resultid="1626" heatid="2160" lane="5" entrytime="00:00:47.06" entrycourse="SCM" />
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="1627" heatid="2144" lane="2" entrytime="00:00:57.92" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Felipe Canalli" birthdate="2015-12-23" gender="M" nation="BRA" license="406749" swrid="5717261" athleteid="1759" externalid="406749">
              <RESULTS>
                <RESULT eventid="1083" points="85" swimtime="00:00:56.66" resultid="1760" heatid="2096" lane="6" entrytime="00:00:55.35" entrycourse="SCM" />
                <RESULT eventid="1067" points="42" swimtime="00:04:44.07" resultid="1761" heatid="2076" lane="4" />
                <RESULT eventid="1127" points="38" swimtime="00:01:05.26" resultid="1762" heatid="2146" lane="5" />
                <RESULT eventid="1114" points="50" swimtime="00:02:13.74" resultid="1763" heatid="2134" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Karam Barbosa Lima" birthdate="2012-12-11" gender="F" nation="BRA" license="376956" swrid="5588758" athleteid="1387" externalid="376956">
              <RESULTS>
                <RESULT eventid="1086" points="331" swimtime="00:01:12.62" resultid="1388" heatid="2102" lane="5" entrytime="00:01:12.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1070" points="282" swimtime="00:03:05.64" resultid="1389" heatid="2082" lane="3" entrytime="00:03:29.66" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.02" />
                    <SPLIT distance="100" swimtime="00:01:27.67" />
                    <SPLIT distance="150" swimtime="00:02:26.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="322" swimtime="00:05:37.27" resultid="1390" heatid="2125" lane="2" entrytime="00:05:52.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:19.23" />
                    <SPLIT distance="150" swimtime="00:02:02.94" />
                    <SPLIT distance="200" swimtime="00:02:46.97" />
                    <SPLIT distance="250" swimtime="00:03:30.56" />
                    <SPLIT distance="300" swimtime="00:04:13.82" />
                    <SPLIT distance="350" swimtime="00:04:56.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="281" swimtime="00:01:23.80" resultid="1391" heatid="2152" lane="2" entrytime="00:01:29.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Fernandes  Dos Reis" birthdate="2012-09-18" gender="M" nation="BRA" license="369279" swrid="5588696" athleteid="1354" externalid="369279">
              <RESULTS>
                <RESULT eventid="1101" points="262" swimtime="00:00:33.97" resultid="1355" heatid="2121" lane="3" entrytime="00:00:36.91" entrycourse="SCM" />
                <RESULT eventid="1073" points="212" swimtime="00:03:03.85" resultid="1356" heatid="2086" lane="1" entrytime="00:03:19.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:26.30" />
                    <SPLIT distance="150" swimtime="00:02:22.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="160" swimtime="00:00:45.93" resultid="1357" heatid="2174" lane="5" entrytime="00:00:49.18" entrycourse="SCM" />
                <RESULT eventid="1117" points="225" swimtime="00:05:48.94" resultid="1358" heatid="2139" lane="6" entrytime="00:05:57.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                    <SPLIT distance="100" swimtime="00:01:19.23" />
                    <SPLIT distance="150" swimtime="00:02:03.17" />
                    <SPLIT distance="200" swimtime="00:02:48.22" />
                    <SPLIT distance="250" swimtime="00:03:33.78" />
                    <SPLIT distance="300" swimtime="00:04:19.12" />
                    <SPLIT distance="350" swimtime="00:05:05.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Moreira Pasqual" birthdate="2014-07-09" gender="M" nation="BRA" license="382125" swrid="5602562" athleteid="1523" externalid="382125">
              <RESULTS>
                <RESULT eventid="1083" points="97" swimtime="00:00:54.26" resultid="1524" heatid="2096" lane="8" entrytime="00:00:58.43" entrycourse="SCM" />
                <RESULT eventid="1067" points="138" swimtime="00:03:12.09" resultid="1525" heatid="2080" lane="7" entrytime="00:03:32.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.29" />
                    <SPLIT distance="100" swimtime="00:01:32.63" />
                    <SPLIT distance="150" swimtime="00:02:22.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="137" swimtime="00:00:39.08" resultid="1526" heatid="2166" lane="2" entrytime="00:00:38.83" entrycourse="SCM" />
                <RESULT eventid="1114" points="108" swimtime="00:01:43.35" resultid="1527" heatid="2135" lane="8" entrytime="00:02:12.02" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Da Cunha Souza" birthdate="2015-05-30" gender="F" nation="BRA" license="400016" swrid="5652883" athleteid="1697" externalid="400016">
              <RESULTS>
                <RESULT eventid="1080" points="84" swimtime="00:01:04.74" resultid="1698" heatid="2091" lane="3" entrytime="00:01:02.80" entrycourse="SCM" />
                <RESULT eventid="1064" points="109" swimtime="00:03:50.61" resultid="1699" heatid="2074" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.76" />
                    <SPLIT distance="100" swimtime="00:01:51.43" />
                    <SPLIT distance="150" swimtime="00:02:54.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="133" swimtime="00:00:44.85" resultid="1700" heatid="2160" lane="6" entrytime="00:00:48.76" entrycourse="SCM" />
                <RESULT eventid="1111" points="94" swimtime="00:02:04.11" resultid="1701" heatid="2128" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Jarenko Gomes" birthdate="2014-05-17" gender="F" nation="BRA" license="407692" athleteid="1808" externalid="407692">
              <RESULTS>
                <RESULT eventid="1092" points="23" swimtime="00:01:25.53" resultid="1809" heatid="2109" lane="3" />
                <RESULT eventid="1080" points="74" swimtime="00:01:07.37" resultid="1810" heatid="2090" lane="1" />
                <RESULT eventid="1136" points="56" swimtime="00:00:59.63" resultid="1811" heatid="2158" lane="6" />
                <RESULT eventid="1124" points="70" swimtime="00:01:01.03" resultid="1812" heatid="2142" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Cunha Moraes" birthdate="2012-11-26" gender="F" nation="BRA" license="406744" athleteid="1736" externalid="406744">
              <RESULTS>
                <RESULT eventid="1098" points="124" swimtime="00:00:48.87" resultid="1737" heatid="2115" lane="8" />
                <RESULT eventid="1142" points="141" swimtime="00:00:54.46" resultid="1738" heatid="2169" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Steven" lastname="Matheussi Viana E Silva" birthdate="2012-05-03" gender="M" nation="BRA" license="376986" swrid="5588810" athleteid="1494" externalid="376986">
              <RESULTS>
                <RESULT eventid="1101" points="182" swimtime="00:00:38.31" resultid="1495" heatid="2120" lane="2" entrytime="00:00:43.02" entrycourse="SCM" />
                <RESULT eventid="1073" points="207" swimtime="00:03:05.24" resultid="1496" heatid="2084" lane="4" />
                <RESULT eventid="1145" points="186" swimtime="00:00:43.66" resultid="1497" heatid="2174" lane="3" entrytime="00:00:49.19" entrycourse="SCM" />
                <RESULT eventid="1117" status="DSQ" swimtime="00:00:00.00" resultid="1498" heatid="2139" lane="7" entrytime="00:06:11.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Pens Correa" birthdate="2015-11-27" gender="M" nation="BRA" license="393262" swrid="5616449" athleteid="1643" externalid="393262">
              <RESULTS>
                <RESULT eventid="1095" points="122" swimtime="00:00:43.77" resultid="1644" heatid="2113" lane="5" entrytime="00:00:41.42" entrycourse="SCM" />
                <RESULT eventid="1067" points="138" swimtime="00:03:12.08" resultid="1645" heatid="2078" lane="8" />
                <RESULT eventid="1139" points="160" swimtime="00:00:37.13" resultid="1646" heatid="2166" lane="3" entrytime="00:00:37.64" entrycourse="SCM" />
                <RESULT eventid="1114" points="136" swimtime="00:01:35.76" resultid="1647" heatid="2133" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Cecilia" lastname="Cabrini Vieira" birthdate="2012-02-11" gender="F" nation="BRA" license="376961" swrid="5588571" athleteid="1397" externalid="376961">
              <RESULTS>
                <RESULT eventid="1098" points="262" swimtime="00:00:38.10" resultid="1398" heatid="2117" lane="3" entrytime="00:00:39.16" entrycourse="SCM" />
                <RESULT eventid="1086" points="413" swimtime="00:01:07.47" resultid="1399" heatid="2102" lane="7" entrytime="00:01:14.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="421" swimtime="00:05:08.61" resultid="1400" heatid="2125" lane="6" entrytime="00:05:47.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                    <SPLIT distance="100" swimtime="00:01:13.15" />
                    <SPLIT distance="150" swimtime="00:01:53.32" />
                    <SPLIT distance="200" swimtime="00:02:34.00" />
                    <SPLIT distance="250" swimtime="00:03:13.67" />
                    <SPLIT distance="300" swimtime="00:03:52.71" />
                    <SPLIT distance="350" swimtime="00:04:31.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="326" swimtime="00:01:19.72" resultid="1401" heatid="2152" lane="3" entrytime="00:01:22.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Marie Silva" birthdate="2014-08-24" gender="F" nation="BRA" license="391025" swrid="5602556" athleteid="1593" externalid="391025">
              <RESULTS>
                <RESULT eventid="1080" points="128" swimtime="00:00:56.29" resultid="1594" heatid="2092" lane="2" entrytime="00:00:57.39" entrycourse="SCM" />
                <RESULT eventid="1064" points="147" swimtime="00:03:28.56" resultid="1595" heatid="2075" lane="8" entrytime="00:03:59.34" entrycourse="SCM" />
                <RESULT eventid="1136" points="139" swimtime="00:00:44.23" resultid="1596" heatid="2161" lane="6" entrytime="00:00:41.68" entrycourse="SCM" />
                <RESULT eventid="1111" points="130" swimtime="00:01:51.47" resultid="1597" heatid="2131" lane="8" entrytime="00:02:13.96" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Jacob Brunetti" birthdate="2015-11-10" gender="M" nation="BRA" license="406837" swrid="5717274" athleteid="1779" externalid="406837">
              <RESULTS>
                <RESULT eventid="1083" points="27" swimtime="00:01:22.21" resultid="1780" heatid="2093" lane="2" />
                <RESULT eventid="1067" points="27" swimtime="00:05:29.32" resultid="1781" heatid="2077" lane="4" />
                <RESULT eventid="1139" points="26" swimtime="00:01:07.36" resultid="1782" heatid="2163" lane="6" entrytime="00:01:12.39" entrycourse="SCM" />
                <RESULT eventid="1127" points="38" swimtime="00:01:05.41" resultid="1783" heatid="2147" lane="8" entrytime="00:01:18.03" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Poletto Abrahao" birthdate="2014-10-20" gender="M" nation="BRA" license="382128" swrid="5602571" athleteid="1533" externalid="382128">
              <RESULTS>
                <RESULT eventid="1095" points="149" swimtime="00:00:41.02" resultid="1534" heatid="2113" lane="3" entrytime="00:00:42.97" entrycourse="SCM" />
                <RESULT eventid="1067" points="144" swimtime="00:03:09.31" resultid="1535" heatid="2080" lane="5" entrytime="00:03:06.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.90" />
                    <SPLIT distance="100" swimtime="00:01:31.35" />
                    <SPLIT distance="150" swimtime="00:02:21.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="185" swimtime="00:00:35.36" resultid="1536" heatid="2166" lane="5" entrytime="00:00:36.40" entrycourse="SCM" />
                <RESULT eventid="1114" points="151" swimtime="00:01:32.44" resultid="1537" heatid="2135" lane="3" entrytime="00:01:49.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Toscani Kim" birthdate="2015-10-02" gender="F" nation="BRA" license="397276" swrid="5641778" athleteid="1682" externalid="397276">
              <RESULTS>
                <RESULT eventid="1092" points="76" swimtime="00:00:57.48" resultid="1683" heatid="2111" lane="2" entrytime="00:00:52.60" entrycourse="SCM" />
                <RESULT eventid="1080" points="132" swimtime="00:00:55.67" resultid="1684" heatid="2091" lane="7" entrytime="00:01:04.05" entrycourse="SCM" />
                <RESULT eventid="1136" points="131" swimtime="00:00:45.08" resultid="1685" heatid="2160" lane="3" entrytime="00:00:47.18" entrycourse="SCM" />
                <RESULT eventid="1111" points="113" swimtime="00:01:56.64" resultid="1686" heatid="2130" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Cabrera Cirino Dos Santos" birthdate="2013-03-30" gender="M" nation="BRA" license="376990" swrid="5588570" athleteid="1479" externalid="376990">
              <RESULTS>
                <RESULT eventid="1101" points="105" swimtime="00:00:46.02" resultid="1480" heatid="2120" lane="6" entrytime="00:00:41.81" entrycourse="SCM" />
                <RESULT eventid="1089" points="178" swimtime="00:01:19.71" resultid="1481" heatid="2107" lane="7" entrytime="00:01:19.82" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="126" swimtime="00:01:36.20" resultid="1482" heatid="2153" lane="5" />
                <RESULT eventid="1117" points="188" swimtime="00:06:10.08" resultid="1483" heatid="2138" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.67" />
                    <SPLIT distance="100" swimtime="00:01:27.70" />
                    <SPLIT distance="150" swimtime="00:02:14.96" />
                    <SPLIT distance="200" swimtime="00:03:03.28" />
                    <SPLIT distance="250" swimtime="00:03:50.68" />
                    <SPLIT distance="300" swimtime="00:04:38.93" />
                    <SPLIT distance="350" swimtime="00:05:25.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cecilia Carvalho" birthdate="2014-10-30" gender="F" nation="BRA" license="391021" swrid="5602525" athleteid="1578" externalid="391021">
              <RESULTS>
                <RESULT eventid="1080" points="78" swimtime="00:01:06.32" resultid="1579" heatid="2090" lane="3" entrytime="00:01:13.89" entrycourse="SCM" />
                <RESULT eventid="1064" points="105" swimtime="00:03:53.76" resultid="1580" heatid="2074" lane="3" entrytime="00:04:18.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.86" />
                    <SPLIT distance="100" swimtime="00:01:47.95" />
                    <SPLIT distance="150" swimtime="00:02:53.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" status="DNS" swimtime="00:00:00.00" resultid="1581" heatid="2144" lane="5" entrytime="00:00:55.17" entrycourse="SCM" />
                <RESULT eventid="1111" status="DNS" swimtime="00:00:00.00" resultid="1582" heatid="2128" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Portes Fabiane" birthdate="2012-12-28" gender="M" nation="BRA" license="376983" swrid="5588864" athleteid="1456" externalid="376983">
              <RESULTS>
                <RESULT eventid="1089" points="78" swimtime="00:01:44.57" resultid="1457" heatid="2105" lane="7" entrytime="00:01:52.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="73" swimtime="00:00:59.61" resultid="1458" heatid="2173" lane="4" entrytime="00:01:01.07" entrycourse="SCM" />
                <RESULT eventid="1133" points="66" swimtime="00:01:59.00" resultid="1459" heatid="2156" lane="6" entrytime="00:02:11.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Livia Bittencourt" birthdate="2015-11-23" gender="F" nation="BRA" license="393260" swrid="5616446" athleteid="1633" externalid="393260">
              <RESULTS>
                <RESULT eventid="1080" points="67" swimtime="00:01:09.72" resultid="1634" heatid="2090" lane="4" entrytime="00:01:12.03" entrycourse="SCM" />
                <RESULT eventid="1064" points="71" swimtime="00:04:26.33" resultid="1635" heatid="2073" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.68" />
                    <SPLIT distance="100" swimtime="00:02:07.54" />
                    <SPLIT distance="150" swimtime="00:03:18.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="66" swimtime="00:01:02.18" resultid="1636" heatid="2142" lane="2" />
                <RESULT eventid="1111" points="73" swimtime="00:02:14.69" resultid="1637" heatid="2128" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Cury Abreu" birthdate="2013-05-17" gender="F" nation="BRA" license="376974" swrid="5588614" athleteid="1426" externalid="376974">
              <RESULTS>
                <RESULT eventid="1098" points="169" swimtime="00:00:44.09" resultid="1427" heatid="2116" lane="8" entrytime="00:00:51.81" entrycourse="SCM" />
                <RESULT eventid="1086" points="295" swimtime="00:01:15.42" resultid="1428" heatid="2101" lane="8" entrytime="00:01:31.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="235" swimtime="00:06:14.69" resultid="1429" heatid="2124" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.14" />
                    <SPLIT distance="100" swimtime="00:01:27.99" />
                    <SPLIT distance="150" swimtime="00:02:15.91" />
                    <SPLIT distance="200" swimtime="00:03:04.80" />
                    <SPLIT distance="250" swimtime="00:03:54.08" />
                    <SPLIT distance="300" swimtime="00:04:43.50" />
                    <SPLIT distance="350" swimtime="00:05:31.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="228" swimtime="00:01:29.79" resultid="1430" heatid="2151" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Prosdocimo" birthdate="2012-11-30" gender="M" nation="BRA" license="369272" swrid="5602575" athleteid="1329" externalid="369272">
              <RESULTS>
                <RESULT eventid="1101" points="185" swimtime="00:00:38.13" resultid="1330" heatid="2119" lane="5" entrytime="00:00:47.52" entrycourse="SCM" />
                <RESULT eventid="1089" points="259" swimtime="00:01:10.28" resultid="1331" heatid="2107" lane="3" entrytime="00:01:17.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="190" swimtime="00:01:23.99" resultid="1332" heatid="2157" lane="1" entrytime="00:01:30.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="275" swimtime="00:05:26.30" resultid="1333" heatid="2139" lane="5" entrytime="00:05:38.64" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.21" />
                    <SPLIT distance="100" swimtime="00:01:16.86" />
                    <SPLIT distance="150" swimtime="00:01:58.49" />
                    <SPLIT distance="200" swimtime="00:02:40.37" />
                    <SPLIT distance="250" swimtime="00:03:22.66" />
                    <SPLIT distance="300" swimtime="00:04:04.77" />
                    <SPLIT distance="350" swimtime="00:04:46.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Spadari Soso" birthdate="2012-12-28" gender="F" nation="BRA" license="377313" swrid="5588921" athleteid="1769" externalid="377313">
              <RESULTS>
                <RESULT eventid="1098" points="163" swimtime="00:00:44.62" resultid="1770" heatid="2114" lane="3" />
                <RESULT eventid="1086" points="324" swimtime="00:01:13.13" resultid="1771" heatid="2101" lane="6" entrytime="00:01:20.81" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="308" swimtime="00:05:42.49" resultid="1772" heatid="2122" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:01:23.82" />
                    <SPLIT distance="150" swimtime="00:02:08.21" />
                    <SPLIT distance="200" swimtime="00:02:52.51" />
                    <SPLIT distance="250" swimtime="00:03:37.20" />
                    <SPLIT distance="300" swimtime="00:04:18.87" />
                    <SPLIT distance="350" swimtime="00:05:00.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="261" swimtime="00:00:44.37" resultid="1773" heatid="2170" lane="4" entrytime="00:00:50.68" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Massimo" lastname="Puppi Cardoso" birthdate="2015-03-30" gender="M" nation="BRA" license="406742" swrid="5717290" athleteid="1727" externalid="406742">
              <RESULTS>
                <RESULT eventid="1083" status="DNS" swimtime="00:00:00.00" resultid="1728" heatid="2095" lane="1" entrytime="00:01:09.85" entrycourse="SCM" />
                <RESULT eventid="1067" status="DNS" swimtime="00:00:00.00" resultid="1729" heatid="2079" lane="3" />
                <RESULT eventid="1127" status="DNS" swimtime="00:00:00.00" resultid="1730" heatid="2148" lane="8" entrytime="00:01:00.99" entrycourse="SCM" />
                <RESULT eventid="1114" status="DNS" swimtime="00:00:00.00" resultid="1731" heatid="2132" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Zagonel Krempel" birthdate="2015-07-27" gender="F" nation="BRA" license="406962" swrid="5717305" athleteid="1794" externalid="406962">
              <RESULTS>
                <RESULT eventid="1080" points="53" swimtime="00:01:15.18" resultid="1795" heatid="2090" lane="6" entrytime="00:01:14.49" entrycourse="SCM" />
                <RESULT eventid="1064" points="49" swimtime="00:05:01.16" resultid="1796" heatid="2072" lane="2" />
                <RESULT eventid="1124" points="44" swimtime="00:01:11.49" resultid="1797" heatid="2143" lane="2" entrytime="00:01:11.43" entrycourse="SCM" />
                <RESULT eventid="1111" points="52" swimtime="00:02:30.90" resultid="1798" heatid="2129" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:14.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Szpak De Vasconcelos" birthdate="2012-06-29" gender="M" nation="BRA" license="369271" swrid="5588928" athleteid="1324" externalid="369271">
              <RESULTS>
                <RESULT eventid="1089" points="296" swimtime="00:01:07.21" resultid="1325" heatid="2108" lane="4" entrytime="00:01:07.57" entrycourse="SCM" />
                <RESULT eventid="1073" points="273" swimtime="00:02:48.99" resultid="1326" heatid="2086" lane="4" entrytime="00:02:53.70" entrycourse="SCM" />
                <RESULT eventid="1145" points="251" swimtime="00:00:39.52" resultid="1327" heatid="2175" lane="4" entrytime="00:00:41.33" entrycourse="SCM" />
                <RESULT eventid="1117" points="292" swimtime="00:05:19.57" resultid="1328" heatid="2139" lane="4" entrytime="00:05:30.78" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Saporiti Salvi" birthdate="2013-06-28" gender="M" nation="BRA" license="377032" swrid="5588896" athleteid="1465" externalid="377032">
              <RESULTS>
                <RESULT eventid="1101" points="157" swimtime="00:00:40.24" resultid="1466" heatid="2120" lane="1" entrytime="00:00:43.82" entrycourse="SCM" />
                <RESULT eventid="1073" status="DSQ" swimtime="00:03:10.23" resultid="1467" heatid="2086" lane="8" entrytime="00:03:19.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.84" />
                    <SPLIT distance="100" swimtime="00:01:31.54" />
                    <SPLIT distance="150" swimtime="00:02:28.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="127" swimtime="00:00:49.56" resultid="1468" heatid="2174" lane="1" entrytime="00:00:55.04" entrycourse="SCM" />
                <RESULT eventid="1117" points="181" swimtime="00:06:15.08" resultid="1469" heatid="2138" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.94" />
                    <SPLIT distance="100" swimtime="00:01:29.95" />
                    <SPLIT distance="150" swimtime="00:02:18.11" />
                    <SPLIT distance="200" swimtime="00:03:07.83" />
                    <SPLIT distance="250" swimtime="00:03:56.53" />
                    <SPLIT distance="300" swimtime="00:04:44.16" />
                    <SPLIT distance="350" swimtime="00:05:30.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Salomao" birthdate="2012-05-07" gender="M" nation="BRA" license="369261" swrid="5602581" athleteid="1294" externalid="369261">
              <RESULTS>
                <RESULT eventid="1101" points="163" swimtime="00:00:39.77" resultid="1295" heatid="2121" lane="6" entrytime="00:00:37.92" entrycourse="SCM" />
                <RESULT eventid="1089" points="244" swimtime="00:01:11.75" resultid="1296" heatid="2108" lane="2" entrytime="00:01:12.13" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="156" swimtime="00:01:29.62" resultid="1297" heatid="2155" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="260" swimtime="00:05:32.29" resultid="1298" heatid="2139" lane="3" entrytime="00:05:46.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                    <SPLIT distance="100" swimtime="00:01:18.57" />
                    <SPLIT distance="150" swimtime="00:02:00.21" />
                    <SPLIT distance="200" swimtime="00:02:41.94" />
                    <SPLIT distance="250" swimtime="00:03:24.73" />
                    <SPLIT distance="300" swimtime="00:04:07.45" />
                    <SPLIT distance="350" swimtime="00:04:51.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giuliana" lastname="Sovierzoski Ferreira" birthdate="2015-01-20" gender="F" nation="BRA" license="397168" swrid="5641776" athleteid="1672" externalid="397168">
              <RESULTS>
                <RESULT eventid="1080" points="130" swimtime="00:00:55.88" resultid="1673" heatid="2092" lane="6" entrytime="00:00:57.38" entrycourse="SCM" />
                <RESULT eventid="1064" points="58" swimtime="00:04:44.34" resultid="1674" heatid="2073" lane="8" />
                <RESULT eventid="1124" points="48" swimtime="00:01:09.29" resultid="1675" heatid="2142" lane="6" />
                <RESULT eventid="1111" points="63" swimtime="00:02:21.28" resultid="1676" heatid="2130" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:12.59" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Martina" lastname="Tallao Benke" birthdate="2012-01-02" gender="F" nation="BRA" license="376984" swrid="5588931" athleteid="1460" externalid="376984">
              <RESULTS>
                <RESULT eventid="1086" points="454" swimtime="00:01:05.38" resultid="1461" heatid="2097" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1070" points="410" swimtime="00:02:43.93" resultid="1462" heatid="2083" lane="4" entrytime="00:02:57.55" entrycourse="SCM" />
                <RESULT eventid="1104" points="462" swimtime="00:04:59.04" resultid="1463" heatid="2125" lane="4" entrytime="00:05:21.10" entrycourse="SCM" />
                <RESULT eventid="1130" points="385" swimtime="00:01:15.45" resultid="1464" heatid="2152" lane="4" entrytime="00:01:18.20" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Shwetz Clivatti" birthdate="2015-03-05" gender="M" nation="BRA" license="406963" swrid="5717297" athleteid="1799" externalid="406963">
              <RESULTS>
                <RESULT eventid="1083" points="36" swimtime="00:01:15.50" resultid="1800" heatid="2094" lane="5" entrytime="00:01:18.59" entrycourse="SCM" />
                <RESULT eventid="1139" points="34" swimtime="00:01:01.73" resultid="1801" heatid="2163" lane="5" entrytime="00:01:06.35" entrycourse="SCM" />
                <RESULT eventid="1127" points="35" swimtime="00:01:07.34" resultid="1802" heatid="2147" lane="1" entrytime="00:01:17.17" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Saber" birthdate="2014-06-04" gender="F" nation="BRA" license="392141" swrid="5602554" athleteid="1618" externalid="392141">
              <RESULTS>
                <RESULT eventid="1080" points="158" swimtime="00:00:52.37" resultid="1619" heatid="2092" lane="3" entrytime="00:00:52.71" entrycourse="SCM" />
                <RESULT eventid="1064" points="146" swimtime="00:03:29.07" resultid="1620" heatid="2075" lane="7" entrytime="00:03:48.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.39" />
                    <SPLIT distance="100" swimtime="00:01:42.35" />
                    <SPLIT distance="150" swimtime="00:02:38.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1124" points="117" swimtime="00:00:51.61" resultid="1621" heatid="2144" lane="7" entrytime="00:00:59.28" entrycourse="SCM" />
                <RESULT eventid="1111" points="128" swimtime="00:01:51.94" resultid="1622" heatid="2130" lane="4" entrytime="00:02:28.45" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Antunes Luzzi" birthdate="2014-02-14" gender="M" nation="BRA" license="391019" swrid="5602510" athleteid="1568" externalid="391019">
              <RESULTS>
                <RESULT eventid="1083" status="DNS" swimtime="00:00:00.00" resultid="1569" heatid="2095" lane="7" entrytime="00:01:08.68" entrycourse="SCM" />
                <RESULT eventid="1067" status="DNS" swimtime="00:00:00.00" resultid="1570" heatid="2078" lane="4" />
                <RESULT eventid="1139" status="DNS" swimtime="00:00:00.00" resultid="1571" heatid="2163" lane="4" entrytime="00:01:05.64" entrycourse="SCM" />
                <RESULT eventid="1114" status="DNS" swimtime="00:00:00.00" resultid="1572" heatid="2132" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Pisani Ferreira" birthdate="2012-08-06" gender="F" nation="BRA" license="376985" swrid="5588862" athleteid="1499" externalid="376985">
              <RESULTS>
                <RESULT eventid="1086" points="165" swimtime="00:01:31.52" resultid="1500" heatid="2099" lane="3" entrytime="00:01:43.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="182" swimtime="00:00:50.04" resultid="1501" heatid="2170" lane="5" entrytime="00:00:52.17" entrycourse="SCM" />
                <RESULT eventid="1130" points="136" swimtime="00:01:46.58" resultid="1502" heatid="2150" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.06" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Schmidt Wozniaki" birthdate="2012-07-07" gender="M" nation="BRA" license="376963" swrid="5588905" athleteid="1407" externalid="376963">
              <RESULTS>
                <RESULT eventid="1089" points="145" swimtime="00:01:25.24" resultid="1408" heatid="2104" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="121" swimtime="00:00:50.35" resultid="1409" heatid="2174" lane="2" entrytime="00:00:53.20" entrycourse="SCM" />
                <RESULT eventid="1133" points="89" swimtime="00:01:47.85" resultid="1410" heatid="2155" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Fortes Traub" birthdate="2012-04-26" gender="M" nation="BRA" license="369532" swrid="5588707" athleteid="1369" externalid="369532">
              <RESULTS>
                <RESULT eventid="1101" points="77" swimtime="00:00:51.01" resultid="1370" heatid="2119" lane="8" />
                <RESULT eventid="1089" points="161" swimtime="00:01:22.35" resultid="1371" heatid="2106" lane="4" entrytime="00:01:23.90" entrycourse="SCM" />
                <RESULT eventid="1133" points="107" swimtime="00:01:41.50" resultid="1372" heatid="2157" lane="8" entrytime="00:01:36.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="154" swimtime="00:06:35.74" resultid="1373" heatid="2139" lane="1" entrytime="00:06:24.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.45" />
                    <SPLIT distance="100" swimtime="00:01:33.77" />
                    <SPLIT distance="150" swimtime="00:02:24.26" />
                    <SPLIT distance="200" swimtime="00:03:15.86" />
                    <SPLIT distance="250" swimtime="00:04:07.31" />
                    <SPLIT distance="300" swimtime="00:04:58.63" />
                    <SPLIT distance="350" swimtime="00:05:49.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Taborda Ribas" birthdate="2015-12-30" gender="M" nation="BRA" license="406748" swrid="5717299" athleteid="1754" externalid="406748">
              <RESULTS>
                <RESULT eventid="1083" points="34" swimtime="00:01:16.71" resultid="1755" heatid="2094" lane="3" entrytime="00:01:21.49" entrycourse="SCM" />
                <RESULT eventid="1067" points="61" swimtime="00:04:12.41" resultid="1756" heatid="2079" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.31" />
                    <SPLIT distance="100" swimtime="00:01:58.98" />
                    <SPLIT distance="150" swimtime="00:03:04.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1127" points="40" swimtime="00:01:04.29" resultid="1757" heatid="2147" lane="7" entrytime="00:01:11.96" entrycourse="SCM" />
                <RESULT eventid="1114" points="40" swimtime="00:02:23.77" resultid="1758" heatid="2132" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Petraglia" birthdate="2012-03-28" gender="M" nation="BRA" license="369282" swrid="5602569" athleteid="1364" externalid="369282">
              <RESULTS>
                <RESULT eventid="1101" status="WDR" swimtime="00:00:00.00" resultid="1365" heatid="2118" lane="3" />
                <RESULT eventid="1089" status="WDR" swimtime="00:00:00.00" resultid="1366" heatid="2107" lane="4" entrytime="00:01:16.50" entrycourse="SCM" />
                <RESULT eventid="1145" points="199" swimtime="00:00:42.72" resultid="1367" heatid="2175" lane="6" entrytime="00:00:44.88" entrycourse="SCM" />
                <RESULT eventid="1117" points="244" swimtime="00:05:39.44" resultid="1368" heatid="2138" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                    <SPLIT distance="100" swimtime="00:01:21.11" />
                    <SPLIT distance="150" swimtime="00:02:05.48" />
                    <SPLIT distance="200" swimtime="00:02:49.70" />
                    <SPLIT distance="250" swimtime="00:03:33.63" />
                    <SPLIT distance="300" swimtime="00:04:16.80" />
                    <SPLIT distance="350" swimtime="00:04:59.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Cavalca Petraglia" birthdate="2015-08-06" gender="M" nation="BRA" license="397275" swrid="5641757" athleteid="1677" externalid="397275">
              <RESULTS>
                <RESULT eventid="1095" points="27" swimtime="00:01:11.81" resultid="1678" heatid="2113" lane="8" entrytime="00:00:55.88" entrycourse="SCM" />
                <RESULT eventid="1083" points="72" swimtime="00:00:59.91" resultid="1679" heatid="2095" lane="2" entrytime="00:01:04.65" entrycourse="SCM" />
                <RESULT eventid="1127" points="69" swimtime="00:00:53.66" resultid="1680" heatid="2148" lane="7" entrytime="00:00:58.56" entrycourse="SCM" />
                <RESULT eventid="1114" points="60" swimtime="00:02:05.67" resultid="1681" heatid="2133" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:02.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Alzamora Calado" birthdate="2013-04-26" gender="F" nation="BRA" license="376960" swrid="5588522" athleteid="1392" externalid="376960">
              <RESULTS>
                <RESULT eventid="1098" status="WDR" swimtime="00:00:00.00" resultid="1393" heatid="2116" lane="5" entrytime="00:00:43.22" entrycourse="SCM" />
                <RESULT eventid="1086" status="WDR" swimtime="00:00:00.00" resultid="1394" heatid="2101" lane="2" entrytime="00:01:21.62" entrycourse="SCM" />
                <RESULT eventid="1104" status="WDR" swimtime="00:00:00.00" resultid="1395" heatid="2124" lane="6" />
                <RESULT eventid="1142" status="WDR" swimtime="00:00:00.00" resultid="1396" heatid="2171" lane="2" entrytime="00:00:47.74" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luigi" lastname="Antoniuk Paganini" birthdate="2014-11-13" gender="M" nation="BRA" license="382127" swrid="5602509" athleteid="1528" externalid="382127">
              <RESULTS>
                <RESULT eventid="1083" points="93" swimtime="00:00:54.89" resultid="1529" heatid="2095" lane="5" entrytime="00:00:59.72" entrycourse="SCM" />
                <RESULT eventid="1067" points="122" swimtime="00:03:20.17" resultid="1530" heatid="2080" lane="2" entrytime="00:03:30.10" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.46" />
                    <SPLIT distance="100" swimtime="00:01:37.57" />
                    <SPLIT distance="150" swimtime="00:02:30.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="143" swimtime="00:00:38.53" resultid="1531" heatid="2165" lane="2" entrytime="00:00:42.83" entrycourse="SCM" />
                <RESULT eventid="1114" points="95" swimtime="00:01:47.99" resultid="1532" heatid="2135" lane="2" entrytime="00:02:00.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Betina" lastname="Vieira Pellanda" birthdate="2014-02-16" gender="F" nation="BRA" license="391041" swrid="5602589" athleteid="1608" externalid="391041">
              <RESULTS>
                <RESULT eventid="1080" points="129" swimtime="00:00:56.10" resultid="1609" heatid="2091" lane="5" entrytime="00:01:02.53" entrycourse="SCM" />
                <RESULT eventid="1064" points="147" swimtime="00:03:28.95" resultid="1610" heatid="2075" lane="2" entrytime="00:03:32.41" entrycourse="SCM" />
                <RESULT eventid="1124" points="124" swimtime="00:00:50.59" resultid="1611" heatid="2145" lane="6" entrytime="00:00:49.00" entrycourse="SCM" />
                <RESULT eventid="1111" points="136" swimtime="00:01:49.88" resultid="1612" heatid="2131" lane="7" entrytime="00:02:10.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maya" lastname="Assahida Moreria" birthdate="2014-02-24" gender="F" nation="BRA" license="391020" swrid="5602512" athleteid="1573" externalid="391020">
              <RESULTS>
                <RESULT eventid="1092" points="140" swimtime="00:00:46.86" resultid="1574" heatid="2111" lane="6" entrytime="00:00:51.30" entrycourse="SCM" />
                <RESULT eventid="1064" points="147" swimtime="00:03:28.63" resultid="1575" heatid="2075" lane="6" entrytime="00:03:27.47" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.59" />
                    <SPLIT distance="100" swimtime="00:01:38.60" />
                    <SPLIT distance="150" swimtime="00:02:35.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="168" swimtime="00:00:41.53" resultid="1576" heatid="2161" lane="7" entrytime="00:00:42.49" entrycourse="SCM" />
                <RESULT eventid="1111" points="146" swimtime="00:01:47.30" resultid="1577" heatid="2131" lane="2" entrytime="00:02:09.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Ribas Omar" birthdate="2014-11-28" gender="M" nation="BRA" license="406746" swrid="5717292" athleteid="1744" externalid="406746">
              <RESULTS>
                <RESULT eventid="1095" points="31" swimtime="00:01:08.91" resultid="1745" heatid="2112" lane="2" />
                <RESULT eventid="1083" points="55" swimtime="00:01:05.44" resultid="1746" heatid="2093" lane="5" />
                <RESULT eventid="1139" points="79" swimtime="00:00:46.80" resultid="1747" heatid="2164" lane="1" entrytime="00:00:51.97" entrycourse="SCM" />
                <RESULT eventid="1114" points="49" swimtime="00:02:14.42" resultid="1748" heatid="2133" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="De Almeida Dias" birthdate="2012-02-18" gender="F" nation="BRA" license="369262" swrid="5588638" athleteid="1299" externalid="369262">
              <RESULTS>
                <RESULT eventid="1086" points="409" swimtime="00:01:07.66" resultid="1300" heatid="2102" lane="4" entrytime="00:01:10.32" entrycourse="SCM" />
                <RESULT eventid="1070" points="351" swimtime="00:02:52.63" resultid="1301" heatid="2083" lane="3" entrytime="00:03:04.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.34" />
                    <SPLIT distance="100" swimtime="00:01:22.69" />
                    <SPLIT distance="150" swimtime="00:02:14.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="423" swimtime="00:05:08.02" resultid="1302" heatid="2123" lane="4" />
                <RESULT eventid="1130" points="343" swimtime="00:01:18.41" resultid="1303" heatid="2152" lane="5" entrytime="00:01:22.58" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Gonçalves Sperandio" birthdate="2013-05-22" gender="M" nation="BRA" license="376980" swrid="5588851" athleteid="1441" externalid="376980">
              <RESULTS>
                <RESULT eventid="1089" points="170" swimtime="00:01:20.90" resultid="1442" heatid="2107" lane="2" entrytime="00:01:19.49" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1073" points="167" swimtime="00:03:18.72" resultid="1443" heatid="2086" lane="7" entrytime="00:03:17.37" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.36" />
                    <SPLIT distance="100" swimtime="00:01:39.01" />
                    <SPLIT distance="150" swimtime="00:02:36.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="133" swimtime="00:00:48.78" resultid="1444" heatid="2174" lane="6" entrytime="00:00:51.03" entrycourse="SCM" />
                <RESULT eventid="1117" points="193" swimtime="00:06:06.71" resultid="1445" heatid="2138" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.94" />
                    <SPLIT distance="100" swimtime="00:01:26.36" />
                    <SPLIT distance="150" swimtime="00:02:12.94" />
                    <SPLIT distance="200" swimtime="00:03:00.51" />
                    <SPLIT distance="250" swimtime="00:03:47.33" />
                    <SPLIT distance="300" swimtime="00:04:34.78" />
                    <SPLIT distance="350" swimtime="00:05:22.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Clara Prado Biscaia" birthdate="2013-10-24" gender="F" nation="BRA" license="391015" swrid="5602526" athleteid="1558" externalid="391015">
              <RESULTS>
                <RESULT eventid="1098" points="167" swimtime="00:00:44.20" resultid="1559" heatid="2115" lane="4" entrytime="00:00:51.97" entrycourse="SCM" />
                <RESULT eventid="1070" points="148" swimtime="00:03:50.12" resultid="1560" heatid="2082" lane="8" entrytime="00:04:08.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.08" />
                    <SPLIT distance="100" swimtime="00:01:51.11" />
                    <SPLIT distance="150" swimtime="00:02:58.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="161" swimtime="00:07:04.52" resultid="1561" heatid="2124" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.58" />
                    <SPLIT distance="100" swimtime="00:01:39.78" />
                    <SPLIT distance="150" swimtime="00:02:33.33" />
                    <SPLIT distance="200" swimtime="00:03:26.63" />
                    <SPLIT distance="250" swimtime="00:04:22.28" />
                    <SPLIT distance="300" swimtime="00:05:16.53" />
                    <SPLIT distance="350" swimtime="00:06:11.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1142" points="114" swimtime="00:00:58.39" resultid="1562" heatid="2169" lane="4" entrytime="00:01:10.37" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Bernardi Pedrosa" birthdate="2013-03-09" gender="F" nation="BRA" license="376977" swrid="5588551" athleteid="1436" externalid="376977">
              <RESULTS>
                <RESULT eventid="1086" points="190" swimtime="00:01:27.32" resultid="1437" heatid="2100" lane="7" entrytime="00:01:37.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1070" points="202" swimtime="00:03:27.68" resultid="1438" heatid="2081" lane="4" entrytime="00:04:14.10" entrycourse="SCM" />
                <RESULT eventid="1104" points="195" swimtime="00:06:38.71" resultid="1439" heatid="2123" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.09" />
                    <SPLIT distance="100" swimtime="00:01:37.41" />
                    <SPLIT distance="150" swimtime="00:02:27.73" />
                    <SPLIT distance="200" swimtime="00:03:19.57" />
                    <SPLIT distance="250" swimtime="00:04:10.54" />
                    <SPLIT distance="300" swimtime="00:05:01.78" />
                    <SPLIT distance="350" swimtime="00:05:52.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1130" points="180" swimtime="00:01:37.16" resultid="1440" heatid="2150" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Baptistella" birthdate="2013-01-23" gender="M" nation="BRA" license="391152" swrid="5602545" athleteid="1613" externalid="391152">
              <RESULTS>
                <RESULT eventid="1089" points="155" swimtime="00:01:23.45" resultid="1614" heatid="2107" lane="8" entrytime="00:01:22.99" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1073" points="149" swimtime="00:03:26.36" resultid="1615" heatid="2085" lane="1" entrytime="00:03:54.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.58" />
                    <SPLIT distance="100" swimtime="00:01:37.50" />
                    <SPLIT distance="150" swimtime="00:02:37.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="153" swimtime="00:01:30.19" resultid="1616" heatid="2153" lane="4" />
                <RESULT eventid="1117" points="182" swimtime="00:06:14.19" resultid="1617" heatid="2138" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                    <SPLIT distance="100" swimtime="00:01:23.37" />
                    <SPLIT distance="150" swimtime="00:02:12.21" />
                    <SPLIT distance="200" swimtime="00:03:02.39" />
                    <SPLIT distance="250" swimtime="00:03:51.96" />
                    <SPLIT distance="300" swimtime="00:04:41.11" />
                    <SPLIT distance="350" swimtime="00:05:30.34" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Cipriani Presiazniuk" birthdate="2012-07-03" gender="M" nation="BRA" license="369267" swrid="5588594" athleteid="1309" externalid="369267">
              <RESULTS>
                <RESULT eventid="1089" points="241" swimtime="00:01:12.05" resultid="1310" heatid="2108" lane="1" entrytime="00:01:13.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1073" points="204" swimtime="00:03:06.22" resultid="1311" heatid="2086" lane="2" entrytime="00:03:17.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.54" />
                    <SPLIT distance="100" swimtime="00:01:28.96" />
                    <SPLIT distance="150" swimtime="00:02:29.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1133" points="172" swimtime="00:01:26.78" resultid="1312" heatid="2157" lane="3" entrytime="00:01:25.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1117" points="230" swimtime="00:05:46.30" resultid="1313" heatid="2139" lane="2" entrytime="00:06:04.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                    <SPLIT distance="100" swimtime="00:01:21.15" />
                    <SPLIT distance="150" swimtime="00:02:05.42" />
                    <SPLIT distance="200" swimtime="00:02:50.89" />
                    <SPLIT distance="250" swimtime="00:03:35.06" />
                    <SPLIT distance="300" swimtime="00:04:19.20" />
                    <SPLIT distance="350" swimtime="00:05:03.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Elisa" lastname="Osternack Almeida" birthdate="2015-04-14" gender="F" nation="BRA" license="406747" swrid="5717286" athleteid="1749" externalid="406747">
              <RESULTS>
                <RESULT eventid="1092" points="65" swimtime="00:01:00.55" resultid="1750" heatid="2110" lane="7" entrytime="00:01:07.04" entrycourse="SCM" />
                <RESULT eventid="1064" points="72" swimtime="00:04:25.09" resultid="1751" heatid="2072" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.99" />
                    <SPLIT distance="100" swimtime="00:02:01.16" />
                    <SPLIT distance="150" swimtime="00:03:15.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1136" points="115" swimtime="00:00:47.03" resultid="1752" heatid="2159" lane="6" entrytime="00:00:55.82" entrycourse="SCM" />
                <RESULT eventid="1111" points="95" swimtime="00:02:03.47" resultid="1753" heatid="2130" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Puppi Cardoso" birthdate="2015-03-30" gender="F" nation="BRA" license="406741" swrid="5717289" athleteid="1722" externalid="406741">
              <RESULTS>
                <RESULT eventid="1092" status="DNS" swimtime="00:00:00.00" resultid="1723" heatid="2109" lane="4" entrytime="00:01:11.34" entrycourse="SCM" />
                <RESULT eventid="1064" status="DNS" swimtime="00:00:00.00" resultid="1724" heatid="2072" lane="6" />
                <RESULT eventid="1124" points="75" swimtime="00:00:59.70" resultid="1725" heatid="2144" lane="3" entrytime="00:00:56.23" entrycourse="SCM" />
                <RESULT eventid="1111" points="67" swimtime="00:02:19.08" resultid="1726" heatid="2129" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:04.94" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Hallage Papp" birthdate="2012-07-02" gender="M" nation="BRA" license="377042" swrid="5588736" athleteid="1475" externalid="377042">
              <RESULTS>
                <RESULT eventid="1089" points="184" swimtime="00:01:18.79" resultid="1476" heatid="2106" lane="8" entrytime="00:01:35.24" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="111" swimtime="00:00:51.88" resultid="1477" heatid="2174" lane="7" entrytime="00:00:53.31" entrycourse="SCM" />
                <RESULT eventid="1133" points="132" swimtime="00:01:34.83" resultid="1478" heatid="2155" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.05" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Liam" lastname="Batista Grise" birthdate="2014-03-27" gender="M" nation="BRA" license="391008" swrid="5602514" athleteid="1548" externalid="391008">
              <RESULTS>
                <RESULT eventid="1083" points="76" swimtime="00:00:58.76" resultid="1549" heatid="2095" lane="3" entrytime="00:01:01.90" entrycourse="SCM" />
                <RESULT eventid="1067" points="34" swimtime="00:05:05.37" resultid="1550" heatid="2076" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:00.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1139" points="89" swimtime="00:00:45.04" resultid="1551" heatid="2165" lane="6" entrytime="00:00:42.24" entrycourse="SCM" />
                <RESULT eventid="1114" points="54" swimtime="00:02:10.30" resultid="1552" heatid="2134" lane="5" entrytime="00:02:30.50" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:06.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Antunes Saboia" birthdate="2012-06-28" gender="M" nation="BRA" license="369278" swrid="5602511" athleteid="1349" externalid="369278">
              <RESULTS>
                <RESULT eventid="1089" points="239" swimtime="00:01:12.24" resultid="1350" heatid="2108" lane="8" entrytime="00:01:14.54" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1073" points="232" swimtime="00:02:58.33" resultid="1351" heatid="2086" lane="6" entrytime="00:03:16.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.11" />
                    <SPLIT distance="100" swimtime="00:01:29.21" />
                    <SPLIT distance="150" swimtime="00:02:20.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1145" points="238" swimtime="00:00:40.22" resultid="1352" heatid="2175" lane="3" entrytime="00:00:44.79" entrycourse="SCM" />
                <RESULT eventid="1133" points="169" swimtime="00:01:27.35" resultid="1353" heatid="2157" lane="7" entrytime="00:01:30.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16131" nation="BRA" region="PR" clubid="1813" swrid="93766" name="Associação Nadar Colombo" shortname="Equipe Nadar">
          <ATHLETES>
            <ATHLETE firstname="Gabriela" lastname="Poli" birthdate="2014-02-27" gender="F" nation="BRA" license="408670" athleteid="1817" externalid="408670">
              <RESULTS>
                <RESULT eventid="1136" points="37" swimtime="00:01:08.80" resultid="1818" heatid="2158" lane="5" />
                <RESULT eventid="1124" points="40" swimtime="00:01:13.79" resultid="1819" heatid="2143" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tayna" lastname="Macedo Gabardo" birthdate="2012-12-01" gender="F" nation="BRA" license="406704" swrid="5717281" athleteid="1814" externalid="406704">
              <RESULTS>
                <RESULT eventid="1098" points="142" swimtime="00:00:46.69" resultid="1815" heatid="2114" lane="6" />
                <RESULT eventid="1086" points="232" swimtime="00:01:21.68" resultid="1816" heatid="2098" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jackson" lastname="Luiz Neto" birthdate="2016-08-18" gender="M" nation="BRA" license="408672" athleteid="1822" externalid="408672">
              <RESULTS>
                <RESULT eventid="1122" points="56" swimtime="00:00:52.48" resultid="1823" heatid="2141" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Weinert Jardwski" birthdate="2013-12-13" gender="F" nation="BRA" license="408671" athleteid="1820" externalid="408671">
              <RESULTS>
                <RESULT eventid="1130" status="DSQ" swimtime="00:02:14.50" resultid="1821" heatid="2150" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:01:01.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
