<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.80168">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Curitiba" name="Troféu Alexandre Viscardi (Infantil/Sênior) 2024" course="LCM" deadline="2024-09-14" entrystartdate="2024-09-09" entrytype="INVITATION" hostclub="Clube Curitibano" hostclub.url="https://clubecuritibano.com.br/" number="38319" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/newInterface/eventos/38319" startmethod="1" timing="AUTOMATIC" touchpad="BOTHSIDE" masters="F" withdrawuntil="2024-09-16" state="PR" nation="BRA" hytek.courseorder="L">
      <AGEDATE value="2024-01-01" type="YEAR" />
      <POOL name="Parque Aquático do Clube Curitibano" lanemin="1" lanemax="8" />
      <FACILITY city="Curitiba" name="Parque Aquático do Clube Curitibano" nation="BRA" state="PR" street="Avenida Presidente Getúlio Vargas, 2857" street2="Água Verde" zip="80240-040" />
      <POINTTABLE pointtableid="3017" name="AQUA Point Scoring" version="2024" />
      <QUALIFY from="2023-09-20" until="2024-09-18" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99252-0598" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99252-0598" street="Avenida do Batel, 1230" street2="Sala 202" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-09-19" daytime="09:10" endtime="12:40" number="1" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1064" daytime="09:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1065" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3850" />
                    <RANKING order="2" place="2" resultid="3331" />
                    <RANKING order="3" place="3" resultid="3338" />
                    <RANKING order="4" place="4" resultid="3796" />
                    <RANKING order="5" place="5" resultid="3745" />
                    <RANKING order="6" place="6" resultid="3778" />
                    <RANKING order="7" place="7" resultid="3930" />
                    <RANKING order="8" place="8" resultid="3408" />
                    <RANKING order="9" place="9" resultid="4112" />
                    <RANKING order="10" place="10" resultid="3758" />
                    <RANKING order="11" place="11" resultid="4624" />
                    <RANKING order="12" place="12" resultid="3121" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1067" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3697" />
                    <RANKING order="2" place="2" resultid="3659" />
                    <RANKING order="3" place="3" resultid="2414" />
                    <RANKING order="4" place="4" resultid="3970" />
                    <RANKING order="5" place="5" resultid="4545" />
                    <RANKING order="6" place="6" resultid="3381" />
                    <RANKING order="7" place="7" resultid="3652" />
                    <RANKING order="8" place="8" resultid="3685" />
                    <RANKING order="9" place="9" resultid="3135" />
                    <RANKING order="10" place="10" resultid="4316" />
                    <RANKING order="11" place="11" resultid="4580" />
                    <RANKING order="12" place="12" resultid="3275" />
                    <RANKING order="13" place="13" resultid="4645" />
                    <RANKING order="14" place="14" resultid="2702" />
                    <RANKING order="15" place="15" resultid="4357" />
                    <RANKING order="16" place="16" resultid="4350" />
                    <RANKING order="17" place="17" resultid="4079" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4419" />
                    <RANKING order="2" place="2" resultid="3524" />
                    <RANKING order="3" place="3" resultid="3462" />
                    <RANKING order="4" place="4" resultid="4506" />
                    <RANKING order="5" place="5" resultid="3229" />
                    <RANKING order="6" place="6" resultid="4067" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5821" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3037" />
                    <RANKING order="2" place="2" resultid="2865" />
                    <RANKING order="3" place="3" resultid="2795" />
                    <RANKING order="4" place="4" resultid="4339" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5822" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3546" />
                    <RANKING order="2" place="2" resultid="3514" />
                    <RANKING order="3" place="3" resultid="4192" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5823" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2773" />
                    <RANKING order="2" place="2" resultid="4433" />
                    <RANKING order="3" place="3" resultid="4305" />
                    <RANKING order="4" place="4" resultid="4055" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5824" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3903" />
                    <RANKING order="2" place="2" resultid="3915" />
                    <RANKING order="3" place="3" resultid="4280" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5825" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3903" />
                    <RANKING order="2" place="2" resultid="4419" />
                    <RANKING order="3" place="3" resultid="3915" />
                    <RANKING order="4" place="4" resultid="3524" />
                    <RANKING order="5" place="5" resultid="3462" />
                    <RANKING order="6" place="6" resultid="3546" />
                    <RANKING order="7" place="7" resultid="3514" />
                    <RANKING order="8" place="8" resultid="3850" />
                    <RANKING order="9" place="9" resultid="2773" />
                    <RANKING order="10" place="10" resultid="3697" />
                    <RANKING order="11" place="11" resultid="4433" />
                    <RANKING order="12" place="12" resultid="3659" />
                    <RANKING order="13" place="13" resultid="2414" />
                    <RANKING order="14" place="14" resultid="3331" />
                    <RANKING order="15" place="15" resultid="3338" />
                    <RANKING order="16" place="16" resultid="3796" />
                    <RANKING order="17" place="17" resultid="3970" />
                    <RANKING order="18" place="18" resultid="3745" />
                    <RANKING order="19" place="19" resultid="4545" />
                    <RANKING order="20" place="20" resultid="3381" />
                    <RANKING order="21" place="21" resultid="3037" />
                    <RANKING order="22" place="22" resultid="3652" />
                    <RANKING order="23" place="23" resultid="3778" />
                    <RANKING order="24" place="24" resultid="3685" />
                    <RANKING order="25" place="25" resultid="3135" />
                    <RANKING order="26" place="26" resultid="4192" />
                    <RANKING order="27" place="27" resultid="2865" />
                    <RANKING order="28" place="28" resultid="2795" />
                    <RANKING order="29" place="29" resultid="4316" />
                    <RANKING order="30" place="30" resultid="3930" />
                    <RANKING order="31" place="31" resultid="3408" />
                    <RANKING order="32" place="32" resultid="4580" />
                    <RANKING order="33" place="33" resultid="3275" />
                    <RANKING order="34" place="34" resultid="4339" />
                    <RANKING order="35" place="35" resultid="4506" />
                    <RANKING order="36" place="36" resultid="4112" />
                    <RANKING order="37" place="37" resultid="3758" />
                    <RANKING order="38" place="38" resultid="4305" />
                    <RANKING order="39" place="39" resultid="4280" />
                    <RANKING order="40" place="40" resultid="4645" />
                    <RANKING order="41" place="41" resultid="2702" />
                    <RANKING order="42" place="42" resultid="3229" />
                    <RANKING order="43" place="43" resultid="4624" />
                    <RANKING order="44" place="44" resultid="4055" />
                    <RANKING order="45" place="45" resultid="4357" />
                    <RANKING order="46" place="46" resultid="4067" />
                    <RANKING order="47" place="47" resultid="3121" />
                    <RANKING order="48" place="48" resultid="4350" />
                    <RANKING order="49" place="49" resultid="4079" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5048" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5049" daytime="09:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5050" daytime="09:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5051" daytime="09:32" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5052" daytime="09:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5053" daytime="09:46" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5054" daytime="09:54" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5055" daytime="10:00" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1072" daytime="10:08" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6182" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3310" />
                    <RANKING order="2" place="2" resultid="3826" />
                    <RANKING order="3" place="3" resultid="3324" />
                    <RANKING order="4" place="4" resultid="3728" />
                    <RANKING order="5" place="5" resultid="3741" />
                    <RANKING order="6" place="6" resultid="3721" />
                    <RANKING order="7" place="7" resultid="4559" />
                    <RANKING order="8" place="8" resultid="4343" />
                    <RANKING order="9" place="9" resultid="4385" />
                    <RANKING order="10" place="10" resultid="3764" />
                    <RANKING order="11" place="11" resultid="3790" />
                    <RANKING order="12" place="12" resultid="4573" />
                    <RANKING order="13" place="13" resultid="3874" />
                    <RANKING order="14" place="14" resultid="4140" />
                    <RANKING order="15" place="15" resultid="4535" />
                    <RANKING order="16" place="16" resultid="3221" />
                    <RANKING order="17" place="17" resultid="4098" />
                    <RANKING order="18" place="18" resultid="2839" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6183" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3665" />
                    <RANKING order="2" place="2" resultid="3289" />
                    <RANKING order="3" place="3" resultid="3678" />
                    <RANKING order="4" place="4" resultid="3815" />
                    <RANKING order="5" place="5" resultid="3387" />
                    <RANKING order="6" place="6" resultid="4652" />
                    <RANKING order="7" place="7" resultid="4527" />
                    <RANKING order="8" place="8" resultid="4593" />
                    <RANKING order="9" place="9" resultid="3704" />
                    <RANKING order="10" place="10" resultid="4269" />
                    <RANKING order="11" place="11" resultid="3296" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6184" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3540" />
                    <RANKING order="2" place="2" resultid="3268" />
                    <RANKING order="3" place="3" resultid="3617" />
                    <RANKING order="4" place="4" resultid="4255" />
                    <RANKING order="5" place="5" resultid="3589" />
                    <RANKING order="6" place="6" resultid="4032" />
                    <RANKING order="7" place="7" resultid="2488" />
                    <RANKING order="8" place="8" resultid="4631" />
                    <RANKING order="9" place="9" resultid="3209" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6185" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3256" />
                    <RANKING order="2" place="2" resultid="3821" />
                    <RANKING order="3" place="3" resultid="3486" />
                    <RANKING order="4" place="4" resultid="3087" />
                    <RANKING order="5" place="5" resultid="3394" />
                    <RANKING order="6" place="6" resultid="3623" />
                    <RANKING order="7" place="7" resultid="4440" />
                    <RANKING order="8" place="8" resultid="4475" />
                    <RANKING order="9" place="9" resultid="3107" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6186" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3518" />
                    <RANKING order="2" place="2" resultid="3552" />
                    <RANKING order="3" place="3" resultid="4426" />
                    <RANKING order="4" place="4" resultid="4365" />
                    <RANKING order="5" place="5" resultid="3094" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6187" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3959" />
                    <RANKING order="2" place="2" resultid="3715" />
                    <RANKING order="3" place="3" resultid="3066" />
                    <RANKING order="4" place="4" resultid="3243" />
                    <RANKING order="5" place="5" resultid="4552" />
                    <RANKING order="6" place="6" resultid="3080" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6188" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4328" />
                    <RANKING order="2" place="2" resultid="2903" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6189" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3518" />
                    <RANKING order="2" place="2" resultid="3959" />
                    <RANKING order="3" place="3" resultid="3552" />
                    <RANKING order="4" place="4" resultid="3256" />
                    <RANKING order="5" place="5" resultid="3821" />
                    <RANKING order="6" place="6" resultid="3540" />
                    <RANKING order="7" place="7" resultid="4426" />
                    <RANKING order="8" place="8" resultid="3268" />
                    <RANKING order="9" place="9" resultid="3486" />
                    <RANKING order="10" place="10" resultid="3715" />
                    <RANKING order="11" place="11" resultid="3665" />
                    <RANKING order="12" place="12" resultid="3087" />
                    <RANKING order="13" place="13" resultid="3617" />
                    <RANKING order="14" place="14" resultid="3394" />
                    <RANKING order="15" place="15" resultid="3289" />
                    <RANKING order="16" place="16" resultid="4255" />
                    <RANKING order="17" place="17" resultid="3066" />
                    <RANKING order="18" place="18" resultid="3678" />
                    <RANKING order="19" place="19" resultid="3243" />
                    <RANKING order="20" place="20" resultid="3310" />
                    <RANKING order="21" place="21" resultid="3623" />
                    <RANKING order="22" place="22" resultid="3815" />
                    <RANKING order="23" place="23" resultid="4552" />
                    <RANKING order="24" place="24" resultid="3826" />
                    <RANKING order="25" place="25" resultid="3589" />
                    <RANKING order="26" place="26" resultid="3387" />
                    <RANKING order="27" place="27" resultid="4365" />
                    <RANKING order="28" place="28" resultid="3080" />
                    <RANKING order="29" place="29" resultid="4328" />
                    <RANKING order="30" place="30" resultid="4440" />
                    <RANKING order="31" place="31" resultid="4475" />
                    <RANKING order="32" place="32" resultid="3107" />
                    <RANKING order="33" place="33" resultid="3324" />
                    <RANKING order="34" place="34" resultid="4652" />
                    <RANKING order="35" place="35" resultid="3728" />
                    <RANKING order="36" place="36" resultid="4527" />
                    <RANKING order="37" place="37" resultid="3741" />
                    <RANKING order="38" place="38" resultid="4593" />
                    <RANKING order="39" place="39" resultid="4032" />
                    <RANKING order="40" place="40" resultid="2903" />
                    <RANKING order="41" place="41" resultid="3721" />
                    <RANKING order="42" place="42" resultid="4559" />
                    <RANKING order="43" place="43" resultid="4343" />
                    <RANKING order="44" place="44" resultid="2488" />
                    <RANKING order="45" place="45" resultid="3704" />
                    <RANKING order="46" place="46" resultid="4385" />
                    <RANKING order="47" place="47" resultid="3764" />
                    <RANKING order="48" place="48" resultid="4269" />
                    <RANKING order="49" place="49" resultid="3296" />
                    <RANKING order="50" place="50" resultid="3790" />
                    <RANKING order="51" place="51" resultid="3094" />
                    <RANKING order="52" place="52" resultid="4573" />
                    <RANKING order="53" place="53" resultid="4631" />
                    <RANKING order="54" place="54" resultid="3874" />
                    <RANKING order="55" place="55" resultid="4140" />
                    <RANKING order="56" place="56" resultid="4535" />
                    <RANKING order="57" place="57" resultid="3221" />
                    <RANKING order="58" place="58" resultid="4098" />
                    <RANKING order="59" place="59" resultid="3209" />
                    <RANKING order="60" place="60" resultid="2839" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5056" daytime="10:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5057" daytime="10:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5058" daytime="10:22" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5059" daytime="10:28" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5060" daytime="10:34" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5061" daytime="10:42" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5062" daytime="10:48" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5063" daytime="10:54" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5064" daytime="11:02" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1080" daytime="11:08" gender="F" number="3" order="3" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5834" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3744" />
                    <RANKING order="2" place="2" resultid="3771" />
                    <RANKING order="3" place="3" resultid="3929" />
                    <RANKING order="4" place="4" resultid="3373" />
                    <RANKING order="5" place="5" resultid="4566" />
                    <RANKING order="6" place="6" resultid="4168" />
                    <RANKING order="7" place="7" resultid="3422" />
                    <RANKING order="8" place="8" resultid="4513" />
                    <RANKING order="9" place="9" resultid="2669" />
                    <RANKING order="10" place="10" resultid="3757" />
                    <RANKING order="11" place="11" resultid="4070" />
                    <RANKING order="12" place="12" resultid="4175" />
                    <RANKING order="13" place="13" resultid="2719" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5835" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4262" />
                    <RANKING order="2" place="2" resultid="3529" />
                    <RANKING order="3" place="3" resultid="4579" />
                    <RANKING order="4" place="4" resultid="3380" />
                    <RANKING order="5" place="5" resultid="4586" />
                    <RANKING order="6" place="6" resultid="2637" />
                    <RANKING order="7" place="7" resultid="4212" />
                    <RANKING order="8" place="8" resultid="3833" />
                    <RANKING order="9" place="9" resultid="2701" />
                    <RANKING order="10" place="10" resultid="4078" />
                    <RANKING order="11" place="-1" resultid="3885" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5836" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3593" />
                    <RANKING order="2" place="2" resultid="2942" />
                    <RANKING order="3" place="3" resultid="3535" />
                    <RANKING order="4" place="4" resultid="3598" />
                    <RANKING order="5" place="5" resultid="2477" />
                    <RANKING order="6" place="6" resultid="3282" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5837" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3458" />
                    <RANKING order="2" place="2" resultid="3467" />
                    <RANKING order="3" place="3" resultid="3846" />
                    <RANKING order="4" place="4" resultid="3317" />
                    <RANKING order="5" place="5" resultid="2585" />
                    <RANKING order="6" place="6" resultid="2713" />
                    <RANKING order="7" place="7" resultid="2407" />
                    <RANKING order="8" place="8" resultid="4447" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5838" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3513" />
                    <RANKING order="2" place="2" resultid="2963" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5839" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3952" />
                    <RANKING order="2" place="2" resultid="2459" />
                    <RANKING order="3" place="3" resultid="4239" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5840" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4028" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5065" daytime="11:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5066" daytime="11:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5067" daytime="11:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5068" daytime="11:18" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5069" daytime="11:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5070" daytime="11:22" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1088" daytime="11:26" gender="M" number="4" order="4" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5866" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3734" />
                    <RANKING order="2" place="2" resultid="3784" />
                    <RANKING order="3" place="3" resultid="2624" />
                    <RANKING order="4" place="4" resultid="3415" />
                    <RANKING order="5" place="5" resultid="4384" />
                    <RANKING order="6" place="6" resultid="3345" />
                    <RANKING order="7" place="7" resultid="2501" />
                    <RANKING order="8" place="8" resultid="3862" />
                    <RANKING order="9" place="9" resultid="3366" />
                    <RANKING order="10" place="10" resultid="2556" />
                    <RANKING order="11" place="11" resultid="3401" />
                    <RANKING order="12" place="12" resultid="4534" />
                    <RANKING order="13" place="13" resultid="3802" />
                    <RANKING order="14" place="14" resultid="3202" />
                    <RANKING order="15" place="15" resultid="2806" />
                    <RANKING order="16" place="16" resultid="2428" />
                    <RANKING order="17" place="17" resultid="4133" />
                    <RANKING order="18" place="18" resultid="3751" />
                    <RANKING order="19" place="19" resultid="2853" />
                    <RANKING order="20" place="20" resultid="4105" />
                    <RANKING order="21" place="21" resultid="2846" />
                    <RANKING order="22" place="22" resultid="4205" />
                    <RANKING order="23" place="-1" resultid="4540" />
                    <RANKING order="24" place="-1" resultid="4619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5867" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4161" />
                    <RANKING order="2" place="2" resultid="4268" />
                    <RANKING order="3" place="3" resultid="3010" />
                    <RANKING order="4" place="4" resultid="4659" />
                    <RANKING order="5" place="5" resultid="2952" />
                    <RANKING order="6" place="6" resultid="2981" />
                    <RANKING order="7" place="7" resultid="3634" />
                    <RANKING order="8" place="8" resultid="4074" />
                    <RANKING order="9" place="9" resultid="3021" />
                    <RANKING order="10" place="-1" resultid="3691" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5868" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2449" />
                    <RANKING order="2" place="2" resultid="4298" />
                    <RANKING order="3" place="3" resultid="3603" />
                    <RANKING order="4" place="4" resultid="4600" />
                    <RANKING order="5" place="5" resultid="2545" />
                    <RANKING order="6" place="6" resultid="2915" />
                    <RANKING order="7" place="7" resultid="4489" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5869" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3507" />
                    <RANKING order="2" place="2" resultid="2601" />
                    <RANKING order="3" place="3" resultid="3857" />
                    <RANKING order="4" place="4" resultid="3492" />
                    <RANKING order="5" place="5" resultid="3868" />
                    <RANKING order="6" place="6" resultid="4396" />
                    <RANKING order="7" place="7" resultid="3359" />
                    <RANKING order="8" place="8" resultid="4311" />
                    <RANKING order="9" place="9" resultid="4147" />
                    <RANKING order="10" place="10" resultid="2550" />
                    <RANKING order="11" place="11" resultid="2663" />
                    <RANKING order="12" place="12" resultid="3114" />
                    <RANKING order="13" place="13" resultid="4275" />
                    <RANKING order="14" place="-1" resultid="4052" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5870" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2400" />
                    <RANKING order="2" place="2" resultid="3558" />
                    <RANKING order="3" place="3" resultid="3517" />
                    <RANKING order="4" place="4" resultid="3303" />
                    <RANKING order="5" place="5" resultid="4182" />
                    <RANKING order="6" place="6" resultid="4403" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5871" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2573" />
                    <RANKING order="2" place="2" resultid="2886" />
                    <RANKING order="3" place="3" resultid="2813" />
                    <RANKING order="4" place="4" resultid="3242" />
                    <RANKING order="5" place="5" resultid="4234" />
                    <RANKING order="6" place="6" resultid="3191" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5872" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2456" />
                    <RANKING order="2" place="2" resultid="2562" />
                    <RANKING order="3" place="-1" resultid="2907" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5078" daytime="11:26" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5079" daytime="11:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5080" daytime="11:32" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5081" daytime="11:36" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5082" daytime="11:38" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5083" daytime="11:40" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5084" daytime="11:44" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5085" daytime="11:46" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5086" daytime="11:48" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5087" daytime="11:52" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1096" daytime="11:54" gender="F" number="5" order="5" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5873" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4169" />
                    <RANKING order="2" place="2" resultid="2657" />
                    <RANKING order="3" place="3" resultid="3779" />
                    <RANKING order="4" place="4" resultid="4047" />
                    <RANKING order="5" place="5" resultid="4113" />
                    <RANKING order="6" place="6" resultid="3922" />
                    <RANKING order="7" place="7" resultid="3772" />
                    <RANKING order="8" place="8" resultid="3839" />
                    <RANKING order="9" place="9" resultid="3197" />
                    <RANKING order="10" place="10" resultid="3000" />
                    <RANKING order="11" place="11" resultid="2630" />
                    <RANKING order="12" place="12" resultid="4514" />
                    <RANKING order="13" place="13" resultid="4243" />
                    <RANKING order="14" place="14" resultid="4176" />
                    <RANKING order="15" place="15" resultid="2738" />
                    <RANKING order="16" place="16" resultid="4625" />
                    <RANKING order="17" place="17" resultid="2761" />
                    <RANKING order="18" place="18" resultid="2720" />
                    <RANKING order="19" place="19" resultid="3122" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5874" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2421" />
                    <RANKING order="2" place="2" resultid="3646" />
                    <RANKING order="3" place="2" resultid="3971" />
                    <RANKING order="4" place="4" resultid="2725" />
                    <RANKING order="5" place="5" resultid="2644" />
                    <RANKING order="6" place="6" resultid="3653" />
                    <RANKING order="7" place="7" resultid="3429" />
                    <RANKING order="8" place="8" resultid="3660" />
                    <RANKING order="9" place="9" resultid="4546" />
                    <RANKING order="10" place="9" resultid="4638" />
                    <RANKING order="11" place="11" resultid="3156" />
                    <RANKING order="12" place="12" resultid="4317" />
                    <RANKING order="13" place="13" resultid="3233" />
                    <RANKING order="14" place="14" resultid="3640" />
                    <RANKING order="15" place="15" resultid="2825" />
                    <RANKING order="16" place="16" resultid="3834" />
                    <RANKING order="17" place="17" resultid="4213" />
                    <RANKING order="18" place="18" resultid="2506" />
                    <RANKING order="19" place="19" resultid="4358" />
                    <RANKING order="20" place="20" resultid="2750" />
                    <RANKING order="21" place="21" resultid="4351" />
                    <RANKING order="22" place="-1" resultid="2517" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5875" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3474" />
                    <RANKING order="2" place="2" resultid="4420" />
                    <RANKING order="3" place="3" resultid="2464" />
                    <RANKING order="4" place="4" resultid="2818" />
                    <RANKING order="5" place="5" resultid="3608" />
                    <RANKING order="6" place="6" resultid="2947" />
                    <RANKING order="7" place="7" resultid="4154" />
                    <RANKING order="8" place="8" resultid="4468" />
                    <RANKING order="9" place="8" resultid="4482" />
                    <RANKING order="10" place="10" resultid="3100" />
                    <RANKING order="11" place="11" resultid="3187" />
                    <RANKING order="12" place="12" resultid="4507" />
                    <RANKING order="13" place="13" resultid="4379" />
                    <RANKING order="14" place="14" resultid="2596" />
                    <RANKING order="15" place="15" resultid="2591" />
                    <RANKING order="16" place="16" resultid="3230" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5876" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4372" />
                    <RANKING order="2" place="2" resultid="3468" />
                    <RANKING order="3" place="3" resultid="2707" />
                    <RANKING order="4" place="4" resultid="2586" />
                    <RANKING order="5" place="5" resultid="2714" />
                    <RANKING order="6" place="6" resultid="4340" />
                    <RANKING order="7" place="7" resultid="2613" />
                    <RANKING order="8" place="8" resultid="2991" />
                    <RANKING order="9" place="9" resultid="4448" />
                    <RANKING order="10" place="10" resultid="2408" />
                    <RANKING order="11" place="11" resultid="4664" />
                    <RANKING order="12" place="12" resultid="2731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5877" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2473" />
                    <RANKING order="2" place="2" resultid="2469" />
                    <RANKING order="3" place="3" resultid="2969" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5878" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2695" />
                    <RANKING order="2" place="2" resultid="4434" />
                    <RANKING order="3" place="3" resultid="3953" />
                    <RANKING order="4" place="4" resultid="2569" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5879" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4285" />
                    <RANKING order="2" place="2" resultid="4281" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5095" daytime="11:54" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5096" daytime="11:56" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5097" daytime="11:58" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5098" daytime="12:00" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5099" daytime="12:02" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5100" daytime="12:04" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5101" daytime="12:06" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5102" daytime="12:08" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5103" daytime="12:10" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5104" daytime="12:12" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="5105" daytime="12:14" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="5106" daytime="12:16" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1104" daytime="12:18" gender="M" number="6" order="6" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5880" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2618" />
                    <RANKING order="2" place="2" resultid="2744" />
                    <RANKING order="3" place="3" resultid="3827" />
                    <RANKING order="4" place="4" resultid="4126" />
                    <RANKING order="5" place="5" resultid="3785" />
                    <RANKING order="6" place="6" resultid="2502" />
                    <RANKING order="7" place="7" resultid="4614" />
                    <RANKING order="8" place="8" resultid="3142" />
                    <RANKING order="9" place="9" resultid="2832" />
                    <RANKING order="10" place="9" resultid="3203" />
                    <RANKING order="11" place="11" resultid="4141" />
                    <RANKING order="12" place="12" resultid="4560" />
                    <RANKING order="13" place="13" resultid="2958" />
                    <RANKING order="14" place="14" resultid="4038" />
                    <RANKING order="15" place="15" resultid="3875" />
                    <RANKING order="16" place="16" resultid="2755" />
                    <RANKING order="17" place="17" resultid="2840" />
                    <RANKING order="18" place="18" resultid="4099" />
                    <RANKING order="19" place="19" resultid="3213" />
                    <RANKING order="20" place="20" resultid="2429" />
                    <RANKING order="21" place="21" resultid="2847" />
                    <RANKING order="22" place="22" resultid="2854" />
                    <RANKING order="23" place="23" resultid="2651" />
                    <RANKING order="24" place="24" resultid="2927" />
                    <RANKING order="25" place="25" resultid="4106" />
                    <RANKING order="26" place="26" resultid="4206" />
                    <RANKING order="27" place="27" resultid="3128" />
                    <RANKING order="28" place="28" resultid="2807" />
                    <RANKING order="29" place="-1" resultid="4620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5881" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2531" />
                    <RANKING order="2" place="2" resultid="3897" />
                    <RANKING order="3" place="3" resultid="3163" />
                    <RANKING order="4" place="4" resultid="3816" />
                    <RANKING order="5" place="5" resultid="3666" />
                    <RANKING order="6" place="6" resultid="3149" />
                    <RANKING order="7" place="7" resultid="3711" />
                    <RANKING order="8" place="8" resultid="3628" />
                    <RANKING order="9" place="9" resultid="3692" />
                    <RANKING order="10" place="10" resultid="4528" />
                    <RANKING order="11" place="11" resultid="4653" />
                    <RANKING order="12" place="12" resultid="3705" />
                    <RANKING order="13" place="13" resultid="2953" />
                    <RANKING order="14" place="14" resultid="2675" />
                    <RANKING order="15" place="15" resultid="3016" />
                    <RANKING order="16" place="16" resultid="3436" />
                    <RANKING order="17" place="17" resultid="2435" />
                    <RANKING order="18" place="18" resultid="4389" />
                    <RANKING order="19" place="19" resultid="2982" />
                    <RANKING order="20" place="20" resultid="3011" />
                    <RANKING order="21" place="21" resultid="4607" />
                    <RANKING order="22" place="22" resultid="3022" />
                    <RANKING order="23" place="-1" resultid="3672" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5882" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3498" />
                    <RANKING order="2" place="2" resultid="2525" />
                    <RANKING order="3" place="3" resultid="2443" />
                    <RANKING order="4" place="4" resultid="3977" />
                    <RANKING order="5" place="5" resultid="2936" />
                    <RANKING order="6" place="6" resultid="3946" />
                    <RANKING order="7" place="7" resultid="2483" />
                    <RANKING order="8" place="8" resultid="4461" />
                    <RANKING order="9" place="9" resultid="2607" />
                    <RANKING order="10" place="10" resultid="4454" />
                    <RANKING order="11" place="11" resultid="4490" />
                    <RANKING order="12" place="12" resultid="4033" />
                    <RANKING order="13" place="13" resultid="2976" />
                    <RANKING order="14" place="14" resultid="4119" />
                    <RANKING order="15" place="15" resultid="4632" />
                    <RANKING order="16" place="16" resultid="3005" />
                    <RANKING order="17" place="17" resultid="2921" />
                    <RANKING order="18" place="18" resultid="4333" />
                    <RANKING order="19" place="19" resultid="4042" />
                    <RANKING order="20" place="20" resultid="3585" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5883" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3935" />
                    <RANKING order="2" place="2" resultid="3881" />
                    <RANKING order="3" place="3" resultid="3575" />
                    <RANKING order="4" place="4" resultid="3052" />
                    <RANKING order="5" place="5" resultid="2538" />
                    <RANKING order="6" place="6" resultid="4476" />
                    <RANKING order="7" place="7" resultid="3581" />
                    <RANKING order="8" place="8" resultid="2801" />
                    <RANKING order="9" place="9" resultid="2870" />
                    <RANKING order="10" place="10" resultid="3569" />
                    <RANKING order="11" place="11" resultid="3910" />
                    <RANKING order="12" place="12" resultid="4441" />
                    <RANKING order="13" place="13" resultid="2995" />
                    <RANKING order="14" place="14" resultid="3564" />
                    <RANKING order="15" place="15" resultid="4148" />
                    <RANKING order="16" place="16" resultid="4397" />
                    <RANKING order="17" place="17" resultid="4081" />
                    <RANKING order="18" place="18" resultid="2768" />
                    <RANKING order="19" place="19" resultid="3108" />
                    <RANKING order="20" place="20" resultid="2986" />
                    <RANKING order="21" place="21" resultid="2664" />
                    <RANKING order="22" place="22" resultid="3179" />
                    <RANKING order="23" place="23" resultid="4276" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5884" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3553" />
                    <RANKING order="2" place="2" resultid="4427" />
                    <RANKING order="3" place="3" resultid="3559" />
                    <RANKING order="4" place="4" resultid="4249" />
                    <RANKING order="5" place="5" resultid="3965" />
                    <RANKING order="6" place="6" resultid="4366" />
                    <RANKING order="7" place="7" resultid="4183" />
                    <RANKING order="8" place="8" resultid="4187" />
                    <RANKING order="9" place="9" resultid="4291" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5885" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3982" />
                    <RANKING order="2" place="2" resultid="3479" />
                    <RANKING order="3" place="3" resultid="3960" />
                    <RANKING order="4" place="4" resultid="2887" />
                    <RANKING order="5" place="5" resultid="4323" />
                    <RANKING order="6" place="6" resultid="4553" />
                    <RANKING order="7" place="7" resultid="2578" />
                    <RANKING order="8" place="8" resultid="2898" />
                    <RANKING order="9" place="9" resultid="3192" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5886" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3808" />
                    <RANKING order="2" place="2" resultid="2563" />
                    <RANKING order="3" place="3" resultid="2790" />
                    <RANKING order="4" place="4" resultid="3891" />
                    <RANKING order="5" place="5" resultid="3048" />
                    <RANKING order="6" place="6" resultid="2780" />
                    <RANKING order="7" place="7" resultid="3059" />
                    <RANKING order="8" place="8" resultid="3073" />
                    <RANKING order="9" place="9" resultid="4329" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5114" daytime="12:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5115" daytime="12:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5116" daytime="12:22" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5117" daytime="12:24" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5118" daytime="12:26" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5119" daytime="12:28" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5120" daytime="12:28" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5121" daytime="12:30" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5122" daytime="12:32" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5123" daytime="12:34" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="5124" daytime="12:36" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="5125" daytime="12:38" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="5126" daytime="12:40" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="5127" daytime="12:42" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="5128" daytime="12:44" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="5129" daytime="12:46" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="5130" daytime="12:46" number="17" order="17" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-09-19" daytime="16:10" endtime="19:16" number="2" officialmeeting="15:30" teamleadermeeting="16:00" warmupfrom="15:00" warmupuntil="16:00">
          <EVENTS>
            <EVENT eventid="1112" daytime="16:40" gender="F" number="7" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6190" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3797" />
                    <RANKING order="2" place="2" resultid="3780" />
                    <RANKING order="3" place="3" resultid="3773" />
                    <RANKING order="4" place="4" resultid="3931" />
                    <RANKING order="5" place="5" resultid="3409" />
                    <RANKING order="6" place="6" resultid="4114" />
                    <RANKING order="7" place="7" resultid="3339" />
                    <RANKING order="8" place="8" resultid="2658" />
                    <RANKING order="9" place="9" resultid="3840" />
                    <RANKING order="10" place="10" resultid="3759" />
                    <RANKING order="11" place="11" resultid="2631" />
                    <RANKING order="12" place="12" resultid="4626" />
                    <RANKING order="13" place="13" resultid="2762" />
                    <RANKING order="14" place="14" resultid="3123" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6191" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3647" />
                    <RANKING order="2" place="2" resultid="2415" />
                    <RANKING order="3" place="3" resultid="3661" />
                    <RANKING order="4" place="4" resultid="3972" />
                    <RANKING order="5" place="5" resultid="3654" />
                    <RANKING order="6" place="6" resultid="2646" />
                    <RANKING order="7" place="7" resultid="3382" />
                    <RANKING order="8" place="8" resultid="4581" />
                    <RANKING order="9" place="9" resultid="3686" />
                    <RANKING order="10" place="10" resultid="4318" />
                    <RANKING order="11" place="11" resultid="3137" />
                    <RANKING order="12" place="12" resultid="4640" />
                    <RANKING order="13" place="13" resultid="4587" />
                    <RANKING order="14" place="14" resultid="3430" />
                    <RANKING order="15" place="15" resultid="2638" />
                    <RANKING order="16" place="16" resultid="4646" />
                    <RANKING order="17" place="17" resultid="2703" />
                    <RANKING order="18" place="-1" resultid="3234" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6192" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3525" />
                    <RANKING order="2" place="2" resultid="3475" />
                    <RANKING order="3" place="3" resultid="4155" />
                    <RANKING order="4" place="4" resultid="2465" />
                    <RANKING order="5" place="5" resultid="4469" />
                    <RANKING order="6" place="6" resultid="4483" />
                    <RANKING order="7" place="7" resultid="3101" />
                    <RANKING order="8" place="8" resultid="2948" />
                    <RANKING order="9" place="9" resultid="4508" />
                    <RANKING order="10" place="10" resultid="2819" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6193" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2709" />
                    <RANKING order="2" place="2" resultid="4341" />
                    <RANKING order="3" place="3" resultid="3039" />
                    <RANKING order="4" place="4" resultid="4373" />
                    <RANKING order="5" place="5" resultid="2866" />
                    <RANKING order="6" place="6" resultid="2796" />
                    <RANKING order="7" place="7" resultid="4665" />
                    <RANKING order="8" place="8" resultid="4449" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6194" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3547" />
                    <RANKING order="2" place="2" resultid="3515" />
                    <RANKING order="3" place="3" resultid="2970" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6195" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2774" />
                    <RANKING order="2" place="2" resultid="2460" />
                    <RANKING order="3" place="3" resultid="4056" />
                    <RANKING order="4" place="4" resultid="4240" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6196" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3904" />
                    <RANKING order="2" place="2" resultid="3916" />
                    <RANKING order="3" place="3" resultid="4282" />
                    <RANKING order="4" place="4" resultid="4286" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6197" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3904" />
                    <RANKING order="2" place="2" resultid="3525" />
                    <RANKING order="3" place="3" resultid="3916" />
                    <RANKING order="4" place="4" resultid="3475" />
                    <RANKING order="5" place="5" resultid="3547" />
                    <RANKING order="6" place="6" resultid="3515" />
                    <RANKING order="7" place="7" resultid="2774" />
                    <RANKING order="8" place="8" resultid="4155" />
                    <RANKING order="9" place="9" resultid="3647" />
                    <RANKING order="10" place="10" resultid="2465" />
                    <RANKING order="11" place="11" resultid="2415" />
                    <RANKING order="12" place="12" resultid="3797" />
                    <RANKING order="13" place="13" resultid="2709" />
                    <RANKING order="14" place="14" resultid="3661" />
                    <RANKING order="15" place="15" resultid="3972" />
                    <RANKING order="16" place="16" resultid="3780" />
                    <RANKING order="17" place="17" resultid="3654" />
                    <RANKING order="18" place="18" resultid="4341" />
                    <RANKING order="19" place="19" resultid="2646" />
                    <RANKING order="20" place="20" resultid="3039" />
                    <RANKING order="21" place="21" resultid="4373" />
                    <RANKING order="22" place="22" resultid="3382" />
                    <RANKING order="23" place="23" resultid="4581" />
                    <RANKING order="24" place="24" resultid="3773" />
                    <RANKING order="25" place="25" resultid="4469" />
                    <RANKING order="26" place="26" resultid="4483" />
                    <RANKING order="27" place="27" resultid="3686" />
                    <RANKING order="28" place="28" resultid="2866" />
                    <RANKING order="29" place="29" resultid="2796" />
                    <RANKING order="30" place="30" resultid="3931" />
                    <RANKING order="31" place="31" resultid="3409" />
                    <RANKING order="32" place="32" resultid="4114" />
                    <RANKING order="33" place="33" resultid="3339" />
                    <RANKING order="34" place="34" resultid="4318" />
                    <RANKING order="35" place="35" resultid="3137" />
                    <RANKING order="36" place="36" resultid="3101" />
                    <RANKING order="37" place="37" resultid="4640" />
                    <RANKING order="38" place="38" resultid="2460" />
                    <RANKING order="39" place="39" resultid="2948" />
                    <RANKING order="40" place="40" resultid="2658" />
                    <RANKING order="41" place="41" resultid="4587" />
                    <RANKING order="42" place="42" resultid="3430" />
                    <RANKING order="43" place="43" resultid="4508" />
                    <RANKING order="44" place="44" resultid="2819" />
                    <RANKING order="45" place="45" resultid="3840" />
                    <RANKING order="46" place="46" resultid="3759" />
                    <RANKING order="47" place="47" resultid="2638" />
                    <RANKING order="48" place="48" resultid="4646" />
                    <RANKING order="49" place="49" resultid="4282" />
                    <RANKING order="50" place="50" resultid="4286" />
                    <RANKING order="51" place="51" resultid="4665" />
                    <RANKING order="52" place="52" resultid="4449" />
                    <RANKING order="53" place="53" resultid="4056" />
                    <RANKING order="54" place="54" resultid="2631" />
                    <RANKING order="55" place="55" resultid="2703" />
                    <RANKING order="56" place="56" resultid="4626" />
                    <RANKING order="57" place="57" resultid="4240" />
                    <RANKING order="58" place="58" resultid="2762" />
                    <RANKING order="59" place="59" resultid="2970" />
                    <RANKING order="60" place="60" resultid="3123" />
                    <RANKING order="61" place="-1" resultid="3234" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5138" daytime="16:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5139" daytime="16:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5140" daytime="16:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5141" daytime="16:52" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5142" daytime="16:56" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5143" daytime="17:00" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5144" daytime="17:04" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5145" daytime="17:08" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5146" daytime="17:12" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1120" daytime="17:18" gender="M" number="8" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6198" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3311" />
                    <RANKING order="2" place="2" resultid="3828" />
                    <RANKING order="3" place="3" resultid="3735" />
                    <RANKING order="4" place="4" resultid="2619" />
                    <RANKING order="5" place="5" resultid="3144" />
                    <RANKING order="6" place="6" resultid="3730" />
                    <RANKING order="7" place="7" resultid="3204" />
                    <RANKING order="8" place="8" resultid="4541" />
                    <RANKING order="9" place="9" resultid="3742" />
                    <RANKING order="10" place="10" resultid="3722" />
                    <RANKING order="11" place="11" resultid="4128" />
                    <RANKING order="12" place="12" resultid="4615" />
                    <RANKING order="13" place="13" resultid="4344" />
                    <RANKING order="14" place="14" resultid="4039" />
                    <RANKING order="15" place="15" resultid="4142" />
                    <RANKING order="16" place="16" resultid="2625" />
                    <RANKING order="17" place="17" resultid="2833" />
                    <RANKING order="18" place="18" resultid="2557" />
                    <RANKING order="19" place="19" resultid="3876" />
                    <RANKING order="20" place="20" resultid="2430" />
                    <RANKING order="21" place="21" resultid="3222" />
                    <RANKING order="22" place="22" resultid="3214" />
                    <RANKING order="23" place="23" resultid="3129" />
                    <RANKING order="24" place="24" resultid="2808" />
                    <RANKING order="25" place="25" resultid="4107" />
                    <RANKING order="26" place="-1" resultid="4621" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6199" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2533" />
                    <RANKING order="2" place="2" resultid="3667" />
                    <RANKING order="3" place="3" resultid="3817" />
                    <RANKING order="4" place="4" resultid="3290" />
                    <RANKING order="5" place="5" resultid="3898" />
                    <RANKING order="6" place="6" resultid="3673" />
                    <RANKING order="7" place="7" resultid="3713" />
                    <RANKING order="8" place="8" resultid="4655" />
                    <RANKING order="9" place="9" resultid="3298" />
                    <RANKING order="10" place="10" resultid="3164" />
                    <RANKING order="11" place="11" resultid="3635" />
                    <RANKING order="12" place="12" resultid="3706" />
                    <RANKING order="13" place="13" resultid="4595" />
                    <RANKING order="14" place="14" resultid="2676" />
                    <RANKING order="15" place="15" resultid="4270" />
                    <RANKING order="16" place="16" resultid="2954" />
                    <RANKING order="17" place="17" resultid="2436" />
                    <RANKING order="18" place="18" resultid="4660" />
                    <RANKING order="19" place="19" resultid="3017" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6200" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3541" />
                    <RANKING order="2" place="2" resultid="2444" />
                    <RANKING order="3" place="3" resultid="3499" />
                    <RANKING order="4" place="4" resultid="3618" />
                    <RANKING order="5" place="5" resultid="4462" />
                    <RANKING order="6" place="6" resultid="3590" />
                    <RANKING order="7" place="7" resultid="4491" />
                    <RANKING order="8" place="8" resultid="2489" />
                    <RANKING order="9" place="9" resultid="4120" />
                    <RANKING order="10" place="10" resultid="4634" />
                    <RANKING order="11" place="11" resultid="4034" />
                    <RANKING order="12" place="12" resultid="4334" />
                    <RANKING order="13" place="13" resultid="2977" />
                    <RANKING order="14" place="14" resultid="3006" />
                    <RANKING order="15" place="15" resultid="4043" />
                    <RANKING order="16" place="16" resultid="3210" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6201" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3487" />
                    <RANKING order="2" place="2" resultid="3257" />
                    <RANKING order="3" place="3" resultid="3822" />
                    <RANKING order="4" place="4" resultid="3882" />
                    <RANKING order="5" place="5" resultid="3624" />
                    <RANKING order="6" place="6" resultid="3360" />
                    <RANKING order="7" place="7" resultid="3582" />
                    <RANKING order="8" place="8" resultid="4477" />
                    <RANKING order="9" place="9" resultid="4059" />
                    <RANKING order="10" place="10" resultid="2996" />
                    <RANKING order="11" place="11" resultid="3053" />
                    <RANKING order="12" place="12" resultid="2802" />
                    <RANKING order="13" place="13" resultid="3115" />
                    <RANKING order="14" place="14" resultid="2551" />
                    <RANKING order="15" place="15" resultid="3180" />
                    <RANKING order="16" place="16" resultid="3219" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6202" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3554" />
                    <RANKING order="2" place="2" resultid="3520" />
                    <RANKING order="3" place="3" resultid="4428" />
                    <RANKING order="4" place="4" resultid="3966" />
                    <RANKING order="5" place="5" resultid="4367" />
                    <RANKING order="6" place="6" resultid="4293" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6203" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3961" />
                    <RANKING order="2" place="2" resultid="4499" />
                    <RANKING order="3" place="3" resultid="3081" />
                    <RANKING order="4" place="4" resultid="2899" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6204" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3892" />
                    <RANKING order="2" place="2" resultid="4330" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6205" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3554" />
                    <RANKING order="2" place="2" resultid="3961" />
                    <RANKING order="3" place="3" resultid="4499" />
                    <RANKING order="4" place="4" resultid="3520" />
                    <RANKING order="5" place="5" resultid="3487" />
                    <RANKING order="6" place="6" resultid="4428" />
                    <RANKING order="7" place="7" resultid="3257" />
                    <RANKING order="8" place="8" resultid="3822" />
                    <RANKING order="9" place="9" resultid="3541" />
                    <RANKING order="10" place="10" resultid="2444" />
                    <RANKING order="11" place="11" resultid="3499" />
                    <RANKING order="12" place="12" resultid="2533" />
                    <RANKING order="13" place="13" resultid="3667" />
                    <RANKING order="14" place="14" resultid="3966" />
                    <RANKING order="15" place="15" resultid="3817" />
                    <RANKING order="16" place="16" resultid="3290" />
                    <RANKING order="17" place="17" resultid="3898" />
                    <RANKING order="18" place="18" resultid="3892" />
                    <RANKING order="19" place="19" resultid="3882" />
                    <RANKING order="20" place="20" resultid="4367" />
                    <RANKING order="21" place="21" resultid="3624" />
                    <RANKING order="22" place="22" resultid="3081" />
                    <RANKING order="23" place="23" resultid="3360" />
                    <RANKING order="24" place="24" resultid="3618" />
                    <RANKING order="25" place="25" resultid="3311" />
                    <RANKING order="26" place="26" resultid="3673" />
                    <RANKING order="27" place="27" resultid="4462" />
                    <RANKING order="28" place="28" resultid="3582" />
                    <RANKING order="29" place="29" resultid="2899" />
                    <RANKING order="30" place="30" resultid="3590" />
                    <RANKING order="31" place="31" resultid="3713" />
                    <RANKING order="32" place="32" resultid="4477" />
                    <RANKING order="33" place="33" resultid="3828" />
                    <RANKING order="34" place="34" resultid="4491" />
                    <RANKING order="35" place="35" resultid="3735" />
                    <RANKING order="36" place="36" resultid="4059" />
                    <RANKING order="37" place="37" resultid="4330" />
                    <RANKING order="38" place="38" resultid="2996" />
                    <RANKING order="39" place="39" resultid="2619" />
                    <RANKING order="40" place="40" resultid="3053" />
                    <RANKING order="41" place="41" resultid="4655" />
                    <RANKING order="42" place="42" resultid="2489" />
                    <RANKING order="43" place="43" resultid="3298" />
                    <RANKING order="44" place="44" resultid="4120" />
                    <RANKING order="45" place="45" resultid="3144" />
                    <RANKING order="46" place="46" resultid="4634" />
                    <RANKING order="47" place="47" resultid="2802" />
                    <RANKING order="48" place="47" resultid="3164" />
                    <RANKING order="49" place="49" resultid="4034" />
                    <RANKING order="50" place="50" resultid="3115" />
                    <RANKING order="51" place="51" resultid="3730" />
                    <RANKING order="52" place="52" resultid="3635" />
                    <RANKING order="53" place="53" resultid="4334" />
                    <RANKING order="54" place="54" resultid="3204" />
                    <RANKING order="55" place="55" resultid="2551" />
                    <RANKING order="56" place="56" resultid="4541" />
                    <RANKING order="57" place="57" resultid="2977" />
                    <RANKING order="58" place="58" resultid="3706" />
                    <RANKING order="59" place="59" resultid="4595" />
                    <RANKING order="60" place="60" resultid="3742" />
                    <RANKING order="61" place="61" resultid="3722" />
                    <RANKING order="62" place="62" resultid="4128" />
                    <RANKING order="63" place="63" resultid="4293" />
                    <RANKING order="64" place="64" resultid="4615" />
                    <RANKING order="65" place="65" resultid="4344" />
                    <RANKING order="66" place="66" resultid="3180" />
                    <RANKING order="67" place="67" resultid="4039" />
                    <RANKING order="68" place="68" resultid="4142" />
                    <RANKING order="69" place="69" resultid="2625" />
                    <RANKING order="70" place="70" resultid="2676" />
                    <RANKING order="71" place="71" resultid="4270" />
                    <RANKING order="72" place="72" resultid="2833" />
                    <RANKING order="73" place="73" resultid="2557" />
                    <RANKING order="74" place="74" resultid="2954" />
                    <RANKING order="75" place="75" resultid="3006" />
                    <RANKING order="76" place="76" resultid="4043" />
                    <RANKING order="77" place="77" resultid="2436" />
                    <RANKING order="78" place="78" resultid="4660" />
                    <RANKING order="79" place="79" resultid="3219" />
                    <RANKING order="80" place="80" resultid="3876" />
                    <RANKING order="81" place="81" resultid="3017" />
                    <RANKING order="82" place="82" resultid="2430" />
                    <RANKING order="83" place="83" resultid="3222" />
                    <RANKING order="84" place="84" resultid="3214" />
                    <RANKING order="85" place="85" resultid="3210" />
                    <RANKING order="86" place="86" resultid="3129" />
                    <RANKING order="87" place="87" resultid="2808" />
                    <RANKING order="88" place="88" resultid="4107" />
                    <RANKING order="89" place="-1" resultid="4621" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5147" daytime="17:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5148" daytime="17:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5149" daytime="17:26" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5150" daytime="17:30" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5151" daytime="17:34" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5152" daytime="17:38" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5153" daytime="17:42" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5154" daytime="17:46" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5155" daytime="17:50" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5156" daytime="17:52" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="5157" daytime="17:56" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="5158" daytime="18:00" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1128" daytime="18:04" gender="F" number="9" order="4" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5887" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3851" />
                    <RANKING order="2" place="2" resultid="4170" />
                    <RANKING order="3" place="3" resultid="3332" />
                    <RANKING order="4" place="4" resultid="3423" />
                    <RANKING order="5" place="5" resultid="3374" />
                    <RANKING order="6" place="6" resultid="2739" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5888" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3698" />
                    <RANKING order="2" place="2" resultid="4547" />
                    <RANKING order="3" place="3" resultid="2645" />
                    <RANKING order="4" place="4" resultid="3136" />
                    <RANKING order="5" place="5" resultid="2422" />
                    <RANKING order="6" place="6" resultid="2826" />
                    <RANKING order="7" place="7" resultid="3835" />
                    <RANKING order="8" place="8" resultid="4639" />
                    <RANKING order="9" place="9" resultid="4359" />
                    <RANKING order="10" place="10" resultid="4352" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5889" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4421" />
                    <RANKING order="2" place="2" resultid="3609" />
                    <RANKING order="3" place="3" resultid="2597" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5890" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3038" />
                    <RANKING order="2" place="2" resultid="2708" />
                    <RANKING order="3" place="3" resultid="2732" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5891" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3249" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5892" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4435" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5893" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5159" daytime="18:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5160" daytime="18:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5161" daytime="18:10" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5162" daytime="18:12" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1135" daytime="18:16" gender="M" number="10" order="5" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5894" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3765" />
                    <RANKING order="2" place="2" resultid="4561" />
                    <RANKING order="3" place="3" resultid="3143" />
                    <RANKING order="4" place="4" resultid="3729" />
                    <RANKING order="5" place="5" resultid="3346" />
                    <RANKING order="6" place="6" resultid="4127" />
                    <RANKING order="7" place="7" resultid="4134" />
                    <RANKING order="8" place="8" resultid="3791" />
                    <RANKING order="9" place="9" resultid="4100" />
                    <RANKING order="10" place="10" resultid="2841" />
                    <RANKING order="11" place="11" resultid="4207" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5895" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2532" />
                    <RANKING order="2" place="2" resultid="3150" />
                    <RANKING order="3" place="3" resultid="4529" />
                    <RANKING order="4" place="4" resultid="3629" />
                    <RANKING order="5" place="5" resultid="3297" />
                    <RANKING order="6" place="6" resultid="3437" />
                    <RANKING order="7" place="7" resultid="4390" />
                    <RANKING order="8" place="8" resultid="3712" />
                    <RANKING order="9" place="9" resultid="4594" />
                    <RANKING order="10" place="10" resultid="4654" />
                    <RANKING order="11" place="11" resultid="4085" />
                    <RANKING order="12" place="12" resultid="4162" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5896" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2526" />
                    <RANKING order="2" place="2" resultid="3947" />
                    <RANKING order="3" place="3" resultid="3352" />
                    <RANKING order="4" place="4" resultid="2450" />
                    <RANKING order="5" place="5" resultid="3269" />
                    <RANKING order="6" place="6" resultid="4455" />
                    <RANKING order="7" place="7" resultid="2608" />
                    <RANKING order="8" place="8" resultid="2484" />
                    <RANKING order="9" place="9" resultid="2916" />
                    <RANKING order="10" place="10" resultid="2922" />
                    <RANKING order="11" place="11" resultid="2546" />
                    <RANKING order="12" place="12" resultid="4633" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5897" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3503" />
                    <RANKING order="2" place="2" resultid="3576" />
                    <RANKING order="3" place="3" resultid="3395" />
                    <RANKING order="4" place="4" resultid="4149" />
                    <RANKING order="5" place="5" resultid="3911" />
                    <RANKING order="6" place="6" resultid="4442" />
                    <RANKING order="7" place="7" resultid="3565" />
                    <RANKING order="8" place="8" resultid="2539" />
                    <RANKING order="9" place="9" resultid="2665" />
                    <RANKING order="10" place="10" resultid="4398" />
                    <RANKING order="11" place="11" resultid="3109" />
                    <RANKING order="12" place="-1" resultid="2987" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5898" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2401" />
                    <RANKING order="2" place="2" resultid="3519" />
                    <RANKING order="3" place="3" resultid="4250" />
                    <RANKING order="4" place="4" resultid="3095" />
                    <RANKING order="5" place="5" resultid="4292" />
                    <RANKING order="6" place="6" resultid="4188" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5899" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3480" />
                    <RANKING order="2" place="2" resultid="3983" />
                    <RANKING order="3" place="3" resultid="3716" />
                    <RANKING order="4" place="4" resultid="3067" />
                    <RANKING order="5" place="5" resultid="4554" />
                    <RANKING order="6" place="6" resultid="3244" />
                    <RANKING order="7" place="7" resultid="4324" />
                    <RANKING order="8" place="8" resultid="2579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="5900" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3809" />
                    <RANKING order="2" place="2" resultid="2564" />
                    <RANKING order="3" place="3" resultid="2785" />
                    <RANKING order="4" place="4" resultid="3060" />
                    <RANKING order="5" place="5" resultid="2781" />
                    <RANKING order="6" place="6" resultid="2910" />
                    <RANKING order="7" place="7" resultid="2893" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5169" daytime="18:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5170" daytime="18:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5171" daytime="18:20" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5172" daytime="18:24" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5173" daytime="18:26" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5174" daytime="18:28" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5175" daytime="18:32" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5176" daytime="18:34" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5177" daytime="18:36" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5178" daytime="18:38" number="10" order="10" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1143" daytime="18:42" gender="F" number="11" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6206" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3852" />
                    <RANKING order="2" place="2" resultid="3333" />
                    <RANKING order="3" place="3" resultid="3746" />
                    <RANKING order="4" place="4" resultid="3841" />
                    <RANKING order="5" place="5" resultid="4171" />
                    <RANKING order="6" place="6" resultid="3923" />
                    <RANKING order="7" place="7" resultid="3375" />
                    <RANKING order="8" place="8" resultid="4567" />
                    <RANKING order="9" place="9" resultid="2670" />
                    <RANKING order="10" place="10" resultid="4071" />
                    <RANKING order="11" place="11" resultid="4177" />
                    <RANKING order="12" place="12" resultid="2721" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6207" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3276" />
                    <RANKING order="2" place="2" resultid="3699" />
                    <RANKING order="3" place="3" resultid="3383" />
                    <RANKING order="4" place="4" resultid="3530" />
                    <RANKING order="5" place="5" resultid="4263" />
                    <RANKING order="6" place="6" resultid="3648" />
                    <RANKING order="7" place="7" resultid="4588" />
                    <RANKING order="8" place="8" resultid="3973" />
                    <RANKING order="9" place="9" resultid="3836" />
                    <RANKING order="10" place="10" resultid="3157" />
                    <RANKING order="11" place="-1" resultid="4647" />
                    <RANKING order="12" place="-1" resultid="3886" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6208" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3463" />
                    <RANKING order="2" place="2" resultid="2876" />
                    <RANKING order="3" place="3" resultid="3283" />
                    <RANKING order="4" place="4" resultid="3536" />
                    <RANKING order="5" place="5" resultid="3599" />
                    <RANKING order="6" place="6" resultid="4156" />
                    <RANKING order="7" place="7" resultid="3594" />
                    <RANKING order="8" place="8" resultid="2943" />
                    <RANKING order="9" place="9" resultid="3188" />
                    <RANKING order="10" place="10" resultid="4068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6209" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3469" />
                    <RANKING order="2" place="2" resultid="3318" />
                    <RANKING order="3" place="3" resultid="3941" />
                    <RANKING order="4" place="4" resultid="2409" />
                    <RANKING order="5" place="5" resultid="2715" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6210" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4193" />
                    <RANKING order="2" place="2" resultid="2964" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6211" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2696" />
                    <RANKING order="2" place="2" resultid="3954" />
                    <RANKING order="3" place="3" resultid="4306" />
                    <RANKING order="4" place="4" resultid="4057" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6212" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3905" />
                    <RANKING order="2" place="2" resultid="4283" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6213" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3905" />
                    <RANKING order="2" place="2" resultid="3469" />
                    <RANKING order="3" place="3" resultid="3318" />
                    <RANKING order="4" place="4" resultid="3852" />
                    <RANKING order="5" place="5" resultid="3463" />
                    <RANKING order="6" place="6" resultid="2876" />
                    <RANKING order="7" place="7" resultid="2696" />
                    <RANKING order="8" place="8" resultid="3276" />
                    <RANKING order="9" place="9" resultid="3699" />
                    <RANKING order="10" place="10" resultid="3283" />
                    <RANKING order="11" place="11" resultid="3536" />
                    <RANKING order="12" place="12" resultid="3599" />
                    <RANKING order="13" place="13" resultid="3333" />
                    <RANKING order="14" place="14" resultid="3954" />
                    <RANKING order="15" place="15" resultid="3383" />
                    <RANKING order="16" place="16" resultid="3746" />
                    <RANKING order="17" place="17" resultid="3941" />
                    <RANKING order="18" place="18" resultid="4156" />
                    <RANKING order="19" place="19" resultid="3594" />
                    <RANKING order="20" place="20" resultid="3530" />
                    <RANKING order="21" place="21" resultid="4263" />
                    <RANKING order="22" place="22" resultid="3648" />
                    <RANKING order="23" place="23" resultid="3841" />
                    <RANKING order="24" place="24" resultid="4588" />
                    <RANKING order="25" place="25" resultid="4193" />
                    <RANKING order="26" place="26" resultid="3973" />
                    <RANKING order="27" place="27" resultid="2943" />
                    <RANKING order="28" place="28" resultid="2409" />
                    <RANKING order="29" place="29" resultid="2715" />
                    <RANKING order="30" place="30" resultid="4171" />
                    <RANKING order="31" place="31" resultid="4306" />
                    <RANKING order="32" place="32" resultid="3923" />
                    <RANKING order="33" place="33" resultid="3836" />
                    <RANKING order="34" place="34" resultid="3157" />
                    <RANKING order="35" place="35" resultid="3375" />
                    <RANKING order="36" place="36" resultid="4567" />
                    <RANKING order="37" place="37" resultid="3188" />
                    <RANKING order="38" place="38" resultid="4283" />
                    <RANKING order="39" place="39" resultid="2670" />
                    <RANKING order="40" place="40" resultid="4071" />
                    <RANKING order="41" place="41" resultid="4057" />
                    <RANKING order="42" place="42" resultid="4177" />
                    <RANKING order="43" place="43" resultid="2964" />
                    <RANKING order="44" place="44" resultid="2721" />
                    <RANKING order="45" place="45" resultid="4068" />
                    <RANKING order="46" place="-1" resultid="4647" />
                    <RANKING order="47" place="-1" resultid="3886" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5186" daytime="18:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5187" daytime="18:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5188" daytime="18:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5189" daytime="18:54" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5190" daytime="19:00" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5191" daytime="19:04" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1151" daytime="19:08" gender="M" number="12" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6214" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3325" />
                    <RANKING order="2" place="2" resultid="3736" />
                    <RANKING order="3" place="3" resultid="3402" />
                    <RANKING order="4" place="4" resultid="3803" />
                    <RANKING order="5" place="5" resultid="3416" />
                    <RANKING order="6" place="6" resultid="3347" />
                    <RANKING order="7" place="7" resultid="4520" />
                    <RANKING order="8" place="8" resultid="3766" />
                    <RANKING order="9" place="9" resultid="3792" />
                    <RANKING order="10" place="10" resultid="3863" />
                    <RANKING order="11" place="11" resultid="4536" />
                    <RANKING order="12" place="12" resultid="3367" />
                    <RANKING order="13" place="13" resultid="4199" />
                    <RANKING order="14" place="14" resultid="2959" />
                    <RANKING order="15" place="15" resultid="3215" />
                    <RANKING order="16" place="16" resultid="3752" />
                    <RANKING order="17" place="17" resultid="2652" />
                    <RANKING order="18" place="18" resultid="2848" />
                    <RANKING order="19" place="-1" resultid="4562" />
                    <RANKING order="20" place="-1" resultid="4574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6215" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3291" />
                    <RANKING order="2" place="2" resultid="2931" />
                    <RANKING order="3" place="3" resultid="3388" />
                    <RANKING order="4" place="4" resultid="3693" />
                    <RANKING order="5" place="5" resultid="3630" />
                    <RANKING order="6" place="6" resultid="3707" />
                    <RANKING order="7" place="7" resultid="4391" />
                    <RANKING order="8" place="8" resultid="4075" />
                    <RANKING order="9" place="9" resultid="4608" />
                    <RANKING order="10" place="10" resultid="4086" />
                    <RANKING order="11" place="-1" resultid="3679" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6216" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2881" />
                    <RANKING order="2" place="2" resultid="2451" />
                    <RANKING order="3" place="3" resultid="4601" />
                    <RANKING order="4" place="4" resultid="4456" />
                    <RANKING order="5" place="5" resultid="3353" />
                    <RANKING order="6" place="6" resultid="4299" />
                    <RANKING order="7" place="7" resultid="4256" />
                    <RANKING order="8" place="8" resultid="3604" />
                    <RANKING order="9" place="9" resultid="4121" />
                    <RANKING order="10" place="10" resultid="4335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6217" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3493" />
                    <RANKING order="2" place="2" resultid="3258" />
                    <RANKING order="3" place="3" resultid="3508" />
                    <RANKING order="4" place="4" resultid="3858" />
                    <RANKING order="5" place="5" resultid="3570" />
                    <RANKING order="6" place="6" resultid="2602" />
                    <RANKING order="7" place="7" resultid="3088" />
                    <RANKING order="8" place="8" resultid="3869" />
                    <RANKING order="9" place="9" resultid="3116" />
                    <RANKING order="10" place="10" resultid="3054" />
                    <RANKING order="11" place="-1" resultid="4053" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6218" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3560" />
                    <RANKING order="2" place="2" resultid="4429" />
                    <RANKING order="3" place="3" resultid="3304" />
                    <RANKING order="4" place="4" resultid="4063" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6219" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4500" />
                    <RANKING order="2" place="2" resultid="4235" />
                    <RANKING order="3" place="3" resultid="3193" />
                    <RANKING order="4" place="-1" resultid="2574" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6220" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4331" />
                    <RANKING order="2" place="2" resultid="3074" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6221" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3493" />
                    <RANKING order="2" place="2" resultid="2881" />
                    <RANKING order="3" place="3" resultid="3560" />
                    <RANKING order="4" place="4" resultid="2451" />
                    <RANKING order="5" place="5" resultid="4429" />
                    <RANKING order="6" place="6" resultid="3291" />
                    <RANKING order="7" place="7" resultid="2931" />
                    <RANKING order="8" place="8" resultid="3258" />
                    <RANKING order="9" place="9" resultid="4500" />
                    <RANKING order="10" place="10" resultid="4601" />
                    <RANKING order="11" place="11" resultid="3508" />
                    <RANKING order="12" place="12" resultid="4456" />
                    <RANKING order="13" place="13" resultid="3353" />
                    <RANKING order="14" place="14" resultid="3858" />
                    <RANKING order="15" place="15" resultid="3304" />
                    <RANKING order="16" place="16" resultid="3570" />
                    <RANKING order="17" place="17" resultid="2602" />
                    <RANKING order="18" place="18" resultid="4299" />
                    <RANKING order="19" place="19" resultid="4256" />
                    <RANKING order="20" place="20" resultid="3088" />
                    <RANKING order="21" place="21" resultid="3388" />
                    <RANKING order="22" place="22" resultid="3604" />
                    <RANKING order="23" place="23" resultid="3325" />
                    <RANKING order="24" place="24" resultid="3869" />
                    <RANKING order="25" place="25" resultid="3736" />
                    <RANKING order="26" place="26" resultid="3693" />
                    <RANKING order="27" place="27" resultid="4121" />
                    <RANKING order="28" place="28" resultid="4331" />
                    <RANKING order="29" place="29" resultid="3116" />
                    <RANKING order="30" place="30" resultid="3630" />
                    <RANKING order="31" place="31" resultid="3402" />
                    <RANKING order="32" place="32" resultid="3074" />
                    <RANKING order="33" place="33" resultid="3054" />
                    <RANKING order="34" place="34" resultid="3803" />
                    <RANKING order="35" place="35" resultid="3416" />
                    <RANKING order="36" place="36" resultid="3707" />
                    <RANKING order="37" place="37" resultid="3347" />
                    <RANKING order="38" place="38" resultid="4235" />
                    <RANKING order="39" place="39" resultid="4520" />
                    <RANKING order="40" place="40" resultid="4335" />
                    <RANKING order="41" place="41" resultid="3766" />
                    <RANKING order="42" place="42" resultid="3792" />
                    <RANKING order="43" place="43" resultid="3863" />
                    <RANKING order="44" place="44" resultid="3193" />
                    <RANKING order="45" place="45" resultid="4391" />
                    <RANKING order="46" place="46" resultid="4536" />
                    <RANKING order="47" place="47" resultid="3367" />
                    <RANKING order="48" place="48" resultid="4075" />
                    <RANKING order="49" place="49" resultid="4063" />
                    <RANKING order="50" place="50" resultid="4608" />
                    <RANKING order="51" place="51" resultid="4199" />
                    <RANKING order="52" place="52" resultid="2959" />
                    <RANKING order="53" place="53" resultid="4086" />
                    <RANKING order="54" place="54" resultid="3215" />
                    <RANKING order="55" place="55" resultid="3752" />
                    <RANKING order="56" place="56" resultid="2652" />
                    <RANKING order="57" place="57" resultid="2848" />
                    <RANKING order="58" place="-1" resultid="3679" />
                    <RANKING order="59" place="-1" resultid="4562" />
                    <RANKING order="60" place="-1" resultid="4574" />
                    <RANKING order="61" place="-1" resultid="2574" />
                    <RANKING order="62" place="-1" resultid="4053" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5192" daytime="19:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5193" daytime="19:14" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5194" daytime="19:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5195" daytime="19:22" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5196" daytime="19:26" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5197" daytime="19:30" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5198" daytime="19:36" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5199" daytime="19:38" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5200" daytime="19:44" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-09-20" daytime="09:10" endtime="11:51" number="3" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1159" daytime="09:10" gender="F" number="13" order="1" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6024" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3781" />
                    <RANKING order="2" place="2" resultid="4173" />
                    <RANKING order="3" place="3" resultid="3410" />
                    <RANKING order="4" place="4" resultid="3747" />
                    <RANKING order="5" place="5" resultid="4115" />
                    <RANKING order="6" place="6" resultid="4048" />
                    <RANKING order="7" place="7" resultid="3843" />
                    <RANKING order="8" place="8" resultid="3925" />
                    <RANKING order="9" place="9" resultid="2633" />
                    <RANKING order="10" place="10" resultid="4245" />
                    <RANKING order="11" place="11" resultid="4515" />
                    <RANKING order="12" place="12" resultid="4628" />
                    <RANKING order="13" place="13" resultid="2764" />
                    <RANKING order="14" place="14" resultid="3124" />
                    <RANKING order="15" place="15" resultid="2722" />
                    <RANKING order="16" place="-1" resultid="3198" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6025" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3649" />
                    <RANKING order="2" place="2" resultid="3974" />
                    <RANKING order="3" place="3" resultid="2417" />
                    <RANKING order="4" place="4" resultid="2647" />
                    <RANKING order="5" place="5" resultid="2727" />
                    <RANKING order="6" place="6" resultid="2424" />
                    <RANKING order="7" place="7" resultid="3656" />
                    <RANKING order="8" place="8" resultid="3531" />
                    <RANKING order="9" place="9" resultid="3663" />
                    <RANKING order="10" place="10" resultid="4582" />
                    <RANKING order="11" place="11" resultid="4548" />
                    <RANKING order="12" place="12" resultid="3432" />
                    <RANKING order="13" place="13" resultid="4641" />
                    <RANKING order="14" place="14" resultid="4589" />
                    <RANKING order="15" place="15" resultid="3642" />
                    <RANKING order="16" place="16" resultid="3235" />
                    <RANKING order="17" place="17" resultid="4214" />
                    <RANKING order="18" place="18" resultid="2518" />
                    <RANKING order="19" place="19" resultid="2704" />
                    <RANKING order="20" place="20" resultid="2498" />
                    <RANKING order="21" place="21" resultid="4360" />
                    <RANKING order="22" place="22" resultid="2507" />
                    <RANKING order="23" place="23" resultid="2752" />
                    <RANKING order="24" place="-1" resultid="3887" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6026" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4422" />
                    <RANKING order="2" place="2" resultid="3476" />
                    <RANKING order="3" place="3" resultid="4157" />
                    <RANKING order="4" place="4" resultid="4470" />
                    <RANKING order="5" place="5" resultid="2821" />
                    <RANKING order="6" place="6" resultid="2949" />
                    <RANKING order="7" place="7" resultid="4485" />
                    <RANKING order="8" place="8" resultid="4509" />
                    <RANKING order="9" place="9" resultid="3103" />
                    <RANKING order="10" place="10" resultid="4381" />
                    <RANKING order="11" place="11" resultid="3231" />
                    <RANKING order="12" place="-1" resultid="2598" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6027" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3471" />
                    <RANKING order="2" place="2" resultid="4374" />
                    <RANKING order="3" place="3" resultid="2711" />
                    <RANKING order="4" place="4" resultid="3319" />
                    <RANKING order="5" place="5" resultid="2992" />
                    <RANKING order="6" place="6" resultid="4450" />
                    <RANKING order="7" place="7" resultid="4666" />
                    <RANKING order="8" place="8" resultid="2734" />
                    <RANKING order="9" place="-1" resultid="3459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6028" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3548" />
                    <RANKING order="2" place="2" resultid="2470" />
                    <RANKING order="3" place="3" resultid="2965" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6029" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2698" />
                    <RANKING order="2" place="2" resultid="2776" />
                    <RANKING order="3" place="3" resultid="4436" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6030" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4287" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5201" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5202" daytime="09:12" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5203" daytime="09:16" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5204" daytime="09:18" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5205" daytime="09:20" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5206" daytime="09:22" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5207" daytime="09:26" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5208" daytime="09:28" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5209" daytime="09:30" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1167" daytime="09:34" gender="M" number="14" order="2" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6031" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2620" />
                    <RANKING order="2" place="2" resultid="3830" />
                    <RANKING order="3" place="3" resultid="3786" />
                    <RANKING order="4" place="4" resultid="2746" />
                    <RANKING order="5" place="5" resultid="3205" />
                    <RANKING order="6" place="6" resultid="3145" />
                    <RANKING order="7" place="7" resultid="4616" />
                    <RANKING order="8" place="8" resultid="2503" />
                    <RANKING order="9" place="9" resultid="3326" />
                    <RANKING order="10" place="10" resultid="4144" />
                    <RANKING order="11" place="11" resultid="4542" />
                    <RANKING order="12" place="12" resultid="4563" />
                    <RANKING order="13" place="13" resultid="2834" />
                    <RANKING order="14" place="14" resultid="3877" />
                    <RANKING order="15" place="15" resultid="4040" />
                    <RANKING order="16" place="16" resultid="2558" />
                    <RANKING order="17" place="17" resultid="2960" />
                    <RANKING order="18" place="18" resultid="4575" />
                    <RANKING order="19" place="19" resultid="2756" />
                    <RANKING order="20" place="20" resultid="2431" />
                    <RANKING order="21" place="21" resultid="2849" />
                    <RANKING order="22" place="21" resultid="2855" />
                    <RANKING order="23" place="23" resultid="2842" />
                    <RANKING order="24" place="24" resultid="2653" />
                    <RANKING order="25" place="25" resultid="3368" />
                    <RANKING order="26" place="26" resultid="3216" />
                    <RANKING order="27" place="27" resultid="4108" />
                    <RANKING order="28" place="28" resultid="2928" />
                    <RANKING order="29" place="29" resultid="2809" />
                    <RANKING order="30" place="30" resultid="4208" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6032" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2534" />
                    <RANKING order="2" place="2" resultid="3668" />
                    <RANKING order="3" place="3" resultid="3900" />
                    <RANKING order="4" place="4" resultid="3818" />
                    <RANKING order="5" place="5" resultid="3166" />
                    <RANKING order="6" place="6" resultid="3675" />
                    <RANKING order="7" place="7" resultid="3694" />
                    <RANKING order="8" place="8" resultid="4530" />
                    <RANKING order="9" place="9" resultid="4656" />
                    <RANKING order="10" place="10" resultid="3631" />
                    <RANKING order="11" place="11" resultid="3708" />
                    <RANKING order="12" place="12" resultid="3299" />
                    <RANKING order="13" place="13" resultid="2677" />
                    <RANKING order="14" place="14" resultid="4163" />
                    <RANKING order="15" place="15" resultid="3438" />
                    <RANKING order="16" place="16" resultid="4610" />
                    <RANKING order="17" place="17" resultid="3018" />
                    <RANKING order="18" place="18" resultid="4076" />
                    <RANKING order="19" place="19" resultid="4661" />
                    <RANKING order="20" place="20" resultid="4392" />
                    <RANKING order="21" place="21" resultid="3012" />
                    <RANKING order="22" place="22" resultid="2983" />
                    <RANKING order="23" place="23" resultid="2437" />
                    <RANKING order="24" place="24" resultid="3023" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6033" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2527" />
                    <RANKING order="2" place="2" resultid="2445" />
                    <RANKING order="3" place="3" resultid="3500" />
                    <RANKING order="4" place="4" resultid="3542" />
                    <RANKING order="5" place="5" resultid="3948" />
                    <RANKING order="6" place="6" resultid="4463" />
                    <RANKING order="7" place="7" resultid="3591" />
                    <RANKING order="8" place="8" resultid="2937" />
                    <RANKING order="9" place="9" resultid="2485" />
                    <RANKING order="10" place="10" resultid="4492" />
                    <RANKING order="11" place="11" resultid="2917" />
                    <RANKING order="12" place="12" resultid="2609" />
                    <RANKING order="13" place="13" resultid="4635" />
                    <RANKING order="14" place="14" resultid="4035" />
                    <RANKING order="15" place="15" resultid="2490" />
                    <RANKING order="16" place="16" resultid="2978" />
                    <RANKING order="17" place="17" resultid="2923" />
                    <RANKING order="18" place="18" resultid="4336" />
                    <RANKING order="19" place="19" resultid="3614" />
                    <RANKING order="20" place="20" resultid="4044" />
                    <RANKING order="21" place="21" resultid="3007" />
                    <RANKING order="22" place="22" resultid="3211" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6034" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3937" />
                    <RANKING order="2" place="2" resultid="3494" />
                    <RANKING order="3" place="3" resultid="3883" />
                    <RANKING order="4" place="4" resultid="3509" />
                    <RANKING order="5" place="5" resultid="3259" />
                    <RANKING order="6" place="5" resultid="4478" />
                    <RANKING order="7" place="7" resultid="3504" />
                    <RANKING order="8" place="8" resultid="3055" />
                    <RANKING order="9" place="9" resultid="3583" />
                    <RANKING order="10" place="10" resultid="3089" />
                    <RANKING order="11" place="11" resultid="2541" />
                    <RANKING order="12" place="12" resultid="3577" />
                    <RANKING order="13" place="13" resultid="2803" />
                    <RANKING order="14" place="14" resultid="4443" />
                    <RANKING order="15" place="15" resultid="3396" />
                    <RANKING order="16" place="16" resultid="2871" />
                    <RANKING order="17" place="17" resultid="4060" />
                    <RANKING order="18" place="18" resultid="3361" />
                    <RANKING order="19" place="19" resultid="2997" />
                    <RANKING order="20" place="20" resultid="3912" />
                    <RANKING order="21" place="21" resultid="4399" />
                    <RANKING order="22" place="22" resultid="3117" />
                    <RANKING order="23" place="23" resultid="3181" />
                    <RANKING order="24" place="24" resultid="3110" />
                    <RANKING order="25" place="25" resultid="2769" />
                    <RANKING order="26" place="26" resultid="4082" />
                    <RANKING order="27" place="27" resultid="4277" />
                    <RANKING order="28" place="-1" resultid="2988" />
                    <RANKING order="29" place="-1" resultid="2552" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6035" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3555" />
                    <RANKING order="2" place="2" resultid="4430" />
                    <RANKING order="3" place="3" resultid="4369" />
                    <RANKING order="4" place="4" resultid="4251" />
                    <RANKING order="5" place="5" resultid="4185" />
                    <RANKING order="6" place="6" resultid="4294" />
                    <RANKING order="7" place="7" resultid="4189" />
                    <RANKING order="8" place="8" resultid="4404" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6036" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3962" />
                    <RANKING order="2" place="2" resultid="3984" />
                    <RANKING order="3" place="3" resultid="4502" />
                    <RANKING order="4" place="4" resultid="3717" />
                    <RANKING order="5" place="5" resultid="4325" />
                    <RANKING order="6" place="6" resultid="4555" />
                    <RANKING order="7" place="7" resultid="2900" />
                    <RANKING order="8" place="8" resultid="2580" />
                    <RANKING order="9" place="9" resultid="3194" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6037" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3811" />
                    <RANKING order="2" place="2" resultid="2791" />
                    <RANKING order="3" place="3" resultid="3893" />
                    <RANKING order="4" place="4" resultid="2911" />
                    <RANKING order="5" place="-1" resultid="3049" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5217" daytime="09:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5218" daytime="09:36" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5219" daytime="09:38" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5220" daytime="09:42" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5221" daytime="09:44" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5222" daytime="09:46" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5223" daytime="09:48" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5224" daytime="09:52" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5225" daytime="09:54" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5226" daytime="09:56" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="5227" daytime="09:58" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="5228" daytime="10:00" number="12" order="12" status="OFFICIAL" />
                <HEAT heatid="5229" daytime="10:04" number="13" order="13" status="OFFICIAL" />
                <HEAT heatid="5230" daytime="10:06" number="14" order="14" status="OFFICIAL" />
                <HEAT heatid="5231" daytime="10:08" number="15" order="15" status="OFFICIAL" />
                <HEAT heatid="5232" daytime="10:10" number="16" order="16" status="OFFICIAL" />
                <HEAT heatid="5233" daytime="10:12" number="17" order="17" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1175" daytime="10:14" gender="F" number="15" order="3" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6038" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3798" />
                    <RANKING order="2" place="2" resultid="2659" />
                    <RANKING order="3" place="3" resultid="3334" />
                    <RANKING order="4" place="4" resultid="2513" />
                    <RANKING order="5" place="5" resultid="3842" />
                    <RANKING order="6" place="6" resultid="3924" />
                    <RANKING order="7" place="7" resultid="4172" />
                    <RANKING order="8" place="8" resultid="4244" />
                    <RANKING order="9" place="9" resultid="3001" />
                    <RANKING order="10" place="10" resultid="4568" />
                    <RANKING order="11" place="11" resultid="2763" />
                    <RANKING order="12" place="12" resultid="2632" />
                    <RANKING order="13" place="13" resultid="4178" />
                    <RANKING order="14" place="14" resultid="4627" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6039" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3277" />
                    <RANKING order="2" place="2" resultid="3384" />
                    <RANKING order="3" place="3" resultid="2416" />
                    <RANKING order="4" place="4" resultid="3655" />
                    <RANKING order="5" place="5" resultid="2726" />
                    <RANKING order="6" place="6" resultid="3641" />
                    <RANKING order="7" place="7" resultid="2639" />
                    <RANKING order="8" place="8" resultid="2423" />
                    <RANKING order="9" place="9" resultid="2827" />
                    <RANKING order="10" place="10" resultid="3662" />
                    <RANKING order="11" place="11" resultid="3158" />
                    <RANKING order="12" place="12" resultid="4648" />
                    <RANKING order="13" place="13" resultid="3431" />
                    <RANKING order="14" place="14" resultid="2497" />
                    <RANKING order="15" place="15" resultid="3837" />
                    <RANKING order="16" place="16" resultid="2751" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6040" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2877" />
                    <RANKING order="2" place="2" resultid="2466" />
                    <RANKING order="3" place="3" resultid="3610" />
                    <RANKING order="4" place="4" resultid="3284" />
                    <RANKING order="5" place="5" resultid="3263" />
                    <RANKING order="6" place="6" resultid="4484" />
                    <RANKING order="7" place="7" resultid="2592" />
                    <RANKING order="8" place="8" resultid="3102" />
                    <RANKING order="9" place="9" resultid="4380" />
                    <RANKING order="10" place="10" resultid="2478" />
                    <RANKING order="11" place="-1" resultid="2820" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6041" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3942" />
                    <RANKING order="2" place="2" resultid="3470" />
                    <RANKING order="3" place="3" resultid="2710" />
                    <RANKING order="4" place="4" resultid="2410" />
                    <RANKING order="5" place="5" resultid="2614" />
                    <RANKING order="6" place="6" resultid="2733" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6042" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2474" />
                    <RANKING order="2" place="2" resultid="4194" />
                    <RANKING order="3" place="3" resultid="2971" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6043" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2697" />
                    <RANKING order="2" place="2" resultid="2775" />
                    <RANKING order="3" place="3" resultid="4307" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6044" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5241" daytime="10:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5242" daytime="10:18" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5243" daytime="10:22" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5244" daytime="10:26" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5245" daytime="10:28" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5246" daytime="10:32" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5247" daytime="10:36" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5248" daytime="10:40" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1182" daytime="10:42" gender="M" number="16" order="4" round="PRE" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6045" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3312" />
                    <RANKING order="2" place="2" resultid="4129" />
                    <RANKING order="3" place="3" resultid="3829" />
                    <RANKING order="4" place="4" resultid="4521" />
                    <RANKING order="5" place="5" resultid="2745" />
                    <RANKING order="6" place="6" resultid="3793" />
                    <RANKING order="7" place="7" resultid="3403" />
                    <RANKING order="8" place="8" resultid="4143" />
                    <RANKING order="9" place="9" resultid="4345" />
                    <RANKING order="10" place="10" resultid="3723" />
                    <RANKING order="11" place="11" resultid="4200" />
                    <RANKING order="12" place="12" resultid="4101" />
                    <RANKING order="13" place="13" resultid="3804" />
                    <RANKING order="14" place="14" resultid="3767" />
                    <RANKING order="15" place="15" resultid="3130" />
                    <RANKING order="16" place="16" resultid="3753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6046" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2932" />
                    <RANKING order="2" place="2" resultid="3151" />
                    <RANKING order="3" place="3" resultid="3292" />
                    <RANKING order="4" place="4" resultid="3389" />
                    <RANKING order="5" place="5" resultid="3899" />
                    <RANKING order="6" place="6" resultid="3165" />
                    <RANKING order="7" place="7" resultid="3674" />
                    <RANKING order="8" place="8" resultid="3636" />
                    <RANKING order="9" place="9" resultid="3680" />
                    <RANKING order="10" place="10" resultid="4609" />
                    <RANKING order="11" place="11" resultid="2955" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6047" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3978" />
                    <RANKING order="2" place="2" resultid="2882" />
                    <RANKING order="3" place="3" resultid="3619" />
                    <RANKING order="4" place="4" resultid="4300" />
                    <RANKING order="5" place="5" resultid="4602" />
                    <RANKING order="6" place="6" resultid="4457" />
                    <RANKING order="7" place="7" resultid="3354" />
                    <RANKING order="8" place="8" resultid="4122" />
                    <RANKING order="9" place="-1" resultid="3586" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6048" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3488" />
                    <RANKING order="2" place="2" resultid="3625" />
                    <RANKING order="3" place="3" resultid="3936" />
                    <RANKING order="4" place="4" resultid="3571" />
                    <RANKING order="5" place="5" resultid="3566" />
                    <RANKING order="6" place="6" resultid="2540" />
                    <RANKING order="7" place="7" resultid="4150" />
                    <RANKING order="8" place="8" resultid="3870" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6049" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3967" />
                    <RANKING order="2" place="2" resultid="2402" />
                    <RANKING order="3" place="3" resultid="4184" />
                    <RANKING order="4" place="4" resultid="3305" />
                    <RANKING order="5" place="5" resultid="4368" />
                    <RANKING order="6" place="-1" resultid="4064" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6050" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3481" />
                    <RANKING order="2" place="2" resultid="4501" />
                    <RANKING order="3" place="3" resultid="3082" />
                    <RANKING order="4" place="4" resultid="3068" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6051" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3810" />
                    <RANKING order="2" place="2" resultid="2786" />
                    <RANKING order="3" place="3" resultid="3061" />
                    <RANKING order="4" place="4" resultid="3238" />
                    <RANKING order="5" place="5" resultid="3075" />
                    <RANKING order="6" place="-1" resultid="2894" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5255" daytime="10:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5256" daytime="10:46" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5257" daytime="10:50" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5258" daytime="10:52" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5259" daytime="10:56" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5260" daytime="10:58" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5261" daytime="11:02" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5262" daytime="11:06" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5263" daytime="11:08" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1190" daytime="11:12" gender="F" number="17" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6222" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3340" />
                    <RANKING order="2" place="2" resultid="3799" />
                    <RANKING order="3" place="3" resultid="3411" />
                    <RANKING order="4" place="4" resultid="3760" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6223" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3700" />
                    <RANKING order="2" place="2" resultid="3687" />
                    <RANKING order="3" place="3" resultid="4319" />
                    <RANKING order="4" place="-1" resultid="3138" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6224" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3464" />
                    <RANKING order="2" place="2" resultid="4471" />
                    <RANKING order="3" place="-1" resultid="3526" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6225" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3040" />
                    <RANKING order="2" place="2" resultid="2867" />
                    <RANKING order="3" place="3" resultid="2797" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6226" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3549" />
                    <RANKING order="2" place="2" resultid="3250" />
                    <RANKING order="3" place="3" resultid="4195" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6227" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6228" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3906" />
                    <RANKING order="2" place="2" resultid="3917" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6229" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3906" />
                    <RANKING order="2" place="2" resultid="3917" />
                    <RANKING order="3" place="3" resultid="3549" />
                    <RANKING order="4" place="4" resultid="3464" />
                    <RANKING order="5" place="5" resultid="3700" />
                    <RANKING order="6" place="6" resultid="3687" />
                    <RANKING order="7" place="7" resultid="3250" />
                    <RANKING order="8" place="8" resultid="4437" />
                    <RANKING order="9" place="9" resultid="3340" />
                    <RANKING order="10" place="10" resultid="3040" />
                    <RANKING order="11" place="11" resultid="4319" />
                    <RANKING order="12" place="12" resultid="2867" />
                    <RANKING order="13" place="13" resultid="4195" />
                    <RANKING order="14" place="14" resultid="3799" />
                    <RANKING order="15" place="15" resultid="3411" />
                    <RANKING order="16" place="16" resultid="2797" />
                    <RANKING order="17" place="17" resultid="4471" />
                    <RANKING order="18" place="18" resultid="3760" />
                    <RANKING order="19" place="-1" resultid="3138" />
                    <RANKING order="20" place="-1" resultid="3526" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5271" daytime="11:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5272" daytime="11:24" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5273" daytime="11:36" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2320" daytime="11:52" gender="M" number="4" order="6" round="FIN" preveventid="1088">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6374" agemax="-1" agemin="13" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5953" />
                    <RANKING order="2" place="2" resultid="5954" />
                    <RANKING order="3" place="3" resultid="5955" />
                    <RANKING order="4" place="4" resultid="5957" />
                    <RANKING order="5" place="5" resultid="5956" />
                    <RANKING order="6" place="6" resultid="5959" />
                    <RANKING order="7" place="7" resultid="5958" />
                    <RANKING order="8" place="8" resultid="5960" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6414" agegroupid="6374" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2312" daytime="11:48" gender="F" number="3" order="7" round="FIN" preveventid="1080">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6373" agemax="-1" agemin="13" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5938" />
                    <RANKING order="2" place="2" resultid="5939" />
                    <RANKING order="3" place="3" resultid="5940" />
                    <RANKING order="4" place="4" resultid="5943" />
                    <RANKING order="5" place="5" resultid="5942" />
                    <RANKING order="6" place="6" resultid="5945" />
                    <RANKING order="7" place="7" resultid="5944" />
                    <RANKING order="8" place="8" resultid="5946" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6416" agegroupid="6373" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-09-20" daytime="16:10" endtime="20:14" number="4" officialmeeting="15:30" teamleadermeeting="16:00" warmupfrom="15:00" warmupuntil="16:00">
          <EVENTS>
            <EVENT eventid="2335" daytime="16:10" gender="M" number="10" order="1" round="FIN" preveventid="1135">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6372" agemax="-1" agemin="13" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6008" />
                    <RANKING order="2" place="2" resultid="6009" />
                    <RANKING order="3" place="3" resultid="6010" />
                    <RANKING order="4" place="4" resultid="6015" />
                    <RANKING order="5" place="5" resultid="6013" />
                    <RANKING order="6" place="6" resultid="6011" />
                    <RANKING order="7" place="7" resultid="6012" />
                    <RANKING order="8" place="8" resultid="6014" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6417" agegroupid="6372" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2328" daytime="16:12" gender="F" number="9" order="2" round="FIN" preveventid="1128">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6371" agemax="-1" agemin="13" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5998" />
                    <RANKING order="2" place="2" resultid="5997" />
                    <RANKING order="3" place="3" resultid="5999" />
                    <RANKING order="4" place="4" resultid="6002" />
                    <RANKING order="5" place="5" resultid="6000" />
                    <RANKING order="6" place="6" resultid="6004" />
                    <RANKING order="7" place="7" resultid="6003" />
                    <RANKING order="8" place="8" resultid="6001" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6418" agegroupid="6371" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1198" daytime="16:16" gender="M" number="18" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6230" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3313" />
                    <RANKING order="2" place="2" resultid="3737" />
                    <RANKING order="3" place="3" resultid="4522" />
                    <RANKING order="4" place="4" resultid="3348" />
                    <RANKING order="5" place="5" resultid="3404" />
                    <RANKING order="6" place="6" resultid="3768" />
                    <RANKING order="7" place="7" resultid="3805" />
                    <RANKING order="8" place="8" resultid="3417" />
                    <RANKING order="9" place="9" resultid="4135" />
                    <RANKING order="10" place="10" resultid="3369" />
                    <RANKING order="11" place="11" resultid="2626" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6231" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3390" />
                    <RANKING order="2" place="2" resultid="2933" />
                    <RANKING order="3" place="3" resultid="3439" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6232" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3270" />
                    <RANKING order="2" place="2" resultid="2452" />
                    <RANKING order="3" place="3" resultid="4257" />
                    <RANKING order="4" place="4" resultid="3355" />
                    <RANKING order="5" place="-1" resultid="4301" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6233" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3495" />
                    <RANKING order="2" place="2" resultid="3397" />
                    <RANKING order="3" place="3" resultid="3572" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6234" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3521" />
                    <RANKING order="2" place="2" resultid="3306" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6235" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3069" />
                    <RANKING order="2" place="2" resultid="3718" />
                    <RANKING order="3" place="3" resultid="2581" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6236" agemax="-1" agemin="20" />
                <AGEGROUP agegroupid="6237" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3521" />
                    <RANKING order="2" place="2" resultid="3495" />
                    <RANKING order="3" place="3" resultid="3270" />
                    <RANKING order="4" place="4" resultid="2452" />
                    <RANKING order="5" place="5" resultid="4257" />
                    <RANKING order="6" place="6" resultid="3355" />
                    <RANKING order="7" place="7" resultid="3069" />
                    <RANKING order="8" place="8" resultid="3306" />
                    <RANKING order="9" place="9" resultid="3397" />
                    <RANKING order="10" place="10" resultid="3313" />
                    <RANKING order="11" place="11" resultid="3390" />
                    <RANKING order="12" place="12" resultid="2933" />
                    <RANKING order="13" place="13" resultid="3572" />
                    <RANKING order="14" place="14" resultid="3737" />
                    <RANKING order="15" place="15" resultid="3718" />
                    <RANKING order="16" place="16" resultid="4522" />
                    <RANKING order="17" place="17" resultid="3439" />
                    <RANKING order="18" place="18" resultid="3348" />
                    <RANKING order="19" place="19" resultid="3404" />
                    <RANKING order="20" place="20" resultid="3768" />
                    <RANKING order="21" place="21" resultid="3805" />
                    <RANKING order="22" place="22" resultid="2581" />
                    <RANKING order="23" place="23" resultid="3417" />
                    <RANKING order="24" place="24" resultid="4135" />
                    <RANKING order="25" place="25" resultid="3369" />
                    <RANKING order="26" place="26" resultid="2626" />
                    <RANKING order="27" place="-1" resultid="4301" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5274" daytime="16:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5275" daytime="16:22" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5276" daytime="16:30" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5277" daytime="16:38" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1205" daytime="16:44" gender="F" number="19" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6238" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3853" />
                    <RANKING order="2" place="2" resultid="3335" />
                    <RANKING order="3" place="3" resultid="3424" />
                    <RANKING order="4" place="4" resultid="3376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6239" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3278" />
                    <RANKING order="2" place="2" resultid="4264" />
                    <RANKING order="3" place="3" resultid="4590" />
                    <RANKING order="4" place="4" resultid="4320" />
                    <RANKING order="5" place="5" resultid="2648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6240" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3285" />
                    <RANKING order="2" place="-1" resultid="3465" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6241" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3320" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6242" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4196" />
                    <RANKING order="2" place="2" resultid="3251" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6243" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4308" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6244" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3907" />
                    <RANKING order="2" place="2" resultid="3918" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6245" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3907" />
                    <RANKING order="2" place="2" resultid="3918" />
                    <RANKING order="3" place="3" resultid="3853" />
                    <RANKING order="4" place="4" resultid="3320" />
                    <RANKING order="5" place="5" resultid="3278" />
                    <RANKING order="6" place="6" resultid="3335" />
                    <RANKING order="7" place="7" resultid="4264" />
                    <RANKING order="8" place="8" resultid="3424" />
                    <RANKING order="9" place="9" resultid="4196" />
                    <RANKING order="10" place="10" resultid="4590" />
                    <RANKING order="11" place="11" resultid="3251" />
                    <RANKING order="12" place="12" resultid="3376" />
                    <RANKING order="13" place="13" resultid="4320" />
                    <RANKING order="14" place="14" resultid="2648" />
                    <RANKING order="15" place="15" resultid="4308" />
                    <RANKING order="16" place="-1" resultid="3285" />
                    <RANKING order="17" place="-1" resultid="3465" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5278" daytime="16:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5279" daytime="16:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5280" daytime="17:00" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1213" daytime="17:08" gender="M" number="20" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6246" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2621" />
                    <RANKING order="2" place="2" resultid="4523" />
                    <RANKING order="3" place="3" resultid="2747" />
                    <RANKING order="4" place="4" resultid="2835" />
                    <RANKING order="5" place="5" resultid="4201" />
                    <RANKING order="6" place="6" resultid="4346" />
                    <RANKING order="7" place="7" resultid="2757" />
                    <RANKING order="8" place="8" resultid="3131" />
                    <RANKING order="9" place="9" resultid="2654" />
                    <RANKING order="10" place="10" resultid="2843" />
                    <RANKING order="11" place="11" resultid="2856" />
                    <RANKING order="12" place="12" resultid="4109" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6247" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3167" />
                    <RANKING order="2" place="2" resultid="3901" />
                    <RANKING order="3" place="3" resultid="3152" />
                    <RANKING order="4" place="4" resultid="3676" />
                    <RANKING order="5" place="5" resultid="3391" />
                    <RANKING order="6" place="6" resultid="3637" />
                    <RANKING order="7" place="7" resultid="3819" />
                    <RANKING order="8" place="8" resultid="4611" />
                    <RANKING order="9" place="9" resultid="2956" />
                    <RANKING order="10" place="10" resultid="3019" />
                    <RANKING order="11" place="11" resultid="2438" />
                    <RANKING order="12" place="12" resultid="4164" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6248" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3979" />
                    <RANKING order="2" place="2" resultid="2446" />
                    <RANKING order="3" place="3" resultid="4302" />
                    <RANKING order="4" place="4" resultid="4458" />
                    <RANKING order="5" place="5" resultid="4464" />
                    <RANKING order="6" place="6" resultid="2938" />
                    <RANKING order="7" place="7" resultid="4036" />
                    <RANKING order="8" place="7" resultid="4493" />
                    <RANKING order="9" place="9" resultid="3008" />
                    <RANKING order="10" place="-1" resultid="2883" />
                    <RANKING order="11" place="-1" resultid="4045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6249" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3489" />
                    <RANKING order="2" place="2" resultid="2603" />
                    <RANKING order="3" place="3" resultid="3260" />
                    <RANKING order="4" place="4" resultid="2542" />
                    <RANKING order="5" place="5" resultid="2872" />
                    <RANKING order="6" place="6" resultid="3056" />
                    <RANKING order="7" place="7" resultid="4444" />
                    <RANKING order="8" place="8" resultid="2770" />
                    <RANKING order="9" place="9" resultid="4479" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6250" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3968" />
                    <RANKING order="2" place="2" resultid="4295" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6251" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2814" />
                    <RANKING order="2" place="-1" resultid="3482" />
                    <RANKING order="3" place="-1" resultid="3985" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6252" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3812" />
                    <RANKING order="2" place="2" resultid="2565" />
                    <RANKING order="3" place="3" resultid="2787" />
                    <RANKING order="4" place="4" resultid="2782" />
                    <RANKING order="5" place="5" resultid="3894" />
                    <RANKING order="6" place="6" resultid="3062" />
                    <RANKING order="7" place="7" resultid="3239" />
                    <RANKING order="8" place="8" resultid="3076" />
                    <RANKING order="9" place="9" resultid="2792" />
                    <RANKING order="10" place="10" resultid="2895" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6253" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3812" />
                    <RANKING order="2" place="2" resultid="2565" />
                    <RANKING order="3" place="3" resultid="3979" />
                    <RANKING order="4" place="4" resultid="2787" />
                    <RANKING order="5" place="5" resultid="3968" />
                    <RANKING order="6" place="6" resultid="3489" />
                    <RANKING order="7" place="7" resultid="2446" />
                    <RANKING order="8" place="8" resultid="2782" />
                    <RANKING order="9" place="9" resultid="3894" />
                    <RANKING order="10" place="10" resultid="3062" />
                    <RANKING order="11" place="11" resultid="3239" />
                    <RANKING order="12" place="12" resultid="4302" />
                    <RANKING order="13" place="13" resultid="4458" />
                    <RANKING order="14" place="14" resultid="4464" />
                    <RANKING order="15" place="15" resultid="2938" />
                    <RANKING order="16" place="16" resultid="2603" />
                    <RANKING order="17" place="17" resultid="3260" />
                    <RANKING order="18" place="18" resultid="3076" />
                    <RANKING order="19" place="19" resultid="3167" />
                    <RANKING order="20" place="20" resultid="2542" />
                    <RANKING order="21" place="21" resultid="3901" />
                    <RANKING order="22" place="22" resultid="3152" />
                    <RANKING order="23" place="23" resultid="2872" />
                    <RANKING order="24" place="24" resultid="3056" />
                    <RANKING order="25" place="24" resultid="3676" />
                    <RANKING order="26" place="26" resultid="4444" />
                    <RANKING order="27" place="27" resultid="2621" />
                    <RANKING order="28" place="28" resultid="2792" />
                    <RANKING order="29" place="29" resultid="2770" />
                    <RANKING order="30" place="30" resultid="4523" />
                    <RANKING order="31" place="31" resultid="3391" />
                    <RANKING order="32" place="32" resultid="2747" />
                    <RANKING order="33" place="33" resultid="2814" />
                    <RANKING order="34" place="34" resultid="4479" />
                    <RANKING order="35" place="35" resultid="4036" />
                    <RANKING order="36" place="35" resultid="4493" />
                    <RANKING order="37" place="37" resultid="2895" />
                    <RANKING order="38" place="38" resultid="3637" />
                    <RANKING order="39" place="39" resultid="3819" />
                    <RANKING order="40" place="40" resultid="4611" />
                    <RANKING order="41" place="41" resultid="2956" />
                    <RANKING order="42" place="42" resultid="2835" />
                    <RANKING order="43" place="43" resultid="4201" />
                    <RANKING order="44" place="44" resultid="3019" />
                    <RANKING order="45" place="45" resultid="4346" />
                    <RANKING order="46" place="46" resultid="4295" />
                    <RANKING order="47" place="47" resultid="2757" />
                    <RANKING order="48" place="48" resultid="2438" />
                    <RANKING order="49" place="49" resultid="4164" />
                    <RANKING order="50" place="50" resultid="3131" />
                    <RANKING order="51" place="51" resultid="2654" />
                    <RANKING order="52" place="52" resultid="2843" />
                    <RANKING order="53" place="53" resultid="3008" />
                    <RANKING order="54" place="54" resultid="2856" />
                    <RANKING order="55" place="55" resultid="4109" />
                    <RANKING order="56" place="-1" resultid="3482" />
                    <RANKING order="57" place="-1" resultid="2883" />
                    <RANKING order="58" place="-1" resultid="3985" />
                    <RANKING order="59" place="-1" resultid="4045" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5281" daytime="17:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5282" daytime="17:10" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5283" daytime="17:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5284" daytime="17:16" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5285" daytime="17:18" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5286" daytime="17:22" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5287" daytime="17:24" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5288" daytime="17:26" number="8" order="8" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1215" daytime="17:28" gender="F" number="21" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6254" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2660" />
                    <RANKING order="2" place="2" resultid="2514" />
                    <RANKING order="3" place="3" resultid="3926" />
                    <RANKING order="4" place="4" resultid="3412" />
                    <RANKING order="5" place="5" resultid="3341" />
                    <RANKING order="6" place="6" resultid="4246" />
                    <RANKING order="7" place="7" resultid="2634" />
                    <RANKING order="8" place="8" resultid="3002" />
                    <RANKING order="9" place="9" resultid="2671" />
                    <RANKING order="10" place="10" resultid="4179" />
                    <RANKING order="11" place="10" resultid="4569" />
                    <RANKING order="12" place="12" resultid="2765" />
                    <RANKING order="13" place="13" resultid="2740" />
                    <RANKING order="14" place="14" resultid="3125" />
                    <RANKING order="15" place="-1" resultid="3199" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6255" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2728" />
                    <RANKING order="2" place="2" resultid="3279" />
                    <RANKING order="3" place="3" resultid="2418" />
                    <RANKING order="4" place="4" resultid="2640" />
                    <RANKING order="5" place="5" resultid="3643" />
                    <RANKING order="6" place="6" resultid="2425" />
                    <RANKING order="7" place="7" resultid="3139" />
                    <RANKING order="8" place="8" resultid="3159" />
                    <RANKING order="9" place="9" resultid="2828" />
                    <RANKING order="10" place="10" resultid="4642" />
                    <RANKING order="11" place="11" resultid="3433" />
                    <RANKING order="12" place="12" resultid="4649" />
                    <RANKING order="13" place="13" resultid="2499" />
                    <RANKING order="14" place="14" resultid="4353" />
                    <RANKING order="15" place="15" resultid="2753" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6256" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2878" />
                    <RANKING order="2" place="2" resultid="2467" />
                    <RANKING order="3" place="3" resultid="4486" />
                    <RANKING order="4" place="4" resultid="3264" />
                    <RANKING order="5" place="5" resultid="3611" />
                    <RANKING order="6" place="6" resultid="2593" />
                    <RANKING order="7" place="7" resultid="4158" />
                    <RANKING order="8" place="8" resultid="2479" />
                    <RANKING order="9" place="9" resultid="3104" />
                    <RANKING order="10" place="10" resultid="2822" />
                    <RANKING order="11" place="11" resultid="4510" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6257" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3943" />
                    <RANKING order="2" place="2" resultid="4375" />
                    <RANKING order="3" place="3" resultid="2798" />
                    <RANKING order="4" place="4" resultid="2587" />
                    <RANKING order="5" place="5" resultid="2615" />
                    <RANKING order="6" place="6" resultid="2735" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6258" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2475" />
                    <RANKING order="2" place="2" resultid="2471" />
                    <RANKING order="3" place="3" resultid="2972" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6259" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2699" />
                    <RANKING order="2" place="2" resultid="2777" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6260" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4288" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6261" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3943" />
                    <RANKING order="2" place="2" resultid="2699" />
                    <RANKING order="3" place="3" resultid="2777" />
                    <RANKING order="4" place="4" resultid="2878" />
                    <RANKING order="5" place="5" resultid="2475" />
                    <RANKING order="6" place="6" resultid="2467" />
                    <RANKING order="7" place="7" resultid="2660" />
                    <RANKING order="8" place="8" resultid="2728" />
                    <RANKING order="9" place="9" resultid="3279" />
                    <RANKING order="10" place="10" resultid="2418" />
                    <RANKING order="11" place="11" resultid="4375" />
                    <RANKING order="12" place="12" resultid="2640" />
                    <RANKING order="13" place="13" resultid="4486" />
                    <RANKING order="14" place="14" resultid="2514" />
                    <RANKING order="15" place="15" resultid="3643" />
                    <RANKING order="16" place="16" resultid="2425" />
                    <RANKING order="17" place="17" resultid="3264" />
                    <RANKING order="18" place="18" resultid="3611" />
                    <RANKING order="19" place="19" resultid="2593" />
                    <RANKING order="20" place="20" resultid="4158" />
                    <RANKING order="21" place="21" resultid="3139" />
                    <RANKING order="22" place="22" resultid="3926" />
                    <RANKING order="23" place="23" resultid="2798" />
                    <RANKING order="24" place="24" resultid="2587" />
                    <RANKING order="25" place="25" resultid="2471" />
                    <RANKING order="26" place="26" resultid="2479" />
                    <RANKING order="27" place="27" resultid="3159" />
                    <RANKING order="28" place="28" resultid="2828" />
                    <RANKING order="29" place="29" resultid="2615" />
                    <RANKING order="30" place="30" resultid="3412" />
                    <RANKING order="31" place="31" resultid="4642" />
                    <RANKING order="32" place="32" resultid="3433" />
                    <RANKING order="33" place="33" resultid="3104" />
                    <RANKING order="34" place="34" resultid="2822" />
                    <RANKING order="35" place="35" resultid="3341" />
                    <RANKING order="36" place="36" resultid="4246" />
                    <RANKING order="37" place="37" resultid="4510" />
                    <RANKING order="38" place="38" resultid="4649" />
                    <RANKING order="39" place="39" resultid="2634" />
                    <RANKING order="40" place="40" resultid="4288" />
                    <RANKING order="41" place="41" resultid="2499" />
                    <RANKING order="42" place="42" resultid="3002" />
                    <RANKING order="43" place="43" resultid="2671" />
                    <RANKING order="44" place="44" resultid="2735" />
                    <RANKING order="45" place="45" resultid="4179" />
                    <RANKING order="46" place="45" resultid="4569" />
                    <RANKING order="47" place="47" resultid="2765" />
                    <RANKING order="48" place="48" resultid="2972" />
                    <RANKING order="49" place="49" resultid="4353" />
                    <RANKING order="50" place="50" resultid="2740" />
                    <RANKING order="51" place="51" resultid="2753" />
                    <RANKING order="52" place="52" resultid="3125" />
                    <RANKING order="53" place="-1" resultid="3199" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5289" daytime="17:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5290" daytime="17:32" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5291" daytime="17:34" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5292" daytime="17:38" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5293" daytime="17:40" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5294" daytime="17:42" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5295" daytime="17:46" number="7" order="7" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1217" daytime="17:48" gender="M" number="22" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6262" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3327" />
                    <RANKING order="2" place="2" resultid="3724" />
                    <RANKING order="3" place="3" resultid="4347" />
                    <RANKING order="4" place="4" resultid="3206" />
                    <RANKING order="5" place="5" resultid="4564" />
                    <RANKING order="6" place="6" resultid="4576" />
                    <RANKING order="7" place="7" resultid="3864" />
                    <RANKING order="8" place="8" resultid="3223" />
                    <RANKING order="9" place="9" resultid="4102" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6263" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3669" />
                    <RANKING order="2" place="2" resultid="3293" />
                    <RANKING order="3" place="3" resultid="3681" />
                    <RANKING order="4" place="4" resultid="4596" />
                    <RANKING order="5" place="5" resultid="4271" />
                    <RANKING order="6" place="6" resultid="2678" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6264" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3271" />
                    <RANKING order="2" place="2" resultid="3543" />
                    <RANKING order="3" place="3" resultid="4258" />
                    <RANKING order="4" place="4" resultid="3620" />
                    <RANKING order="5" place="5" resultid="4123" />
                    <RANKING order="6" place="6" resultid="4337" />
                    <RANKING order="7" place="7" resultid="2491" />
                    <RANKING order="8" place="-1" resultid="3587" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6265" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3090" />
                    <RANKING order="2" place="2" resultid="3362" />
                    <RANKING order="3" place="3" resultid="3111" />
                    <RANKING order="4" place="4" resultid="4312" />
                    <RANKING order="5" place="5" resultid="3118" />
                    <RANKING order="6" place="6" resultid="3182" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6266" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3556" />
                    <RANKING order="2" place="2" resultid="3096" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6267" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3963" />
                    <RANKING order="2" place="2" resultid="4503" />
                    <RANKING order="3" place="3" resultid="3245" />
                    <RANKING order="4" place="4" resultid="3083" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6268" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2904" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6269" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3963" />
                    <RANKING order="2" place="2" resultid="3556" />
                    <RANKING order="3" place="3" resultid="3669" />
                    <RANKING order="4" place="4" resultid="3271" />
                    <RANKING order="5" place="5" resultid="4503" />
                    <RANKING order="6" place="6" resultid="3543" />
                    <RANKING order="7" place="7" resultid="4258" />
                    <RANKING order="8" place="8" resultid="3620" />
                    <RANKING order="9" place="9" resultid="3293" />
                    <RANKING order="10" place="10" resultid="3090" />
                    <RANKING order="11" place="11" resultid="3681" />
                    <RANKING order="12" place="12" resultid="3245" />
                    <RANKING order="13" place="13" resultid="3362" />
                    <RANKING order="14" place="14" resultid="3083" />
                    <RANKING order="15" place="15" resultid="3327" />
                    <RANKING order="16" place="16" resultid="3724" />
                    <RANKING order="17" place="17" resultid="3111" />
                    <RANKING order="18" place="18" resultid="4123" />
                    <RANKING order="19" place="19" resultid="4347" />
                    <RANKING order="20" place="20" resultid="4596" />
                    <RANKING order="21" place="21" resultid="3096" />
                    <RANKING order="22" place="22" resultid="4337" />
                    <RANKING order="23" place="23" resultid="3206" />
                    <RANKING order="24" place="24" resultid="4564" />
                    <RANKING order="25" place="25" resultid="4312" />
                    <RANKING order="26" place="26" resultid="2491" />
                    <RANKING order="27" place="27" resultid="4271" />
                    <RANKING order="28" place="28" resultid="2904" />
                    <RANKING order="29" place="29" resultid="3118" />
                    <RANKING order="30" place="30" resultid="4576" />
                    <RANKING order="31" place="31" resultid="3864" />
                    <RANKING order="32" place="32" resultid="2678" />
                    <RANKING order="33" place="33" resultid="3182" />
                    <RANKING order="34" place="34" resultid="3223" />
                    <RANKING order="35" place="35" resultid="4102" />
                    <RANKING order="36" place="-1" resultid="3587" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5296" daytime="17:48" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5297" daytime="18:00" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5298" daytime="18:14" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5299" daytime="18:26" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5300" daytime="18:38" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1219" daytime="18:48" gender="F" number="23" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1220" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3989" />
                    <RANKING order="2" place="2" resultid="4013" />
                    <RANKING order="3" place="3" resultid="3444" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5301" daytime="18:48" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1221" daytime="18:56" gender="F" number="24" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1222" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3988" />
                    <RANKING order="2" place="2" resultid="3443" />
                    <RANKING order="3" place="3" resultid="4012" />
                    <RANKING order="4" place="4" resultid="4669" />
                    <RANKING order="5" place="5" resultid="2681" />
                    <RANKING order="6" place="6" resultid="2519" />
                    <RANKING order="7" place="7" resultid="4406" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5302" daytime="18:56" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1223" daytime="19:02" gender="F" number="25" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1224" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3987" />
                    <RANKING order="2" place="2" resultid="4668" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5303" daytime="19:02" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1225" daytime="19:08" gender="F" number="26" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1226" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3990" />
                    <RANKING order="2" place="2" resultid="3025" />
                    <RANKING order="3" place="3" resultid="2682" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5304" daytime="19:08" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1227" daytime="19:14" gender="F" number="27" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1228" agemax="19" agemin="17" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1229" daytime="19:14" gender="F" number="28" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1230" agemax="-1" agemin="20" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1231" daytime="19:14" gender="M" number="29" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1232" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3999" />
                    <RANKING order="2" place="2" resultid="3449" />
                    <RANKING order="3" place="3" resultid="4673" />
                    <RANKING order="4" place="4" resultid="2686" />
                    <RANKING order="5" place="5" resultid="4018" />
                    <RANKING order="6" place="6" resultid="2860" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5305" daytime="19:14" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1233" daytime="19:20" gender="M" number="30" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1234" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3998" />
                    <RANKING order="2" place="2" resultid="4017" />
                    <RANKING order="3" place="3" resultid="3448" />
                    <RANKING order="4" place="4" resultid="4672" />
                    <RANKING order="5" place="5" resultid="3171" />
                    <RANKING order="6" place="6" resultid="4410" />
                    <RANKING order="7" place="7" resultid="3029" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5306" daytime="19:20" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1235" daytime="19:26" gender="M" number="31" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1236" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3997" />
                    <RANKING order="2" place="2" resultid="2520" />
                    <RANKING order="3" place="3" resultid="3028" />
                    <RANKING order="4" place="4" resultid="4671" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5307" daytime="19:26" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1237" daytime="19:32" gender="M" number="32" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1238" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3995" />
                    <RANKING order="2" place="2" resultid="3447" />
                    <RANKING order="3" place="3" resultid="3169" />
                    <RANKING order="4" place="4" resultid="2685" />
                    <RANKING order="5" place="5" resultid="4408" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5308" daytime="19:32" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1239" daytime="19:38" gender="M" number="33" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1240" agemax="19" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4016" />
                    <RANKING order="2" place="2" resultid="3996" />
                    <RANKING order="3" place="3" resultid="4409" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5309" daytime="19:38" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1241" daytime="19:42" gender="M" number="34" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="FREE" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1242" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2859" />
                    <RANKING order="2" place="2" resultid="3170" />
                    <RANKING order="3" place="3" resultid="3027" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5310" daytime="19:42" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-09-21" daytime="09:10" endtime="13:02" number="5" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="2343" daytime="09:10" gender="F" number="13" order="1" round="FIN" preveventid="1159">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6370" agemax="-1" agemin="13" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6101" />
                    <RANKING order="2" place="2" resultid="6102" />
                    <RANKING order="3" place="3" resultid="6103" />
                    <RANKING order="4" place="4" resultid="6107" />
                    <RANKING order="5" place="5" resultid="6105" />
                    <RANKING order="6" place="6" resultid="6104" />
                    <RANKING order="7" place="7" resultid="6108" />
                    <RANKING order="8" place="8" resultid="6106" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6421" agegroupid="6370" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2351" daytime="09:12" gender="M" number="14" order="2" round="FIN" preveventid="1167">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6369" agemax="-1" agemin="13" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6116" />
                    <RANKING order="2" place="2" resultid="6118" />
                    <RANKING order="3" place="3" resultid="6117" />
                    <RANKING order="4" place="4" resultid="6119" />
                    <RANKING order="5" place="5" resultid="6121" />
                    <RANKING order="6" place="6" resultid="6120" />
                    <RANKING order="7" place="7" resultid="6122" />
                    <RANKING order="8" place="8" resultid="6123" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6422" agegroupid="6369" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1243" daytime="09:14" gender="F" number="35" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6270" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3854" />
                    <RANKING order="2" place="2" resultid="3748" />
                    <RANKING order="3" place="3" resultid="3377" />
                    <RANKING order="4" place="4" resultid="3774" />
                    <RANKING order="5" place="5" resultid="3932" />
                    <RANKING order="6" place="6" resultid="3426" />
                    <RANKING order="7" place="7" resultid="4570" />
                    <RANKING order="8" place="8" resultid="4517" />
                    <RANKING order="9" place="9" resultid="2672" />
                    <RANKING order="10" place="10" resultid="4117" />
                    <RANKING order="11" place="-1" resultid="3761" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6271" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3385" />
                    <RANKING order="2" place="2" resultid="3533" />
                    <RANKING order="3" place="3" resultid="4583" />
                    <RANKING order="4" place="4" resultid="4265" />
                    <RANKING order="5" place="5" resultid="4591" />
                    <RANKING order="6" place="-1" resultid="3888" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6272" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3595" />
                    <RANKING order="2" place="2" resultid="2944" />
                    <RANKING order="3" place="3" resultid="3600" />
                    <RANKING order="4" place="4" resultid="3537" />
                    <RANKING order="5" place="5" resultid="3286" />
                    <RANKING order="6" place="6" resultid="2480" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6273" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3460" />
                    <RANKING order="2" place="2" resultid="3847" />
                    <RANKING order="3" place="3" resultid="2716" />
                    <RANKING order="4" place="4" resultid="2411" />
                    <RANKING order="5" place="5" resultid="4451" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6274" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2967" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6275" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3956" />
                    <RANKING order="2" place="2" resultid="2461" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6276" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4029" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6277" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3956" />
                    <RANKING order="2" place="2" resultid="3460" />
                    <RANKING order="3" place="3" resultid="3595" />
                    <RANKING order="4" place="4" resultid="3847" />
                    <RANKING order="5" place="5" resultid="3385" />
                    <RANKING order="6" place="6" resultid="3854" />
                    <RANKING order="7" place="7" resultid="2944" />
                    <RANKING order="8" place="8" resultid="4029" />
                    <RANKING order="9" place="9" resultid="3748" />
                    <RANKING order="10" place="10" resultid="2461" />
                    <RANKING order="11" place="11" resultid="3533" />
                    <RANKING order="12" place="12" resultid="3600" />
                    <RANKING order="13" place="13" resultid="4583" />
                    <RANKING order="14" place="14" resultid="3537" />
                    <RANKING order="15" place="15" resultid="4265" />
                    <RANKING order="16" place="16" resultid="3377" />
                    <RANKING order="17" place="17" resultid="3774" />
                    <RANKING order="18" place="18" resultid="4591" />
                    <RANKING order="19" place="19" resultid="2716" />
                    <RANKING order="20" place="20" resultid="3932" />
                    <RANKING order="21" place="21" resultid="3286" />
                    <RANKING order="22" place="22" resultid="3426" />
                    <RANKING order="23" place="23" resultid="4570" />
                    <RANKING order="24" place="24" resultid="2411" />
                    <RANKING order="25" place="25" resultid="4517" />
                    <RANKING order="26" place="26" resultid="2672" />
                    <RANKING order="27" place="27" resultid="2480" />
                    <RANKING order="28" place="28" resultid="4117" />
                    <RANKING order="29" place="29" resultid="4451" />
                    <RANKING order="30" place="30" resultid="2967" />
                    <RANKING order="31" place="-1" resultid="3761" />
                    <RANKING order="32" place="-1" resultid="3888" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5311" daytime="09:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5312" daytime="09:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5313" daytime="09:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5314" daytime="09:28" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1251" daytime="09:34" gender="M" number="36" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6278" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3738" />
                    <RANKING order="2" place="2" resultid="3419" />
                    <RANKING order="3" place="3" resultid="3349" />
                    <RANKING order="4" place="4" resultid="3787" />
                    <RANKING order="5" place="5" resultid="4386" />
                    <RANKING order="6" place="6" resultid="3865" />
                    <RANKING order="7" place="7" resultid="3370" />
                    <RANKING order="8" place="8" resultid="3806" />
                    <RANKING order="9" place="9" resultid="2559" />
                    <RANKING order="10" place="10" resultid="4537" />
                    <RANKING order="11" place="11" resultid="3405" />
                    <RANKING order="12" place="12" resultid="2810" />
                    <RANKING order="13" place="13" resultid="2627" />
                    <RANKING order="14" place="14" resultid="4137" />
                    <RANKING order="15" place="15" resultid="2432" />
                    <RANKING order="16" place="16" resultid="3132" />
                    <RANKING order="17" place="17" resultid="3754" />
                    <RANKING order="18" place="18" resultid="2857" />
                    <RANKING order="19" place="19" resultid="2850" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6279" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4165" />
                    <RANKING order="2" place="2" resultid="3013" />
                    <RANKING order="3" place="-1" resultid="4272" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6280" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2453" />
                    <RANKING order="2" place="2" resultid="3605" />
                    <RANKING order="3" place="3" resultid="4603" />
                    <RANKING order="4" place="4" resultid="2918" />
                    <RANKING order="5" place="5" resultid="2547" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6281" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3496" />
                    <RANKING order="2" place="2" resultid="2604" />
                    <RANKING order="3" place="3" resultid="3510" />
                    <RANKING order="4" place="4" resultid="3859" />
                    <RANKING order="5" place="5" resultid="3871" />
                    <RANKING order="6" place="6" resultid="3363" />
                    <RANKING order="7" place="7" resultid="3091" />
                    <RANKING order="8" place="8" resultid="3119" />
                    <RANKING order="9" place="-1" resultid="4313" />
                    <RANKING order="10" place="-1" resultid="2553" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6282" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2404" />
                    <RANKING order="2" place="2" resultid="3307" />
                    <RANKING order="3" place="-1" resultid="3561" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6283" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2575" />
                    <RANKING order="2" place="2" resultid="3247" />
                    <RANKING order="3" place="3" resultid="4236" />
                    <RANKING order="4" place="-1" resultid="2815" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6284" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2890" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6285" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2404" />
                    <RANKING order="2" place="2" resultid="3496" />
                    <RANKING order="3" place="3" resultid="2604" />
                    <RANKING order="4" place="4" resultid="3510" />
                    <RANKING order="5" place="5" resultid="2453" />
                    <RANKING order="6" place="6" resultid="3859" />
                    <RANKING order="7" place="7" resultid="2575" />
                    <RANKING order="8" place="8" resultid="3605" />
                    <RANKING order="9" place="9" resultid="4603" />
                    <RANKING order="10" place="10" resultid="2890" />
                    <RANKING order="11" place="11" resultid="3307" />
                    <RANKING order="12" place="12" resultid="3871" />
                    <RANKING order="13" place="13" resultid="3247" />
                    <RANKING order="14" place="14" resultid="2918" />
                    <RANKING order="15" place="15" resultid="2547" />
                    <RANKING order="16" place="16" resultid="4165" />
                    <RANKING order="17" place="17" resultid="3363" />
                    <RANKING order="18" place="18" resultid="3738" />
                    <RANKING order="19" place="19" resultid="3091" />
                    <RANKING order="20" place="20" resultid="3419" />
                    <RANKING order="21" place="21" resultid="3349" />
                    <RANKING order="22" place="22" resultid="3787" />
                    <RANKING order="23" place="23" resultid="4386" />
                    <RANKING order="24" place="24" resultid="3865" />
                    <RANKING order="25" place="25" resultid="3370" />
                    <RANKING order="26" place="26" resultid="3806" />
                    <RANKING order="27" place="27" resultid="4236" />
                    <RANKING order="28" place="28" resultid="2559" />
                    <RANKING order="29" place="29" resultid="4537" />
                    <RANKING order="30" place="30" resultid="3013" />
                    <RANKING order="31" place="31" resultid="3405" />
                    <RANKING order="32" place="32" resultid="3119" />
                    <RANKING order="33" place="33" resultid="2810" />
                    <RANKING order="34" place="34" resultid="2627" />
                    <RANKING order="35" place="35" resultid="4137" />
                    <RANKING order="36" place="36" resultid="2432" />
                    <RANKING order="37" place="37" resultid="3132" />
                    <RANKING order="38" place="38" resultid="3754" />
                    <RANKING order="39" place="39" resultid="2857" />
                    <RANKING order="40" place="40" resultid="2850" />
                    <RANKING order="41" place="-1" resultid="3561" />
                    <RANKING order="42" place="-1" resultid="4313" />
                    <RANKING order="43" place="-1" resultid="2815" />
                    <RANKING order="44" place="-1" resultid="4272" />
                    <RANKING order="45" place="-1" resultid="2553" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5315" daytime="09:34" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5316" daytime="09:38" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5317" daytime="09:44" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5318" daytime="09:48" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5319" daytime="09:52" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5320" daytime="09:56" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1259" daytime="10:00" gender="F" number="37" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6286" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2661" />
                    <RANKING order="2" place="2" resultid="2515" />
                    <RANKING order="3" place="3" resultid="4049" />
                    <RANKING order="4" place="4" resultid="2511" />
                    <RANKING order="5" place="5" resultid="3425" />
                    <RANKING order="6" place="6" resultid="2635" />
                    <RANKING order="7" place="7" resultid="2741" />
                    <RANKING order="8" place="8" resultid="4116" />
                    <RANKING order="9" place="9" resultid="4072" />
                    <RANKING order="10" place="10" resultid="4516" />
                    <RANKING order="11" place="11" resultid="4180" />
                    <RANKING order="12" place="12" resultid="2766" />
                    <RANKING order="13" place="13" resultid="4629" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6287" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2426" />
                    <RANKING order="2" place="2" resultid="3701" />
                    <RANKING order="3" place="3" resultid="2649" />
                    <RANKING order="4" place="4" resultid="2829" />
                    <RANKING order="5" place="5" resultid="4549" />
                    <RANKING order="6" place="6" resultid="4361" />
                    <RANKING order="7" place="7" resultid="2729" />
                    <RANKING order="8" place="8" resultid="3532" />
                    <RANKING order="9" place="9" resultid="4643" />
                    <RANKING order="10" place="10" resultid="4354" />
                    <RANKING order="11" place="11" resultid="2508" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6288" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4423" />
                    <RANKING order="2" place="2" resultid="3477" />
                    <RANKING order="3" place="2" resultid="4159" />
                    <RANKING order="4" place="4" resultid="2950" />
                    <RANKING order="5" place="5" resultid="2599" />
                    <RANKING order="6" place="6" resultid="4472" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6289" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3472" />
                    <RANKING order="2" place="2" resultid="3321" />
                    <RANKING order="3" place="3" resultid="2588" />
                    <RANKING order="4" place="4" resultid="4376" />
                    <RANKING order="5" place="5" resultid="4363" />
                    <RANKING order="6" place="6" resultid="2993" />
                    <RANKING order="7" place="7" resultid="2616" />
                    <RANKING order="8" place="8" resultid="2736" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6290" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3252" />
                    <RANKING order="2" place="2" resultid="2973" />
                    <RANKING order="3" place="3" resultid="2966" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6291" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4438" />
                    <RANKING order="2" place="2" resultid="3955" />
                    <RANKING order="3" place="3" resultid="3044" />
                    <RANKING order="4" place="4" resultid="4309" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6292" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4496" />
                    <RANKING order="2" place="2" resultid="4289" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6293" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4423" />
                    <RANKING order="2" place="2" resultid="3472" />
                    <RANKING order="3" place="3" resultid="3321" />
                    <RANKING order="4" place="4" resultid="3477" />
                    <RANKING order="5" place="4" resultid="4159" />
                    <RANKING order="6" place="6" resultid="2588" />
                    <RANKING order="7" place="7" resultid="2426" />
                    <RANKING order="8" place="8" resultid="4438" />
                    <RANKING order="9" place="9" resultid="3701" />
                    <RANKING order="10" place="10" resultid="2661" />
                    <RANKING order="11" place="11" resultid="4496" />
                    <RANKING order="12" place="12" resultid="2515" />
                    <RANKING order="13" place="13" resultid="4376" />
                    <RANKING order="14" place="14" resultid="2649" />
                    <RANKING order="15" place="14" resultid="3252" />
                    <RANKING order="16" place="16" resultid="3955" />
                    <RANKING order="17" place="17" resultid="4049" />
                    <RANKING order="18" place="18" resultid="3044" />
                    <RANKING order="19" place="19" resultid="2950" />
                    <RANKING order="20" place="20" resultid="2829" />
                    <RANKING order="21" place="21" resultid="2599" />
                    <RANKING order="22" place="22" resultid="4549" />
                    <RANKING order="23" place="23" resultid="4361" />
                    <RANKING order="24" place="24" resultid="4472" />
                    <RANKING order="25" place="25" resultid="2511" />
                    <RANKING order="26" place="26" resultid="2729" />
                    <RANKING order="27" place="27" resultid="4363" />
                    <RANKING order="28" place="28" resultid="2993" />
                    <RANKING order="29" place="29" resultid="3532" />
                    <RANKING order="30" place="30" resultid="2616" />
                    <RANKING order="31" place="31" resultid="3425" />
                    <RANKING order="32" place="32" resultid="4643" />
                    <RANKING order="33" place="33" resultid="4309" />
                    <RANKING order="34" place="34" resultid="4289" />
                    <RANKING order="35" place="35" resultid="2635" />
                    <RANKING order="36" place="36" resultid="2741" />
                    <RANKING order="37" place="37" resultid="4116" />
                    <RANKING order="38" place="38" resultid="4072" />
                    <RANKING order="39" place="39" resultid="2736" />
                    <RANKING order="40" place="40" resultid="4516" />
                    <RANKING order="41" place="41" resultid="4180" />
                    <RANKING order="42" place="42" resultid="2973" />
                    <RANKING order="43" place="43" resultid="2766" />
                    <RANKING order="44" place="44" resultid="2966" />
                    <RANKING order="45" place="45" resultid="4629" />
                    <RANKING order="46" place="46" resultid="4354" />
                    <RANKING order="47" place="47" resultid="2508" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5321" daytime="10:00" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5322" daytime="10:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5323" daytime="10:04" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5324" daytime="10:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5325" daytime="10:08" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5326" daytime="10:10" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1267" daytime="10:12" gender="M" number="38" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6294" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2622" />
                    <RANKING order="2" place="2" resultid="4617" />
                    <RANKING order="3" place="3" resultid="3146" />
                    <RANKING order="4" place="4" resultid="3731" />
                    <RANKING order="5" place="5" resultid="3418" />
                    <RANKING order="6" place="6" resultid="3769" />
                    <RANKING order="7" place="7" resultid="2836" />
                    <RANKING order="8" place="8" resultid="4136" />
                    <RANKING order="9" place="9" resultid="3217" />
                    <RANKING order="10" place="10" resultid="2758" />
                    <RANKING order="11" place="11" resultid="2844" />
                    <RANKING order="12" place="12" resultid="2655" />
                    <RANKING order="13" place="13" resultid="2929" />
                    <RANKING order="14" place="14" resultid="2961" />
                    <RANKING order="15" place="15" resultid="4209" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6295" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2535" />
                    <RANKING order="2" place="2" resultid="4531" />
                    <RANKING order="3" place="3" resultid="3632" />
                    <RANKING order="4" place="4" resultid="3300" />
                    <RANKING order="5" place="5" resultid="4657" />
                    <RANKING order="6" place="6" resultid="3709" />
                    <RANKING order="7" place="7" resultid="3670" />
                    <RANKING order="8" place="8" resultid="2679" />
                    <RANKING order="9" place="9" resultid="4087" />
                    <RANKING order="10" place="10" resultid="2439" />
                    <RANKING order="11" place="11" resultid="4393" />
                    <RANKING order="12" place="12" resultid="3440" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6296" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2528" />
                    <RANKING order="2" place="2" resultid="2447" />
                    <RANKING order="3" place="3" resultid="3949" />
                    <RANKING order="4" place="4" resultid="4459" />
                    <RANKING order="5" place="5" resultid="2610" />
                    <RANKING order="6" place="6" resultid="2939" />
                    <RANKING order="7" place="7" resultid="2486" />
                    <RANKING order="8" place="8" resultid="3544" />
                    <RANKING order="9" place="9" resultid="3501" />
                    <RANKING order="10" place="10" resultid="4465" />
                    <RANKING order="11" place="11" resultid="3272" />
                    <RANKING order="12" place="12" resultid="2924" />
                    <RANKING order="13" place="13" resultid="2979" />
                    <RANKING order="14" place="14" resultid="3615" />
                    <RANKING order="15" place="-1" resultid="4636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6297" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3578" />
                    <RANKING order="2" place="2" resultid="3505" />
                    <RANKING order="3" place="3" resultid="3938" />
                    <RANKING order="4" place="4" resultid="3823" />
                    <RANKING order="5" place="5" resultid="3913" />
                    <RANKING order="6" place="6" resultid="4151" />
                    <RANKING order="7" place="7" resultid="3398" />
                    <RANKING order="8" place="7" resultid="4445" />
                    <RANKING order="9" place="9" resultid="4061" />
                    <RANKING order="10" place="10" resultid="4480" />
                    <RANKING order="11" place="11" resultid="2543" />
                    <RANKING order="12" place="12" resultid="2666" />
                    <RANKING order="13" place="13" resultid="3057" />
                    <RANKING order="14" place="14" resultid="2998" />
                    <RANKING order="15" place="15" resultid="2989" />
                    <RANKING order="16" place="16" resultid="4400" />
                    <RANKING order="17" place="-1" resultid="2873" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6298" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2403" />
                    <RANKING order="2" place="2" resultid="4431" />
                    <RANKING order="3" place="3" resultid="4252" />
                    <RANKING order="4" place="4" resultid="3097" />
                    <RANKING order="5" place="5" resultid="4296" />
                    <RANKING order="6" place="6" resultid="4190" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6299" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3483" />
                    <RANKING order="2" place="2" resultid="3986" />
                    <RANKING order="3" place="3" resultid="3719" />
                    <RANKING order="4" place="4" resultid="4504" />
                    <RANKING order="5" place="5" resultid="4326" />
                    <RANKING order="6" place="6" resultid="4556" />
                    <RANKING order="7" place="7" resultid="2494" />
                    <RANKING order="8" place="8" resultid="3246" />
                    <RANKING order="9" place="9" resultid="2582" />
                    <RANKING order="10" place="10" resultid="3185" />
                    <RANKING order="11" place="11" resultid="2901" />
                    <RANKING order="12" place="12" resultid="3195" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6300" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2566" />
                    <RANKING order="2" place="2" resultid="2788" />
                    <RANKING order="3" place="3" resultid="2783" />
                    <RANKING order="4" place="4" resultid="3895" />
                    <RANKING order="5" place="5" resultid="3063" />
                    <RANKING order="6" place="6" resultid="2912" />
                    <RANKING order="7" place="7" resultid="3077" />
                    <RANKING order="8" place="8" resultid="2896" />
                    <RANKING order="9" place="9" resultid="3226" />
                    <RANKING order="10" place="-1" resultid="2793" />
                    <RANKING order="11" place="-1" resultid="3050" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6301" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2566" />
                    <RANKING order="2" place="2" resultid="2788" />
                    <RANKING order="3" place="3" resultid="3483" />
                    <RANKING order="4" place="4" resultid="3986" />
                    <RANKING order="5" place="5" resultid="2403" />
                    <RANKING order="6" place="6" resultid="3719" />
                    <RANKING order="7" place="7" resultid="2528" />
                    <RANKING order="8" place="8" resultid="3578" />
                    <RANKING order="9" place="9" resultid="2783" />
                    <RANKING order="10" place="10" resultid="2535" />
                    <RANKING order="11" place="11" resultid="3895" />
                    <RANKING order="12" place="12" resultid="2447" />
                    <RANKING order="13" place="13" resultid="4431" />
                    <RANKING order="14" place="14" resultid="4504" />
                    <RANKING order="15" place="15" resultid="3505" />
                    <RANKING order="16" place="16" resultid="4326" />
                    <RANKING order="17" place="17" resultid="3949" />
                    <RANKING order="18" place="17" resultid="4556" />
                    <RANKING order="19" place="19" resultid="3063" />
                    <RANKING order="20" place="20" resultid="2494" />
                    <RANKING order="21" place="21" resultid="4252" />
                    <RANKING order="22" place="22" resultid="4459" />
                    <RANKING order="23" place="23" resultid="2912" />
                    <RANKING order="24" place="24" resultid="2610" />
                    <RANKING order="25" place="24" resultid="3938" />
                    <RANKING order="26" place="26" resultid="3823" />
                    <RANKING order="27" place="27" resultid="3913" />
                    <RANKING order="28" place="28" resultid="2939" />
                    <RANKING order="29" place="29" resultid="2486" />
                    <RANKING order="30" place="30" resultid="4151" />
                    <RANKING order="31" place="31" resultid="3398" />
                    <RANKING order="32" place="31" resultid="4445" />
                    <RANKING order="33" place="33" resultid="3246" />
                    <RANKING order="34" place="34" resultid="3544" />
                    <RANKING order="35" place="35" resultid="2582" />
                    <RANKING order="36" place="36" resultid="3501" />
                    <RANKING order="37" place="37" resultid="3077" />
                    <RANKING order="38" place="38" resultid="4465" />
                    <RANKING order="39" place="39" resultid="4061" />
                    <RANKING order="40" place="40" resultid="4480" />
                    <RANKING order="41" place="40" resultid="4531" />
                    <RANKING order="42" place="42" resultid="2896" />
                    <RANKING order="43" place="43" resultid="3272" />
                    <RANKING order="44" place="44" resultid="2543" />
                    <RANKING order="45" place="45" resultid="3185" />
                    <RANKING order="46" place="46" resultid="2901" />
                    <RANKING order="47" place="47" resultid="2622" />
                    <RANKING order="48" place="48" resultid="2666" />
                    <RANKING order="49" place="49" resultid="3057" />
                    <RANKING order="50" place="50" resultid="2924" />
                    <RANKING order="51" place="50" resultid="2998" />
                    <RANKING order="52" place="52" resultid="2989" />
                    <RANKING order="53" place="53" resultid="4617" />
                    <RANKING order="54" place="54" resultid="3195" />
                    <RANKING order="55" place="55" resultid="3146" />
                    <RANKING order="56" place="56" resultid="3632" />
                    <RANKING order="57" place="57" resultid="3097" />
                    <RANKING order="58" place="57" resultid="3731" />
                    <RANKING order="59" place="59" resultid="4400" />
                    <RANKING order="60" place="60" resultid="2979" />
                    <RANKING order="61" place="60" resultid="3300" />
                    <RANKING order="62" place="62" resultid="4657" />
                    <RANKING order="63" place="63" resultid="4296" />
                    <RANKING order="64" place="64" resultid="3226" />
                    <RANKING order="65" place="65" resultid="3615" />
                    <RANKING order="66" place="66" resultid="3709" />
                    <RANKING order="67" place="67" resultid="3670" />
                    <RANKING order="68" place="68" resultid="3418" />
                    <RANKING order="69" place="69" resultid="2679" />
                    <RANKING order="70" place="70" resultid="4087" />
                    <RANKING order="71" place="71" resultid="2439" />
                    <RANKING order="72" place="72" resultid="4393" />
                    <RANKING order="73" place="73" resultid="3440" />
                    <RANKING order="74" place="74" resultid="3769" />
                    <RANKING order="75" place="75" resultid="4190" />
                    <RANKING order="76" place="76" resultid="2836" />
                    <RANKING order="77" place="77" resultid="4136" />
                    <RANKING order="78" place="78" resultid="3217" />
                    <RANKING order="79" place="79" resultid="2758" />
                    <RANKING order="80" place="80" resultid="2844" />
                    <RANKING order="81" place="81" resultid="2655" />
                    <RANKING order="82" place="82" resultid="2929" />
                    <RANKING order="83" place="83" resultid="2961" />
                    <RANKING order="84" place="84" resultid="4209" />
                    <RANKING order="85" place="-1" resultid="2873" />
                    <RANKING order="86" place="-1" resultid="2793" />
                    <RANKING order="87" place="-1" resultid="3050" />
                    <RANKING order="88" place="-1" resultid="4636" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5327" daytime="10:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5328" daytime="10:16" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5329" daytime="10:18" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5330" daytime="10:20" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5331" daytime="10:22" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5332" daytime="10:24" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5333" daytime="10:26" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5334" daytime="10:28" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5335" daytime="10:30" number="9" order="9" status="OFFICIAL" />
                <HEAT heatid="5336" daytime="10:32" number="10" order="10" status="OFFICIAL" />
                <HEAT heatid="5337" daytime="10:32" number="11" order="11" status="OFFICIAL" />
                <HEAT heatid="5338" daytime="10:34" number="12" order="12" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1275" daytime="10:36" gender="F" number="39" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6302" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3800" />
                    <RANKING order="2" place="2" resultid="3844" />
                    <RANKING order="3" place="3" resultid="3927" />
                    <RANKING order="4" place="4" resultid="3782" />
                    <RANKING order="5" place="5" resultid="3413" />
                    <RANKING order="6" place="6" resultid="4247" />
                    <RANKING order="7" place="7" resultid="3003" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6303" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3280" />
                    <RANKING order="2" place="2" resultid="2419" />
                    <RANKING order="3" place="3" resultid="3650" />
                    <RANKING order="4" place="4" resultid="3657" />
                    <RANKING order="5" place="5" resultid="3644" />
                    <RANKING order="6" place="6" resultid="2641" />
                    <RANKING order="7" place="7" resultid="3975" />
                    <RANKING order="8" place="8" resultid="3688" />
                    <RANKING order="9" place="9" resultid="3160" />
                    <RANKING order="10" place="10" resultid="2830" />
                    <RANKING order="11" place="11" resultid="3434" />
                    <RANKING order="12" place="12" resultid="4650" />
                    <RANKING order="13" place="13" resultid="4355" />
                    <RANKING order="14" place="-1" resultid="4227" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6304" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2879" />
                    <RANKING order="2" place="2" resultid="3265" />
                    <RANKING order="3" place="3" resultid="3287" />
                    <RANKING order="4" place="4" resultid="4382" />
                    <RANKING order="5" place="5" resultid="3105" />
                    <RANKING order="6" place="6" resultid="2594" />
                    <RANKING order="7" place="7" resultid="4511" />
                    <RANKING order="8" place="-1" resultid="3612" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6305" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3944" />
                    <RANKING order="2" place="2" resultid="3041" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6306" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2974" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6307" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2778" />
                    <RANKING order="2" place="2" resultid="2570" />
                    <RANKING order="3" place="3" resultid="3045" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6308" agemax="-1" agemin="20" />
                <AGEGROUP agegroupid="6309" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3944" />
                    <RANKING order="2" place="2" resultid="2879" />
                    <RANKING order="3" place="3" resultid="3280" />
                    <RANKING order="4" place="4" resultid="2778" />
                    <RANKING order="5" place="5" resultid="3800" />
                    <RANKING order="6" place="6" resultid="2419" />
                    <RANKING order="7" place="7" resultid="3041" />
                    <RANKING order="8" place="8" resultid="3650" />
                    <RANKING order="9" place="9" resultid="3265" />
                    <RANKING order="10" place="10" resultid="3657" />
                    <RANKING order="11" place="11" resultid="3644" />
                    <RANKING order="12" place="12" resultid="3287" />
                    <RANKING order="13" place="13" resultid="3844" />
                    <RANKING order="14" place="14" resultid="3927" />
                    <RANKING order="15" place="15" resultid="3782" />
                    <RANKING order="16" place="16" resultid="2570" />
                    <RANKING order="17" place="17" resultid="2641" />
                    <RANKING order="18" place="18" resultid="3413" />
                    <RANKING order="19" place="19" resultid="4382" />
                    <RANKING order="20" place="20" resultid="3975" />
                    <RANKING order="21" place="21" resultid="3105" />
                    <RANKING order="22" place="22" resultid="3688" />
                    <RANKING order="23" place="23" resultid="3160" />
                    <RANKING order="24" place="24" resultid="3045" />
                    <RANKING order="25" place="25" resultid="2594" />
                    <RANKING order="26" place="26" resultid="2830" />
                    <RANKING order="27" place="27" resultid="3434" />
                    <RANKING order="28" place="28" resultid="4650" />
                    <RANKING order="29" place="29" resultid="4247" />
                    <RANKING order="30" place="30" resultid="4511" />
                    <RANKING order="31" place="31" resultid="3003" />
                    <RANKING order="32" place="32" resultid="4355" />
                    <RANKING order="33" place="33" resultid="2974" />
                    <RANKING order="34" place="-1" resultid="4227" />
                    <RANKING order="35" place="-1" resultid="3612" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5339" daytime="10:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5340" daytime="10:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5341" daytime="10:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5342" daytime="10:52" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5343" daytime="10:58" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1277" daytime="11:02" gender="M" number="40" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6310" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3314" />
                    <RANKING order="2" place="2" resultid="3831" />
                    <RANKING order="3" place="3" resultid="3328" />
                    <RANKING order="4" place="4" resultid="4130" />
                    <RANKING order="5" place="5" resultid="2748" />
                    <RANKING order="6" place="6" resultid="4524" />
                    <RANKING order="7" place="7" resultid="3794" />
                    <RANKING order="8" place="8" resultid="4202" />
                    <RANKING order="9" place="9" resultid="3406" />
                    <RANKING order="10" place="10" resultid="4145" />
                    <RANKING order="11" place="11" resultid="3866" />
                    <RANKING order="12" place="12" resultid="4103" />
                    <RANKING order="13" place="13" resultid="3878" />
                    <RANKING order="14" place="-1" resultid="3725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6311" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3294" />
                    <RANKING order="2" place="2" resultid="3392" />
                    <RANKING order="3" place="3" resultid="3153" />
                    <RANKING order="4" place="4" resultid="3682" />
                    <RANKING order="5" place="5" resultid="3168" />
                    <RANKING order="6" place="6" resultid="3638" />
                    <RANKING order="7" place="7" resultid="4612" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6312" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2884" />
                    <RANKING order="2" place="2" resultid="3980" />
                    <RANKING order="3" place="3" resultid="4604" />
                    <RANKING order="4" place="4" resultid="3356" />
                    <RANKING order="5" place="5" resultid="4259" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6313" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3490" />
                    <RANKING order="2" place="2" resultid="3261" />
                    <RANKING order="3" place="3" resultid="3626" />
                    <RANKING order="4" place="4" resultid="3573" />
                    <RANKING order="5" place="5" resultid="3567" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6314" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4370" />
                    <RANKING order="2" place="2" resultid="4065" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6315" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3484" />
                    <RANKING order="2" place="2" resultid="3070" />
                    <RANKING order="3" place="3" resultid="3084" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6316" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3813" />
                    <RANKING order="2" place="2" resultid="3064" />
                    <RANKING order="3" place="3" resultid="3240" />
                    <RANKING order="4" place="4" resultid="2891" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6317" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3813" />
                    <RANKING order="2" place="2" resultid="3484" />
                    <RANKING order="3" place="3" resultid="2884" />
                    <RANKING order="4" place="4" resultid="3490" />
                    <RANKING order="5" place="5" resultid="3980" />
                    <RANKING order="6" place="6" resultid="3261" />
                    <RANKING order="7" place="7" resultid="3626" />
                    <RANKING order="8" place="8" resultid="3064" />
                    <RANKING order="9" place="9" resultid="3294" />
                    <RANKING order="10" place="10" resultid="4604" />
                    <RANKING order="11" place="11" resultid="3573" />
                    <RANKING order="12" place="12" resultid="3356" />
                    <RANKING order="13" place="13" resultid="3070" />
                    <RANKING order="14" place="14" resultid="3240" />
                    <RANKING order="15" place="15" resultid="3314" />
                    <RANKING order="16" place="16" resultid="3831" />
                    <RANKING order="17" place="17" resultid="3392" />
                    <RANKING order="18" place="18" resultid="3084" />
                    <RANKING order="19" place="19" resultid="3153" />
                    <RANKING order="20" place="20" resultid="3567" />
                    <RANKING order="21" place="20" resultid="4259" />
                    <RANKING order="22" place="22" resultid="2891" />
                    <RANKING order="23" place="23" resultid="3682" />
                    <RANKING order="24" place="24" resultid="3168" />
                    <RANKING order="25" place="25" resultid="4370" />
                    <RANKING order="26" place="26" resultid="3638" />
                    <RANKING order="27" place="27" resultid="3328" />
                    <RANKING order="28" place="28" resultid="4130" />
                    <RANKING order="29" place="29" resultid="2748" />
                    <RANKING order="30" place="30" resultid="4524" />
                    <RANKING order="31" place="31" resultid="3794" />
                    <RANKING order="32" place="31" resultid="4612" />
                    <RANKING order="33" place="33" resultid="4202" />
                    <RANKING order="34" place="34" resultid="3406" />
                    <RANKING order="35" place="35" resultid="4145" />
                    <RANKING order="36" place="36" resultid="4065" />
                    <RANKING order="37" place="37" resultid="3866" />
                    <RANKING order="38" place="38" resultid="4103" />
                    <RANKING order="39" place="39" resultid="3878" />
                    <RANKING order="40" place="-1" resultid="3725" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5344" daytime="11:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5345" daytime="11:06" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5346" daytime="11:12" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5347" daytime="11:16" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5348" daytime="11:20" number="5" order="5" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1279" daytime="11:24" gender="F" number="41" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6318" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3342" />
                    <RANKING order="2" place="2" resultid="3775" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6319" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4321" />
                    <RANKING order="2" place="2" resultid="3140" />
                    <RANKING order="3" place="3" resultid="3689" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6320" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="3527" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6321" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2868" />
                    <RANKING order="2" place="2" resultid="2799" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6322" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3550" />
                    <RANKING order="2" place="2" resultid="3253" />
                    <RANKING order="3" place="3" resultid="4197" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6323" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="6324" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3908" />
                    <RANKING order="2" place="2" resultid="3919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6325" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3908" />
                    <RANKING order="2" place="2" resultid="3919" />
                    <RANKING order="3" place="3" resultid="3550" />
                    <RANKING order="4" place="4" resultid="3342" />
                    <RANKING order="5" place="5" resultid="4321" />
                    <RANKING order="6" place="6" resultid="3140" />
                    <RANKING order="7" place="7" resultid="3689" />
                    <RANKING order="8" place="8" resultid="3253" />
                    <RANKING order="9" place="9" resultid="2868" />
                    <RANKING order="10" place="10" resultid="3775" />
                    <RANKING order="11" place="11" resultid="4197" />
                    <RANKING order="12" place="12" resultid="2799" />
                    <RANKING order="13" place="-1" resultid="3527" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5349" daytime="11:24" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5350" daytime="11:48" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1281" daytime="12:10" gender="X" number="42" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1282" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4011" />
                    <RANKING order="2" place="2" resultid="4025" />
                    <RANKING order="3" place="3" resultid="3455" />
                    <RANKING order="4" place="4" resultid="2692" />
                    <RANKING order="5" place="5" resultid="4680" />
                    <RANKING order="6" place="6" resultid="3442" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5351" daytime="12:10" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1283" daytime="12:16" gender="X" number="43" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1284" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4010" />
                    <RANKING order="2" place="2" resultid="3454" />
                    <RANKING order="3" place="3" resultid="4679" />
                    <RANKING order="4" place="4" resultid="4024" />
                    <RANKING order="5" place="5" resultid="3176" />
                    <RANKING order="6" place="6" resultid="2691" />
                    <RANKING order="7" place="7" resultid="4682" />
                    <RANKING order="8" place="8" resultid="4416" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5352" daytime="12:16" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1285" daytime="12:24" gender="X" number="44" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1286" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3034" />
                    <RANKING order="2" place="2" resultid="4009" />
                    <RANKING order="3" place="3" resultid="4678" />
                    <RANKING order="4" place="4" resultid="4023" />
                    <RANKING order="5" place="5" resultid="4681" />
                    <RANKING order="6" place="6" resultid="3453" />
                    <RANKING order="7" place="7" resultid="2690" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5353" daytime="12:24" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1287" daytime="12:30" gender="X" number="45" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1288" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4006" />
                    <RANKING order="2" place="2" resultid="4022" />
                    <RANKING order="3" place="3" resultid="2689" />
                    <RANKING order="4" place="4" resultid="3175" />
                    <RANKING order="5" place="5" resultid="4414" />
                    <RANKING order="6" place="6" resultid="4677" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5354" daytime="12:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1289" daytime="12:36" gender="X" number="46" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1290" agemax="19" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4007" />
                    <RANKING order="2" place="2" resultid="4415" />
                    <RANKING order="3" place="3" resultid="3033" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5355" daytime="12:36" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1291" daytime="12:42" gender="X" number="47" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1292" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4008" />
                    <RANKING order="2" place="2" resultid="2522" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5356" daytime="12:42" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-09-21" daytime="16:10" endtime="19:30" number="6" officialmeeting="15:30" teamleadermeeting="16:00" warmupfrom="15:00" warmupuntil="16:00">
          <EVENTS>
            <EVENT eventid="2359" daytime="16:10" gender="M" number="16" order="1" round="FIN" preveventid="1182">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6368" agemax="-1" agemin="13" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6141" />
                    <RANKING order="2" place="2" resultid="6142" />
                    <RANKING order="3" place="3" resultid="6144" />
                    <RANKING order="4" place="4" resultid="6143" />
                    <RANKING order="5" place="5" resultid="6147" />
                    <RANKING order="6" place="6" resultid="6448" />
                    <RANKING order="7" place="7" resultid="6149" />
                    <RANKING order="8" place="8" resultid="6148" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6423" agegroupid="6368" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2391" daytime="16:12" gender="F" number="15" order="2" round="FIN" preveventid="1175">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6367" agemax="-1" agemin="13" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="6129" />
                    <RANKING order="2" place="2" resultid="6128" />
                    <RANKING order="3" place="3" resultid="6127" />
                    <RANKING order="4" place="4" resultid="6131" />
                    <RANKING order="5" place="5" resultid="6465" />
                    <RANKING order="6" place="6" resultid="6132" />
                    <RANKING order="7" place="7" resultid="6134" />
                    <RANKING order="8" place="8" resultid="6135" />
                    <RANKING order="9" place="8" resultid="6136" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6424" agegroupid="6367" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1293" daytime="16:16" gender="M" number="48" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6326" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3315" />
                    <RANKING order="2" place="2" resultid="3350" />
                    <RANKING order="3" place="3" resultid="3732" />
                    <RANKING order="4" place="4" resultid="4525" />
                    <RANKING order="5" place="5" resultid="4138" />
                    <RANKING order="6" place="-1" resultid="3147" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6327" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2934" />
                    <RANKING order="2" place="2" resultid="2536" />
                    <RANKING order="3" place="3" resultid="4532" />
                    <RANKING order="4" place="4" resultid="3301" />
                    <RANKING order="5" place="5" resultid="4598" />
                    <RANKING order="6" place="6" resultid="4394" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6328" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3273" />
                    <RANKING order="2" place="2" resultid="3357" />
                    <RANKING order="3" place="3" resultid="3950" />
                    <RANKING order="4" place="4" resultid="2529" />
                    <RANKING order="5" place="5" resultid="2611" />
                    <RANKING order="6" place="6" resultid="2925" />
                    <RANKING order="7" place="-1" resultid="2454" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6329" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3399" />
                    <RANKING order="2" place="2" resultid="3824" />
                    <RANKING order="3" place="-1" resultid="3579" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6330" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3522" />
                    <RANKING order="2" place="2" resultid="4253" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6331" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3071" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6332" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2913" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6333" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3522" />
                    <RANKING order="2" place="2" resultid="3399" />
                    <RANKING order="3" place="3" resultid="3273" />
                    <RANKING order="4" place="4" resultid="3357" />
                    <RANKING order="5" place="5" resultid="3071" />
                    <RANKING order="6" place="6" resultid="3950" />
                    <RANKING order="7" place="7" resultid="3824" />
                    <RANKING order="8" place="8" resultid="2934" />
                    <RANKING order="9" place="9" resultid="3315" />
                    <RANKING order="10" place="10" resultid="2529" />
                    <RANKING order="11" place="11" resultid="2913" />
                    <RANKING order="12" place="12" resultid="2611" />
                    <RANKING order="13" place="13" resultid="4253" />
                    <RANKING order="14" place="14" resultid="2536" />
                    <RANKING order="15" place="15" resultid="2925" />
                    <RANKING order="16" place="16" resultid="4532" />
                    <RANKING order="17" place="17" resultid="3350" />
                    <RANKING order="18" place="18" resultid="3301" />
                    <RANKING order="19" place="19" resultid="3732" />
                    <RANKING order="20" place="20" resultid="4525" />
                    <RANKING order="21" place="21" resultid="4598" />
                    <RANKING order="22" place="22" resultid="4138" />
                    <RANKING order="23" place="23" resultid="4394" />
                    <RANKING order="24" place="-1" resultid="2454" />
                    <RANKING order="25" place="-1" resultid="3147" />
                    <RANKING order="26" place="-1" resultid="3579" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5357" daytime="16:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5358" daytime="16:20" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5359" daytime="16:24" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5360" daytime="16:28" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1295" daytime="16:32" gender="F" number="49" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6334" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3855" />
                    <RANKING order="2" place="2" resultid="3336" />
                    <RANKING order="3" place="3" resultid="3343" />
                    <RANKING order="4" place="4" resultid="3427" />
                    <RANKING order="5" place="5" resultid="3378" />
                    <RANKING order="6" place="6" resultid="2742" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6335" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3702" />
                    <RANKING order="2" place="2" resultid="4550" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6336" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6337" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="6338" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3254" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6339" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="6340" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3920" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6341" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4424" />
                    <RANKING order="2" place="2" resultid="3855" />
                    <RANKING order="3" place="3" resultid="3920" />
                    <RANKING order="4" place="4" resultid="3336" />
                    <RANKING order="5" place="5" resultid="3702" />
                    <RANKING order="6" place="6" resultid="4550" />
                    <RANKING order="7" place="7" resultid="3254" />
                    <RANKING order="8" place="8" resultid="3343" />
                    <RANKING order="9" place="9" resultid="3427" />
                    <RANKING order="10" place="10" resultid="3378" />
                    <RANKING order="11" place="11" resultid="2742" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5361" daytime="16:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5362" daytime="16:38" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1297" daytime="16:42" gender="M" number="50" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6342" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2628" />
                    <RANKING order="2" place="2" resultid="3788" />
                    <RANKING order="3" place="3" resultid="2504" />
                    <RANKING order="4" place="4" resultid="3329" />
                    <RANKING order="5" place="5" resultid="3739" />
                    <RANKING order="6" place="6" resultid="4387" />
                    <RANKING order="7" place="7" resultid="3420" />
                    <RANKING order="8" place="8" resultid="4538" />
                    <RANKING order="9" place="9" resultid="2560" />
                    <RANKING order="10" place="10" resultid="4543" />
                    <RANKING order="11" place="11" resultid="2433" />
                    <RANKING order="12" place="12" resultid="2811" />
                    <RANKING order="13" place="13" resultid="2837" />
                    <RANKING order="14" place="14" resultid="3755" />
                    <RANKING order="15" place="15" resultid="4203" />
                    <RANKING order="16" place="16" resultid="2858" />
                    <RANKING order="17" place="17" resultid="4110" />
                    <RANKING order="18" place="18" resultid="2759" />
                    <RANKING order="19" place="19" resultid="3133" />
                    <RANKING order="20" place="20" resultid="2851" />
                    <RANKING order="21" place="21" resultid="4210" />
                    <RANKING order="22" place="-1" resultid="3371" />
                    <RANKING order="23" place="-1" resultid="4622" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6343" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4166" />
                    <RANKING order="2" place="2" resultid="3014" />
                    <RANKING order="3" place="3" resultid="3441" />
                    <RANKING order="4" place="4" resultid="4662" />
                    <RANKING order="5" place="5" resultid="3695" />
                    <RANKING order="6" place="6" resultid="2984" />
                    <RANKING order="7" place="7" resultid="2680" />
                    <RANKING order="8" place="8" resultid="2440" />
                    <RANKING order="9" place="9" resultid="3154" />
                    <RANKING order="10" place="-1" resultid="3024" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6344" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4303" />
                    <RANKING order="2" place="2" resultid="4605" />
                    <RANKING order="3" place="3" resultid="2940" />
                    <RANKING order="4" place="4" resultid="3606" />
                    <RANKING order="5" place="5" resultid="2548" />
                    <RANKING order="6" place="6" resultid="4494" />
                    <RANKING order="7" place="7" resultid="2919" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6345" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3511" />
                    <RANKING order="2" place="2" resultid="2605" />
                    <RANKING order="3" place="3" resultid="3939" />
                    <RANKING order="4" place="4" resultid="3860" />
                    <RANKING order="5" place="5" resultid="2804" />
                    <RANKING order="6" place="6" resultid="3872" />
                    <RANKING order="7" place="7" resultid="4401" />
                    <RANKING order="8" place="8" resultid="2554" />
                    <RANKING order="9" place="9" resultid="4152" />
                    <RANKING order="10" place="10" resultid="2667" />
                    <RANKING order="11" place="11" resultid="4314" />
                    <RANKING order="12" place="12" resultid="3364" />
                    <RANKING order="13" place="13" resultid="4083" />
                    <RANKING order="14" place="-1" resultid="4278" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6346" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2405" />
                    <RANKING order="2" place="2" resultid="3562" />
                    <RANKING order="3" place="3" resultid="3308" />
                    <RANKING order="4" place="4" resultid="4405" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6347" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2888" />
                    <RANKING order="2" place="2" resultid="2576" />
                    <RANKING order="3" place="3" resultid="2816" />
                    <RANKING order="4" place="4" resultid="4557" />
                    <RANKING order="5" place="5" resultid="2495" />
                    <RANKING order="6" place="6" resultid="2583" />
                    <RANKING order="7" place="7" resultid="4237" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6348" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2457" />
                    <RANKING order="2" place="2" resultid="2567" />
                    <RANKING order="3" place="3" resultid="2908" />
                    <RANKING order="4" place="4" resultid="3078" />
                    <RANKING order="5" place="-1" resultid="3227" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6349" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2457" />
                    <RANKING order="2" place="2" resultid="2567" />
                    <RANKING order="3" place="3" resultid="2405" />
                    <RANKING order="4" place="4" resultid="2888" />
                    <RANKING order="5" place="5" resultid="3511" />
                    <RANKING order="6" place="6" resultid="2605" />
                    <RANKING order="7" place="7" resultid="3939" />
                    <RANKING order="8" place="8" resultid="2576" />
                    <RANKING order="9" place="9" resultid="3562" />
                    <RANKING order="10" place="10" resultid="3860" />
                    <RANKING order="11" place="11" resultid="4303" />
                    <RANKING order="12" place="12" resultid="2816" />
                    <RANKING order="13" place="13" resultid="4605" />
                    <RANKING order="14" place="14" resultid="4557" />
                    <RANKING order="15" place="15" resultid="2940" />
                    <RANKING order="16" place="16" resultid="2495" />
                    <RANKING order="17" place="17" resultid="2908" />
                    <RANKING order="18" place="18" resultid="3606" />
                    <RANKING order="19" place="19" resultid="2548" />
                    <RANKING order="20" place="20" resultid="2804" />
                    <RANKING order="21" place="20" resultid="4494" />
                    <RANKING order="22" place="22" resultid="4166" />
                    <RANKING order="23" place="23" resultid="3872" />
                    <RANKING order="24" place="24" resultid="2919" />
                    <RANKING order="25" place="25" resultid="4401" />
                    <RANKING order="26" place="26" resultid="3308" />
                    <RANKING order="27" place="27" resultid="2554" />
                    <RANKING order="28" place="28" resultid="2583" />
                    <RANKING order="29" place="29" resultid="2628" />
                    <RANKING order="30" place="30" resultid="3788" />
                    <RANKING order="31" place="31" resultid="4152" />
                    <RANKING order="32" place="32" resultid="4237" />
                    <RANKING order="33" place="33" resultid="2667" />
                    <RANKING order="34" place="34" resultid="4314" />
                    <RANKING order="35" place="35" resultid="2504" />
                    <RANKING order="36" place="36" resultid="3329" />
                    <RANKING order="37" place="37" resultid="3739" />
                    <RANKING order="38" place="38" resultid="3078" />
                    <RANKING order="39" place="39" resultid="4405" />
                    <RANKING order="40" place="40" resultid="3364" />
                    <RANKING order="41" place="41" resultid="4387" />
                    <RANKING order="42" place="42" resultid="4083" />
                    <RANKING order="43" place="43" resultid="3014" />
                    <RANKING order="44" place="44" resultid="3420" />
                    <RANKING order="45" place="45" resultid="3441" />
                    <RANKING order="46" place="46" resultid="4662" />
                    <RANKING order="47" place="47" resultid="4538" />
                    <RANKING order="48" place="48" resultid="2560" />
                    <RANKING order="49" place="49" resultid="4543" />
                    <RANKING order="50" place="50" resultid="3695" />
                    <RANKING order="51" place="51" resultid="2433" />
                    <RANKING order="52" place="52" resultid="2984" />
                    <RANKING order="53" place="53" resultid="2811" />
                    <RANKING order="54" place="54" resultid="2680" />
                    <RANKING order="55" place="55" resultid="2440" />
                    <RANKING order="56" place="56" resultid="3154" />
                    <RANKING order="57" place="57" resultid="2837" />
                    <RANKING order="58" place="58" resultid="3755" />
                    <RANKING order="59" place="59" resultid="4203" />
                    <RANKING order="60" place="60" resultid="2858" />
                    <RANKING order="61" place="61" resultid="4110" />
                    <RANKING order="62" place="62" resultid="2759" />
                    <RANKING order="63" place="63" resultid="3133" />
                    <RANKING order="64" place="64" resultid="2851" />
                    <RANKING order="65" place="65" resultid="4210" />
                    <RANKING order="66" place="-1" resultid="3371" />
                    <RANKING order="67" place="-1" resultid="3024" />
                    <RANKING order="68" place="-1" resultid="3227" />
                    <RANKING order="69" place="-1" resultid="4622" />
                    <RANKING order="70" place="-1" resultid="4278" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5363" daytime="16:42" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5364" daytime="16:44" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5365" daytime="16:48" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5366" daytime="16:50" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5367" daytime="16:52" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5368" daytime="16:54" number="6" order="6" status="OFFICIAL" />
                <HEAT heatid="5369" daytime="16:56" number="7" order="7" status="OFFICIAL" />
                <HEAT heatid="5370" daytime="16:58" number="8" order="8" status="OFFICIAL" />
                <HEAT heatid="5371" daytime="17:00" number="9" order="9" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1305" daytime="17:02" gender="F" number="51" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6350" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3749" />
                    <RANKING order="2" place="2" resultid="3933" />
                    <RANKING order="3" place="3" resultid="4571" />
                    <RANKING order="4" place="4" resultid="3776" />
                    <RANKING order="5" place="5" resultid="3762" />
                    <RANKING order="6" place="6" resultid="2673" />
                    <RANKING order="7" place="7" resultid="4518" />
                    <RANKING order="8" place="8" resultid="2723" />
                    <RANKING order="9" place="9" resultid="3126" />
                    <RANKING order="10" place="-1" resultid="3200" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6351" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4266" />
                    <RANKING order="2" place="2" resultid="4584" />
                    <RANKING order="3" place="3" resultid="2642" />
                    <RANKING order="4" place="4" resultid="4215" />
                    <RANKING order="5" place="5" resultid="3161" />
                    <RANKING order="6" place="6" resultid="2509" />
                    <RANKING order="7" place="7" resultid="2705" />
                    <RANKING order="8" place="-1" resultid="3889" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6352" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2945" />
                    <RANKING order="2" place="2" resultid="3601" />
                    <RANKING order="3" place="3" resultid="3596" />
                    <RANKING order="4" place="4" resultid="3538" />
                    <RANKING order="5" place="5" resultid="2481" />
                    <RANKING order="6" place="6" resultid="2823" />
                    <RANKING order="7" place="7" resultid="3266" />
                    <RANKING order="8" place="8" resultid="3189" />
                    <RANKING order="9" place="9" resultid="4487" />
                    <RANKING order="10" place="-1" resultid="4473" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6353" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2589" />
                    <RANKING order="2" place="2" resultid="3322" />
                    <RANKING order="3" place="3" resultid="4377" />
                    <RANKING order="4" place="4" resultid="3848" />
                    <RANKING order="5" place="5" resultid="2717" />
                    <RANKING order="6" place="6" resultid="4452" />
                    <RANKING order="7" place="7" resultid="2412" />
                    <RANKING order="8" place="8" resultid="3042" />
                    <RANKING order="9" place="9" resultid="4667" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6354" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="6355" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3957" />
                    <RANKING order="2" place="2" resultid="2462" />
                    <RANKING order="3" place="3" resultid="4241" />
                    <RANKING order="4" place="4" resultid="2571" />
                    <RANKING order="5" place="5" resultid="3046" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6356" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4030" />
                    <RANKING order="2" place="-1" resultid="4497" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6357" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3957" />
                    <RANKING order="2" place="2" resultid="4030" />
                    <RANKING order="3" place="3" resultid="4266" />
                    <RANKING order="4" place="4" resultid="2589" />
                    <RANKING order="5" place="5" resultid="2945" />
                    <RANKING order="6" place="6" resultid="3322" />
                    <RANKING order="7" place="7" resultid="4584" />
                    <RANKING order="8" place="8" resultid="3601" />
                    <RANKING order="9" place="9" resultid="4377" />
                    <RANKING order="10" place="10" resultid="3848" />
                    <RANKING order="11" place="11" resultid="3596" />
                    <RANKING order="12" place="12" resultid="3538" />
                    <RANKING order="13" place="13" resultid="3749" />
                    <RANKING order="14" place="14" resultid="2462" />
                    <RANKING order="15" place="15" resultid="3933" />
                    <RANKING order="16" place="16" resultid="2717" />
                    <RANKING order="17" place="17" resultid="2481" />
                    <RANKING order="18" place="18" resultid="2823" />
                    <RANKING order="19" place="19" resultid="4571" />
                    <RANKING order="20" place="20" resultid="2642" />
                    <RANKING order="21" place="21" resultid="3776" />
                    <RANKING order="22" place="22" resultid="3762" />
                    <RANKING order="23" place="23" resultid="3266" />
                    <RANKING order="24" place="24" resultid="4452" />
                    <RANKING order="25" place="25" resultid="3189" />
                    <RANKING order="26" place="26" resultid="4215" />
                    <RANKING order="27" place="27" resultid="2412" />
                    <RANKING order="28" place="28" resultid="3042" />
                    <RANKING order="29" place="29" resultid="4487" />
                    <RANKING order="30" place="30" resultid="4241" />
                    <RANKING order="31" place="31" resultid="2673" />
                    <RANKING order="32" place="32" resultid="2571" />
                    <RANKING order="33" place="33" resultid="3161" />
                    <RANKING order="34" place="34" resultid="4518" />
                    <RANKING order="35" place="35" resultid="2509" />
                    <RANKING order="36" place="36" resultid="4667" />
                    <RANKING order="37" place="37" resultid="2723" />
                    <RANKING order="38" place="38" resultid="3126" />
                    <RANKING order="39" place="39" resultid="3046" />
                    <RANKING order="40" place="40" resultid="2705" />
                    <RANKING order="41" place="-1" resultid="3200" />
                    <RANKING order="42" place="-1" resultid="4473" />
                    <RANKING order="43" place="-1" resultid="4497" />
                    <RANKING order="44" place="-1" resultid="3889" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5372" daytime="17:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5373" daytime="17:04" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5374" daytime="17:06" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="5375" daytime="17:08" number="4" order="4" status="OFFICIAL" />
                <HEAT heatid="5376" daytime="17:10" number="5" order="5" status="OFFICIAL" />
                <HEAT heatid="5377" daytime="17:12" number="6" order="6" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2383" daytime="17:14" gender="M" number="6" order="7" round="FIN" preveventid="1104">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6375" agemax="-1" agemin="13" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5981" />
                    <RANKING order="2" place="2" resultid="5979" />
                    <RANKING order="3" place="3" resultid="5980" />
                    <RANKING order="4" place="4" resultid="5982" />
                    <RANKING order="5" place="5" resultid="5984" />
                    <RANKING order="6" place="6" resultid="5983" />
                    <RANKING order="7" place="7" resultid="5986" />
                    <RANKING order="8" place="8" resultid="5985" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="6425" agegroupid="6375" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="2375" daytime="17:16" gender="F" number="5" order="8" round="FIN" preveventid="1096">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="5399" agemax="-1" agemin="13" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="5968" />
                    <RANKING order="2" place="2" resultid="5969" />
                    <RANKING order="3" place="3" resultid="5970" />
                    <RANKING order="4" place="4" resultid="5974" />
                    <RANKING order="5" place="5" resultid="5971" />
                    <RANKING order="6" place="6" resultid="5973" />
                    <RANKING order="7" place="7" resultid="5977" />
                    <RANKING order="8" place="8" resultid="5976" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5978" agegroupid="5399" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1312" daytime="17:18" gender="M" number="52" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="1500" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="3100" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="6358" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3726" />
                    <RANKING order="2" place="2" resultid="4348" />
                    <RANKING order="3" place="3" resultid="3207" />
                    <RANKING order="4" place="4" resultid="4577" />
                    <RANKING order="5" place="5" resultid="3879" />
                    <RANKING order="6" place="6" resultid="4131" />
                    <RANKING order="7" place="7" resultid="3224" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6359" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3683" />
                    <RANKING order="2" place="2" resultid="4597" />
                    <RANKING order="3" place="3" resultid="4273" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6360" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4260" />
                    <RANKING order="2" place="2" resultid="4466" />
                    <RANKING order="3" place="3" resultid="3621" />
                    <RANKING order="4" place="4" resultid="4124" />
                    <RANKING order="5" place="-1" resultid="2492" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6361" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3092" />
                    <RANKING order="2" place="2" resultid="3112" />
                    <RANKING order="3" place="3" resultid="3183" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6362" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3098" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6363" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3085" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6364" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2905" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="6365" agemax="-1" agemin="-1" name="Troféu Paraná (Infantil/Sênior) 2024">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4260" />
                    <RANKING order="2" place="2" resultid="4466" />
                    <RANKING order="3" place="3" resultid="3621" />
                    <RANKING order="4" place="4" resultid="3092" />
                    <RANKING order="5" place="5" resultid="3683" />
                    <RANKING order="6" place="6" resultid="3085" />
                    <RANKING order="7" place="7" resultid="4124" />
                    <RANKING order="8" place="8" resultid="4597" />
                    <RANKING order="9" place="9" resultid="3112" />
                    <RANKING order="10" place="10" resultid="3726" />
                    <RANKING order="11" place="11" resultid="4348" />
                    <RANKING order="12" place="12" resultid="4273" />
                    <RANKING order="13" place="13" resultid="2905" />
                    <RANKING order="14" place="14" resultid="3098" />
                    <RANKING order="15" place="15" resultid="3207" />
                    <RANKING order="16" place="16" resultid="4577" />
                    <RANKING order="17" place="17" resultid="3879" />
                    <RANKING order="18" place="18" resultid="4131" />
                    <RANKING order="19" place="19" resultid="3224" />
                    <RANKING order="20" place="20" resultid="3183" />
                    <RANKING order="21" place="-1" resultid="2492" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5378" daytime="17:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="5379" daytime="17:42" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="5380" daytime="18:08" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1320" daytime="18:28" gender="F" number="53" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1321" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3994" />
                    <RANKING order="2" place="2" resultid="4015" />
                    <RANKING order="3" place="3" resultid="3446" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5381" daytime="18:28" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1322" daytime="18:36" gender="F" number="54" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1323" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3993" />
                    <RANKING order="2" place="2" resultid="3445" />
                    <RANKING order="3" place="3" resultid="2684" />
                    <RANKING order="4" place="4" resultid="4014" />
                    <RANKING order="5" place="5" resultid="4670" />
                    <RANKING order="6" place="6" resultid="4407" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5382" daytime="18:36" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1324" daytime="18:44" gender="F" number="55" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1325" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3992" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5383" daytime="18:44" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1326" daytime="18:50" gender="F" number="56" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1327" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="3026" />
                    <RANKING order="2" place="2" resultid="2683" />
                    <RANKING order="3" place="-1" resultid="3991" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5384" daytime="18:50" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1328" daytime="18:56" gender="F" number="57" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1329" agemax="19" agemin="17" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1330" daytime="18:56" gender="F" number="58" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1331" agemax="-1" agemin="20" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1332" daytime="18:56" gender="M" number="59" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1333" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4002" />
                    <RANKING order="2" place="2" resultid="4674" />
                    <RANKING order="3" place="3" resultid="4020" />
                    <RANKING order="4" place="4" resultid="2862" />
                    <RANKING order="5" place="-1" resultid="3450" />
                    <RANKING order="6" place="-1" resultid="2687" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5385" daytime="18:56" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1334" daytime="19:02" gender="M" number="60" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1335" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4003" />
                    <RANKING order="2" place="2" resultid="4021" />
                    <RANKING order="3" place="3" resultid="3031" />
                    <RANKING order="4" place="4" resultid="4675" />
                    <RANKING order="5" place="5" resultid="3173" />
                    <RANKING order="6" place="6" resultid="4412" />
                    <RANKING order="7" place="-1" resultid="3451" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5386" daytime="19:02" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1336" daytime="19:10" gender="M" number="61" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1337" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4005" />
                    <RANKING order="2" place="2" resultid="3032" />
                    <RANKING order="3" place="-1" resultid="4676" />
                    <RANKING order="4" place="-1" resultid="2521" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5387" daytime="19:10" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1338" daytime="19:16" gender="M" number="62" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1339" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4004" />
                    <RANKING order="2" place="2" resultid="3452" />
                    <RANKING order="3" place="3" resultid="2688" />
                    <RANKING order="4" place="4" resultid="4413" />
                    <RANKING order="5" place="5" resultid="3174" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5388" daytime="19:16" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1340" daytime="19:22" gender="M" number="63" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1341" agemax="19" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="4001" />
                    <RANKING order="2" place="2" resultid="4411" />
                    <RANKING order="3" place="-1" resultid="4019" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5389" daytime="19:22" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1342" daytime="19:28" gender="M" number="64" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="4" stroke="MEDLEY" />
              <FEE currency="BRL" value="12400" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1343" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="2861" />
                    <RANKING order="2" place="2" resultid="3172" />
                    <RANKING order="3" place="3" resultid="3030" />
                    <RANKING order="4" place="-1" resultid="4000" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="5390" daytime="19:28" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="1007" nation="BRA" region="PR" clubid="4417" swrid="93785" name="Santa Mônica Clube De Campo" shortname="Santa Mônica">
          <ATHLETES>
            <ATHLETE firstname="Henrique" lastname="Blansky Hagebock" birthdate="2008-08-15" gender="M" nation="BRA" license="339123" swrid="5455418" athleteid="4474" externalid="339123">
              <RESULTS>
                <RESULT eventid="1072" points="442" swimtime="00:04:48.87" resultid="4475" heatid="5061" lane="3" entrytime="00:04:42.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="100" swimtime="00:01:07.09" />
                    <SPLIT distance="150" swimtime="00:01:43.76" />
                    <SPLIT distance="200" swimtime="00:02:21.36" />
                    <SPLIT distance="250" swimtime="00:02:58.40" />
                    <SPLIT distance="300" swimtime="00:03:35.84" />
                    <SPLIT distance="350" swimtime="00:04:13.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="513" swimtime="00:00:26.11" resultid="4476" heatid="5125" lane="4" entrytime="00:00:25.73" entrycourse="LCM" />
                <RESULT eventid="1120" points="454" swimtime="00:02:12.70" resultid="4477" heatid="5155" lane="5" entrytime="00:02:09.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                    <SPLIT distance="100" swimtime="00:01:04.59" />
                    <SPLIT distance="150" swimtime="00:01:39.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="578" swimtime="00:00:56.23" resultid="4478" heatid="5229" lane="5" entrytime="00:00:57.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="366" swimtime="00:00:32.91" resultid="4479" heatid="5285" lane="2" entrytime="00:00:34.22" entrycourse="LCM" />
                <RESULT eventid="1267" points="447" swimtime="00:00:29.11" resultid="4480" heatid="5335" lane="8" entrytime="00:00:28.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Giuseppe Bulla Lanaro" birthdate="2007-05-22" gender="M" nation="BRA" license="331630" swrid="5600174" athleteid="4425" externalid="331630">
              <RESULTS>
                <RESULT eventid="1072" points="578" swimtime="00:04:24.07" resultid="4426" heatid="5064" lane="5" entrytime="00:04:12.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.45" />
                    <SPLIT distance="100" swimtime="00:01:00.82" />
                    <SPLIT distance="150" swimtime="00:01:33.98" />
                    <SPLIT distance="200" swimtime="00:02:07.80" />
                    <SPLIT distance="250" swimtime="00:02:42.53" />
                    <SPLIT distance="300" swimtime="00:03:17.22" />
                    <SPLIT distance="350" swimtime="00:03:52.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="567" swimtime="00:00:25.25" resultid="4427" heatid="5129" lane="6" entrytime="00:00:25.08" entrycourse="LCM" />
                <RESULT eventid="1120" points="620" swimtime="00:01:59.58" resultid="4428" heatid="5158" lane="6" entrytime="00:01:57.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.65" />
                    <SPLIT distance="100" swimtime="00:00:57.83" />
                    <SPLIT distance="150" swimtime="00:01:28.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="530" swimtime="00:02:20.85" resultid="4429" heatid="5199" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="150" swimtime="00:01:50.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="663" swimtime="00:00:53.74" resultid="4430" heatid="5233" lane="1" entrytime="00:00:53.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="540" swimtime="00:00:27.34" resultid="4431" heatid="5336" lane="8" entrytime="00:00:27.81" entrycourse="LCM" />
                <RESULT eventid="2351" points="650" swimtime="00:00:54.08" resultid="6122" heatid="6422" lane="1" entrytime="00:00:53.74">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Marcos Morais" birthdate="2010-01-30" gender="M" nation="BRA" license="416736" athleteid="4658" externalid="416736">
              <RESULTS>
                <RESULT eventid="1088" points="273" swimtime="00:01:27.64" resultid="4659" heatid="5078" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="275" swimtime="00:02:36.73" resultid="4660" heatid="5148" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:01:14.00" />
                    <SPLIT distance="150" swimtime="00:01:56.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="324" swimtime="00:01:08.18" resultid="4661" heatid="5218" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="299" swimtime="00:00:38.78" resultid="4662" heatid="5364" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="F" nation="BRA" license="344301" swrid="5569976" athleteid="4418" externalid="344301">
              <RESULTS>
                <RESULT eventid="1064" points="607" swimtime="00:04:37.93" resultid="4419" heatid="5053" lane="5" entrytime="00:04:41.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                    <SPLIT distance="100" swimtime="00:01:08.04" />
                    <SPLIT distance="150" swimtime="00:01:44.00" />
                    <SPLIT distance="200" swimtime="00:02:19.74" />
                    <SPLIT distance="250" swimtime="00:02:54.98" />
                    <SPLIT distance="300" swimtime="00:03:30.29" />
                    <SPLIT distance="350" swimtime="00:04:04.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="595" swimtime="00:00:28.06" resultid="4420" heatid="5104" lane="3" entrytime="00:00:28.49" entrycourse="LCM" />
                <RESULT eventid="1128" points="608" swimtime="00:01:05.47" resultid="4421" heatid="5161" lane="4" entrytime="00:01:04.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="634" swimtime="00:01:00.19" resultid="4422" heatid="5208" lane="5" entrytime="00:01:00.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="546" swimtime="00:00:29.88" resultid="4423" heatid="5326" lane="4" entrytime="00:00:29.79" entrycourse="LCM" />
                <RESULT eventid="1295" points="526" swimtime="00:02:30.87" resultid="4424" heatid="5362" lane="5" entrytime="00:02:27.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                    <SPLIT distance="100" swimtime="00:01:12.48" />
                    <SPLIT distance="150" swimtime="00:01:53.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2375" points="570" swimtime="00:00:28.46" resultid="5970" heatid="5978" lane="3" entrytime="00:00:28.06" />
                <RESULT eventid="2328" points="610" swimtime="00:01:05.40" resultid="5998" heatid="6418" lane="5" entrytime="00:01:05.47">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2343" points="622" swimtime="00:01:00.55" resultid="6102" heatid="6421" lane="5" entrytime="00:01:00.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.84" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emily" lastname="Sayuri Tangueria De Lima" birthdate="2010-06-11" gender="F" nation="BRA" license="367215" swrid="5588901" athleteid="4544" externalid="367215">
              <RESULTS>
                <RESULT eventid="1064" points="449" swimtime="00:05:07.21" resultid="4545" heatid="5051" lane="8" entrytime="00:05:05.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:12.93" />
                    <SPLIT distance="150" swimtime="00:01:52.38" />
                    <SPLIT distance="200" swimtime="00:02:32.41" />
                    <SPLIT distance="250" swimtime="00:03:11.86" />
                    <SPLIT distance="300" swimtime="00:03:51.73" />
                    <SPLIT distance="350" swimtime="00:04:31.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="413" swimtime="00:00:31.68" resultid="4546" heatid="5098" lane="3" entrytime="00:00:32.31" entrycourse="LCM" />
                <RESULT eventid="1128" points="382" swimtime="00:01:16.41" resultid="4547" heatid="5160" lane="6" entrytime="00:01:15.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="426" swimtime="00:01:08.68" resultid="4548" heatid="5203" lane="1" entrytime="00:01:10.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="356" swimtime="00:00:34.46" resultid="4549" heatid="5326" lane="7" entrytime="00:00:32.97" entrycourse="LCM" />
                <RESULT eventid="1295" points="331" swimtime="00:02:55.98" resultid="4550" heatid="5362" lane="7" entrytime="00:02:53.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.32" />
                    <SPLIT distance="100" swimtime="00:01:21.46" />
                    <SPLIT distance="150" swimtime="00:02:10.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Schlickmann Assis" birthdate="2003-07-24" gender="F" nation="BRA" license="303874" swrid="5600257" athleteid="4495" externalid="303874">
              <RESULTS>
                <RESULT eventid="1259" points="403" swimtime="00:00:33.05" resultid="4496" heatid="5322" lane="8" />
                <RESULT eventid="1305" status="DNS" swimtime="00:00:00.00" resultid="4497" heatid="5377" lane="2" entrytime="00:00:36.93" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Inoue Kuroda" birthdate="2009-04-18" gender="M" nation="BRA" license="324700" swrid="5600190" athleteid="4460" externalid="324700">
              <RESULTS>
                <RESULT eventid="1104" points="485" swimtime="00:00:26.61" resultid="4461" heatid="5124" lane="3" entrytime="00:00:26.81" entrycourse="LCM" />
                <RESULT eventid="1120" points="485" swimtime="00:02:09.76" resultid="4462" heatid="5156" lane="7" entrytime="00:02:06.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.65" />
                    <SPLIT distance="100" swimtime="00:01:02.81" />
                    <SPLIT distance="150" swimtime="00:01:36.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="540" swimtime="00:00:57.53" resultid="4463" heatid="5230" lane="1" entrytime="00:00:56.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="446" swimtime="00:00:30.82" resultid="4464" heatid="5282" lane="8" />
                <RESULT eventid="1267" points="450" swimtime="00:00:29.04" resultid="4465" heatid="5330" lane="6" />
                <RESULT eventid="1312" points="539" swimtime="00:17:49.98" resultid="4466" heatid="5380" lane="5" entrytime="00:17:30.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.00" />
                    <SPLIT distance="100" swimtime="00:01:05.07" />
                    <SPLIT distance="150" swimtime="00:01:40.11" />
                    <SPLIT distance="200" swimtime="00:02:15.61" />
                    <SPLIT distance="250" swimtime="00:02:51.71" />
                    <SPLIT distance="300" swimtime="00:03:27.29" />
                    <SPLIT distance="350" swimtime="00:04:02.73" />
                    <SPLIT distance="400" swimtime="00:04:38.32" />
                    <SPLIT distance="450" swimtime="00:05:14.00" />
                    <SPLIT distance="500" swimtime="00:05:49.50" />
                    <SPLIT distance="550" swimtime="00:06:24.98" />
                    <SPLIT distance="600" swimtime="00:07:01.14" />
                    <SPLIT distance="650" swimtime="00:07:37.17" />
                    <SPLIT distance="700" swimtime="00:08:13.19" />
                    <SPLIT distance="750" swimtime="00:08:50.27" />
                    <SPLIT distance="800" swimtime="00:09:26.63" />
                    <SPLIT distance="850" swimtime="00:10:03.47" />
                    <SPLIT distance="900" swimtime="00:10:40.16" />
                    <SPLIT distance="950" swimtime="00:11:16.30" />
                    <SPLIT distance="1000" swimtime="00:11:52.71" />
                    <SPLIT distance="1050" swimtime="00:12:29.26" />
                    <SPLIT distance="1100" swimtime="00:13:05.91" />
                    <SPLIT distance="1150" swimtime="00:13:42.88" />
                    <SPLIT distance="1200" swimtime="00:14:19.26" />
                    <SPLIT distance="1250" swimtime="00:14:55.52" />
                    <SPLIT distance="1300" swimtime="00:15:31.14" />
                    <SPLIT distance="1350" swimtime="00:16:07.35" />
                    <SPLIT distance="1400" swimtime="00:16:42.82" />
                    <SPLIT distance="1450" swimtime="00:17:18.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Araujo Felix" birthdate="2010-05-27" gender="F" nation="BRA" license="393157" swrid="5622260" athleteid="4637" externalid="393157">
              <RESULTS>
                <RESULT eventid="1096" points="413" swimtime="00:00:31.68" resultid="4638" heatid="5098" lane="4" entrytime="00:00:31.83" entrycourse="LCM" />
                <RESULT eventid="1128" points="219" swimtime="00:01:32.03" resultid="4639" heatid="5159" lane="5" entrytime="00:01:31.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="418" swimtime="00:02:30.86" resultid="4640" heatid="5139" lane="3" entrytime="00:02:32.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="100" swimtime="00:01:13.21" />
                    <SPLIT distance="150" swimtime="00:01:51.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="416" swimtime="00:01:09.23" resultid="4641" heatid="5203" lane="3" entrytime="00:01:09.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="352" swimtime="00:00:38.04" resultid="4642" heatid="5291" lane="5" entrytime="00:00:44.08" entrycourse="LCM" />
                <RESULT eventid="1259" points="283" swimtime="00:00:37.19" resultid="4643" heatid="5324" lane="8" entrytime="00:00:37.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Helena Vieira Jussen" birthdate="2011-12-29" gender="F" nation="BRA" license="372282" swrid="5588740" athleteid="4565" externalid="372282">
              <RESULTS>
                <RESULT eventid="1080" points="366" swimtime="00:01:29.63" resultid="4566" heatid="5066" lane="2" entrytime="00:01:31.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="290" swimtime="00:03:10.33" resultid="4567" heatid="5186" lane="3" entrytime="00:03:31.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.53" />
                    <SPLIT distance="100" swimtime="00:01:33.06" />
                    <SPLIT distance="150" swimtime="00:02:25.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="267" swimtime="00:01:28.98" resultid="4568" heatid="5242" lane="2" entrytime="00:01:27.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="258" swimtime="00:00:42.18" resultid="4569" heatid="5291" lane="4" entrytime="00:00:44.03" entrycourse="LCM" />
                <RESULT eventid="1243" points="345" swimtime="00:03:16.01" resultid="4570" heatid="5311" lane="3" entrytime="00:03:18.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.40" />
                    <SPLIT distance="100" swimtime="00:01:36.64" />
                    <SPLIT distance="150" swimtime="00:02:26.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="368" swimtime="00:00:40.68" resultid="4571" heatid="5375" lane="8" entrytime="00:00:43.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Larissa" lastname="Garcia Reschetti Rubbo" birthdate="2011-08-06" gender="F" nation="BRA" license="367053" swrid="5588720" athleteid="4512" externalid="367053" level="DCOMP IT">
              <RESULTS>
                <RESULT eventid="1080" points="337" swimtime="00:01:32.09" resultid="4513" heatid="5066" lane="7" entrytime="00:01:31.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="334" swimtime="00:00:34.00" resultid="4514" heatid="5098" lane="1" entrytime="00:00:33.09" entrycourse="LCM" />
                <RESULT eventid="1159" points="307" swimtime="00:01:16.60" resultid="4515" heatid="5202" lane="3" entrytime="00:01:14.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="184" swimtime="00:00:42.92" resultid="4516" heatid="5323" lane="3" entrytime="00:00:41.52" entrycourse="LCM" />
                <RESULT eventid="1243" points="324" swimtime="00:03:20.19" resultid="4517" heatid="5312" lane="8" entrytime="00:03:15.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.95" />
                    <SPLIT distance="100" swimtime="00:01:36.04" />
                    <SPLIT distance="150" swimtime="00:02:29.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="309" swimtime="00:00:43.09" resultid="4518" heatid="5374" lane="6" entrytime="00:00:44.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Vianna" birthdate="2011-01-31" gender="M" nation="BRA" license="371380" swrid="5588947" athleteid="4558" externalid="371380">
              <RESULTS>
                <RESULT eventid="1072" points="389" swimtime="00:05:01.32" resultid="4559" heatid="5058" lane="6" entrytime="00:05:00.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:11.99" />
                    <SPLIT distance="150" swimtime="00:01:51.35" />
                    <SPLIT distance="200" swimtime="00:02:30.72" />
                    <SPLIT distance="250" swimtime="00:03:09.15" />
                    <SPLIT distance="300" swimtime="00:03:48.91" />
                    <SPLIT distance="350" swimtime="00:04:25.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="334" swimtime="00:00:30.12" resultid="4560" heatid="5118" lane="7" entrytime="00:00:29.69" entrycourse="LCM" />
                <RESULT eventid="1135" points="326" swimtime="00:01:11.79" resultid="4561" heatid="5171" lane="6" entrytime="00:01:10.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 18:47), Na volta dos 150m (Medley Individual, Peito)." eventid="1151" status="DSQ" swimtime="00:02:51.42" resultid="4562" heatid="5193" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                    <SPLIT distance="100" swimtime="00:01:18.45" />
                    <SPLIT distance="150" swimtime="00:02:16.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="381" swimtime="00:01:04.61" resultid="4563" heatid="5221" lane="4" entrytime="00:01:04.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="359" swimtime="00:10:35.87" resultid="4564" heatid="5298" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="100" swimtime="00:01:15.42" />
                    <SPLIT distance="150" swimtime="00:01:55.90" />
                    <SPLIT distance="200" swimtime="00:02:36.59" />
                    <SPLIT distance="250" swimtime="00:03:16.81" />
                    <SPLIT distance="300" swimtime="00:03:56.60" />
                    <SPLIT distance="350" swimtime="00:04:36.84" />
                    <SPLIT distance="400" swimtime="00:05:17.61" />
                    <SPLIT distance="450" swimtime="00:05:58.44" />
                    <SPLIT distance="500" swimtime="00:06:38.71" />
                    <SPLIT distance="550" swimtime="00:07:19.94" />
                    <SPLIT distance="600" swimtime="00:08:01.15" />
                    <SPLIT distance="650" swimtime="00:08:41.74" />
                    <SPLIT distance="700" swimtime="00:09:21.69" />
                    <SPLIT distance="750" swimtime="00:10:01.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Marques Machado" birthdate="2010-02-17" gender="M" nation="BRA" license="390918" swrid="5600212" athleteid="4592" externalid="390918">
              <RESULTS>
                <RESULT eventid="1072" points="396" swimtime="00:04:59.53" resultid="4593" heatid="5056" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:08.74" />
                    <SPLIT distance="150" swimtime="00:01:47.51" />
                    <SPLIT distance="200" swimtime="00:02:25.42" />
                    <SPLIT distance="250" swimtime="00:03:03.72" />
                    <SPLIT distance="300" swimtime="00:03:42.47" />
                    <SPLIT distance="350" swimtime="00:04:21.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="265" swimtime="00:01:16.96" resultid="4594" heatid="5171" lane="1" entrytime="00:01:12.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="370" swimtime="00:02:22.06" resultid="4595" heatid="5151" lane="2" entrytime="00:02:19.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.51" />
                    <SPLIT distance="100" swimtime="00:01:09.04" />
                    <SPLIT distance="150" swimtime="00:01:45.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="362" swimtime="00:10:33.93" resultid="4596" heatid="5298" lane="3" entrytime="00:10:36.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                    <SPLIT distance="100" swimtime="00:01:09.91" />
                    <SPLIT distance="150" swimtime="00:01:48.10" />
                    <SPLIT distance="200" swimtime="00:02:27.56" />
                    <SPLIT distance="250" swimtime="00:03:07.53" />
                    <SPLIT distance="300" swimtime="00:03:48.64" />
                    <SPLIT distance="350" swimtime="00:04:30.20" />
                    <SPLIT distance="400" swimtime="00:05:10.97" />
                    <SPLIT distance="450" swimtime="00:05:52.70" />
                    <SPLIT distance="500" swimtime="00:06:34.31" />
                    <SPLIT distance="550" swimtime="00:07:15.77" />
                    <SPLIT distance="600" swimtime="00:07:57.12" />
                    <SPLIT distance="650" swimtime="00:08:38.14" />
                    <SPLIT distance="700" swimtime="00:09:18.97" />
                    <SPLIT distance="750" swimtime="00:09:57.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="410" swimtime="00:19:32.36" resultid="4597" heatid="5379" lane="2" entrytime="00:20:18.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:11.50" />
                    <SPLIT distance="150" swimtime="00:01:49.58" />
                    <SPLIT distance="200" swimtime="00:02:29.32" />
                    <SPLIT distance="250" swimtime="00:03:07.16" />
                    <SPLIT distance="300" swimtime="00:03:46.65" />
                    <SPLIT distance="350" swimtime="00:04:25.61" />
                    <SPLIT distance="400" swimtime="00:05:06.02" />
                    <SPLIT distance="450" swimtime="00:05:43.84" />
                    <SPLIT distance="500" swimtime="00:06:23.66" />
                    <SPLIT distance="550" swimtime="00:07:03.07" />
                    <SPLIT distance="600" swimtime="00:07:42.95" />
                    <SPLIT distance="650" swimtime="00:08:22.70" />
                    <SPLIT distance="700" swimtime="00:09:02.83" />
                    <SPLIT distance="750" swimtime="00:09:41.62" />
                    <SPLIT distance="800" swimtime="00:10:22.49" />
                    <SPLIT distance="850" swimtime="00:11:01.29" />
                    <SPLIT distance="900" swimtime="00:11:40.47" />
                    <SPLIT distance="950" swimtime="00:12:19.78" />
                    <SPLIT distance="1000" swimtime="00:13:00.12" />
                    <SPLIT distance="1050" swimtime="00:13:39.38" />
                    <SPLIT distance="1100" swimtime="00:14:19.03" />
                    <SPLIT distance="1150" swimtime="00:14:59.77" />
                    <SPLIT distance="1200" swimtime="00:15:39.69" />
                    <SPLIT distance="1250" swimtime="00:16:19.12" />
                    <SPLIT distance="1300" swimtime="00:16:58.76" />
                    <SPLIT distance="1350" swimtime="00:17:38.58" />
                    <SPLIT distance="1400" swimtime="00:18:18.36" />
                    <SPLIT distance="1450" swimtime="00:18:56.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1293" points="269" swimtime="00:02:50.77" resultid="4598" heatid="5358" lane="6" entrytime="00:02:49.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.69" />
                    <SPLIT distance="100" swimtime="00:01:21.92" />
                    <SPLIT distance="150" swimtime="00:02:08.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabio" lastname="C Burak" birthdate="2009-08-29" gender="M" nation="BRA" license="343297" swrid="5600126" athleteid="4599" externalid="343297">
              <RESULTS>
                <RESULT eventid="1088" points="479" swimtime="00:01:12.69" resultid="4600" heatid="5085" lane="1" entrytime="00:01:11.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="502" swimtime="00:02:23.44" resultid="4601" heatid="5198" lane="2" entrytime="00:02:21.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                    <SPLIT distance="100" swimtime="00:01:07.65" />
                    <SPLIT distance="150" swimtime="00:01:49.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="465" swimtime="00:01:06.56" resultid="4602" heatid="5260" lane="4" entrytime="00:01:06.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="467" swimtime="00:02:41.66" resultid="4603" heatid="5320" lane="8" entrytime="00:02:39.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:17.31" />
                    <SPLIT distance="150" swimtime="00:01:59.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="472" swimtime="00:02:23.73" resultid="4604" heatid="5346" lane="5" entrytime="00:02:30.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                    <SPLIT distance="100" swimtime="00:01:09.98" />
                    <SPLIT distance="150" swimtime="00:01:47.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="491" swimtime="00:00:32.89" resultid="4605" heatid="5369" lane="6" entrytime="00:00:34.98" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Dallastra" birthdate="2010-08-21" gender="M" nation="BRA" license="408024" swrid="5723028" athleteid="4651" externalid="408024">
              <RESULTS>
                <RESULT eventid="1072" points="423" swimtime="00:04:52.98" resultid="4652" heatid="5056" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="100" swimtime="00:01:08.15" />
                    <SPLIT distance="150" swimtime="00:01:45.24" />
                    <SPLIT distance="200" swimtime="00:02:23.68" />
                    <SPLIT distance="250" swimtime="00:03:02.47" />
                    <SPLIT distance="300" swimtime="00:03:40.68" />
                    <SPLIT distance="350" swimtime="00:04:17.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="384" swimtime="00:00:28.76" resultid="4653" heatid="5118" lane="5" entrytime="00:00:28.80" entrycourse="LCM" />
                <RESULT eventid="1135" points="249" swimtime="00:01:18.52" resultid="4654" heatid="5170" lane="6" entrytime="00:01:18.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="414" swimtime="00:02:16.76" resultid="4655" heatid="5151" lane="5" entrytime="00:02:17.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                    <SPLIT distance="100" swimtime="00:01:05.00" />
                    <SPLIT distance="150" swimtime="00:01:41.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="436" swimtime="00:01:01.77" resultid="4656" heatid="5222" lane="7" entrytime="00:01:02.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="335" swimtime="00:00:32.04" resultid="4657" heatid="5331" lane="6" entrytime="00:00:35.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Augusto Vaz" birthdate="2011-06-25" gender="M" nation="BRA" license="401737" swrid="5661339" athleteid="4613" externalid="401737">
              <RESULTS>
                <RESULT eventid="1104" points="366" swimtime="00:00:29.23" resultid="4614" heatid="5118" lane="1" entrytime="00:00:29.83" entrycourse="LCM" />
                <RESULT eventid="1120" points="347" swimtime="00:02:25.03" resultid="4615" heatid="5149" lane="8" entrytime="00:02:46.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.94" />
                    <SPLIT distance="100" swimtime="00:01:09.39" />
                    <SPLIT distance="150" swimtime="00:01:48.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="391" swimtime="00:01:04.03" resultid="4616" heatid="5221" lane="7" entrytime="00:01:05.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="373" swimtime="00:00:30.92" resultid="4617" heatid="5333" lane="8" entrytime="00:00:31.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Novakoski" birthdate="2009-03-05" gender="F" nation="BRA" license="339136" swrid="5600225" athleteid="4467" externalid="339136">
              <RESULTS>
                <RESULT eventid="1096" points="474" swimtime="00:00:30.28" resultid="4468" heatid="5103" lane="2" entrytime="00:00:30.14" entrycourse="LCM" />
                <RESULT eventid="1112" points="448" swimtime="00:02:27.48" resultid="4469" heatid="5143" lane="5" entrytime="00:02:27.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:11.36" />
                    <SPLIT distance="150" swimtime="00:01:50.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="504" swimtime="00:01:04.97" resultid="4470" heatid="5208" lane="8" entrytime="00:01:05.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="345" swimtime="00:11:30.61" resultid="4471" heatid="5272" lane="7" entrytime="00:11:16.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.11" />
                    <SPLIT distance="100" swimtime="00:01:15.75" />
                    <SPLIT distance="150" swimtime="00:01:57.82" />
                    <SPLIT distance="200" swimtime="00:02:40.84" />
                    <SPLIT distance="250" swimtime="00:03:23.81" />
                    <SPLIT distance="300" swimtime="00:04:07.59" />
                    <SPLIT distance="350" swimtime="00:04:50.96" />
                    <SPLIT distance="400" swimtime="00:05:35.58" />
                    <SPLIT distance="450" swimtime="00:06:19.67" />
                    <SPLIT distance="500" swimtime="00:07:04.30" />
                    <SPLIT distance="550" swimtime="00:07:48.93" />
                    <SPLIT distance="600" swimtime="00:08:34.24" />
                    <SPLIT distance="650" swimtime="00:09:19.74" />
                    <SPLIT distance="700" swimtime="00:10:05.76" />
                    <SPLIT distance="750" swimtime="00:10:50.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="351" swimtime="00:00:34.63" resultid="4472" heatid="5325" lane="3" entrytime="00:00:34.67" entrycourse="LCM" />
                <RESULT eventid="1305" status="DNS" swimtime="00:00:00.00" resultid="4473" heatid="5374" lane="3" entrytime="00:00:44.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Cavassin Ieger" birthdate="2011-08-31" gender="M" nation="BRA" license="367149" swrid="5588743" athleteid="4533" externalid="367149">
              <RESULTS>
                <RESULT eventid="1088" points="265" swimtime="00:01:28.55" resultid="4534" heatid="5080" lane="5" entrytime="00:01:30.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="314" swimtime="00:05:23.52" resultid="4535" heatid="5057" lane="1" entrytime="00:05:50.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:13.64" />
                    <SPLIT distance="150" swimtime="00:01:54.64" />
                    <SPLIT distance="200" swimtime="00:02:35.55" />
                    <SPLIT distance="250" swimtime="00:03:17.58" />
                    <SPLIT distance="300" swimtime="00:03:58.60" />
                    <SPLIT distance="350" swimtime="00:04:41.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="282" swimtime="00:02:53.83" resultid="4536" heatid="5193" lane="4" entrytime="00:02:54.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:01:24.84" />
                    <SPLIT distance="150" swimtime="00:02:13.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="287" swimtime="00:03:10.11" resultid="4537" heatid="5316" lane="4" entrytime="00:03:15.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.63" />
                    <SPLIT distance="100" swimtime="00:01:30.56" />
                    <SPLIT distance="150" swimtime="00:02:21.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="296" swimtime="00:00:38.92" resultid="4538" heatid="5366" lane="4" entrytime="00:00:41.26" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucca" lastname="Maceno Araujo" birthdate="2010-09-29" gender="M" nation="BRA" license="367056" swrid="5588788" athleteid="4526" externalid="367056">
              <RESULTS>
                <RESULT eventid="1072" points="422" swimtime="00:04:53.26" resultid="4527" heatid="5056" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                    <SPLIT distance="100" swimtime="00:01:06.60" />
                    <SPLIT distance="150" swimtime="00:01:44.79" />
                    <SPLIT distance="200" swimtime="00:02:22.54" />
                    <SPLIT distance="250" swimtime="00:03:01.39" />
                    <SPLIT distance="300" swimtime="00:03:39.89" />
                    <SPLIT distance="350" swimtime="00:04:18.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="390" swimtime="00:00:28.61" resultid="4528" heatid="5119" lane="1" entrytime="00:00:28.63" entrycourse="LCM" />
                <RESULT eventid="1135" points="402" swimtime="00:01:06.99" resultid="4529" heatid="5171" lane="5" entrytime="00:01:06.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="445" swimtime="00:01:01.36" resultid="4530" heatid="5222" lane="6" entrytime="00:01:01.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="447" swimtime="00:00:29.11" resultid="4531" heatid="5334" lane="3" entrytime="00:00:29.18" entrycourse="LCM" />
                <RESULT eventid="1293" points="341" swimtime="00:02:37.85" resultid="4532" heatid="5358" lane="5" entrytime="00:02:44.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:01:15.73" />
                    <SPLIT distance="150" swimtime="00:01:59.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Ieger" birthdate="2009-02-20" gender="M" nation="BRA" license="356888" swrid="5600180" athleteid="4488" externalid="356888">
              <RESULTS>
                <RESULT eventid="1088" points="398" swimtime="00:01:17.31" resultid="4489" heatid="5084" lane="8" entrytime="00:01:19.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="442" swimtime="00:00:27.44" resultid="4490" heatid="5124" lane="1" entrytime="00:00:27.18" entrycourse="LCM" />
                <RESULT eventid="1120" points="437" swimtime="00:02:14.36" resultid="4491" heatid="5154" lane="5" entrytime="00:02:17.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.67" />
                    <SPLIT distance="100" swimtime="00:01:03.27" />
                    <SPLIT distance="150" swimtime="00:01:39.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="484" swimtime="00:00:59.65" resultid="4492" heatid="5228" lane="8" entrytime="00:00:59.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="356" swimtime="00:00:33.22" resultid="4493" heatid="5282" lane="2" />
                <RESULT eventid="1297" points="439" swimtime="00:00:34.12" resultid="4494" heatid="5369" lane="5" entrytime="00:00:34.68" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Gelenski Pelaio" birthdate="2005-10-10" gender="M" nation="BRA" license="281473" swrid="5600173" athleteid="4551" externalid="281473" level="UNIDOMBOSC">
              <RESULTS>
                <RESULT eventid="1072" points="476" swimtime="00:04:41.83" resultid="4552" heatid="5063" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                    <SPLIT distance="100" swimtime="00:01:03.35" />
                    <SPLIT distance="150" swimtime="00:01:38.40" />
                    <SPLIT distance="200" swimtime="00:02:14.21" />
                    <SPLIT distance="250" swimtime="00:02:50.44" />
                    <SPLIT distance="300" swimtime="00:03:27.51" />
                    <SPLIT distance="350" swimtime="00:04:05.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="541" swimtime="00:00:25.66" resultid="4553" heatid="5129" lane="3" entrytime="00:00:24.92" entrycourse="LCM" />
                <RESULT eventid="1135" points="516" swimtime="00:01:01.62" resultid="4554" heatid="5177" lane="5" entrytime="00:01:00.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="537" swimtime="00:00:57.65" resultid="4555" heatid="5232" lane="2" entrytime="00:00:56.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="529" swimtime="00:00:27.52" resultid="4556" heatid="5338" lane="8" entrytime="00:00:26.80" entrycourse="LCM" />
                <RESULT eventid="1297" points="479" swimtime="00:00:33.16" resultid="4557" heatid="5370" lane="7" entrytime="00:00:33.59" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juliana" lastname="Moreira Furtado" birthdate="2011-01-27" gender="F" nation="BRA" license="403783" swrid="5684587" athleteid="4623" externalid="403783">
              <RESULTS>
                <RESULT eventid="1064" points="290" swimtime="00:05:55.21" resultid="4624" heatid="5048" lane="4" entrytime="00:05:59.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                    <SPLIT distance="100" swimtime="00:01:19.94" />
                    <SPLIT distance="150" swimtime="00:02:04.16" />
                    <SPLIT distance="200" swimtime="00:02:50.61" />
                    <SPLIT distance="250" swimtime="00:03:38.11" />
                    <SPLIT distance="300" swimtime="00:04:24.71" />
                    <SPLIT distance="350" swimtime="00:05:11.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="297" swimtime="00:00:35.38" resultid="4625" heatid="5097" lane="8" entrytime="00:00:36.10" entrycourse="LCM" />
                <RESULT eventid="1112" points="288" swimtime="00:02:50.70" resultid="4626" heatid="5138" lane="2" entrytime="00:02:49.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.27" />
                    <SPLIT distance="100" swimtime="00:01:22.34" />
                    <SPLIT distance="150" swimtime="00:02:07.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="207" swimtime="00:01:36.80" resultid="4627" heatid="5241" lane="3" entrytime="00:01:37.77" entrycourse="LCM" />
                <RESULT eventid="1159" points="303" swimtime="00:01:16.91" resultid="4628" heatid="5202" lane="1" entrytime="00:01:18.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="139" swimtime="00:00:47.14" resultid="4629" heatid="5322" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Analyce" lastname="Nunes Porto Luz" birthdate="2006-10-29" gender="F" nation="BRA" license="369322" swrid="5600226" athleteid="4432" externalid="369322">
              <RESULTS>
                <RESULT eventid="1064" points="466" swimtime="00:05:03.54" resultid="4433" heatid="5055" lane="2" entrytime="00:04:50.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                    <SPLIT distance="100" swimtime="00:01:10.72" />
                    <SPLIT distance="150" swimtime="00:01:49.04" />
                    <SPLIT distance="200" swimtime="00:02:27.86" />
                    <SPLIT distance="250" swimtime="00:03:06.55" />
                    <SPLIT distance="300" swimtime="00:03:46.06" />
                    <SPLIT distance="350" swimtime="00:04:25.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="508" swimtime="00:00:29.58" resultid="4434" heatid="5106" lane="6" entrytime="00:00:29.48" entrycourse="LCM" />
                <RESULT eventid="1128" points="464" swimtime="00:01:11.64" resultid="4435" heatid="5162" lane="4" entrytime="00:01:11.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="542" swimtime="00:01:03.42" resultid="4436" heatid="5209" lane="6" entrytime="00:01:03.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="432" swimtime="00:10:40.87" resultid="4437" heatid="5273" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.09" />
                    <SPLIT distance="100" swimtime="00:01:14.41" />
                    <SPLIT distance="150" swimtime="00:01:54.83" />
                    <SPLIT distance="200" swimtime="00:02:35.75" />
                    <SPLIT distance="250" swimtime="00:03:16.90" />
                    <SPLIT distance="300" swimtime="00:03:58.37" />
                    <SPLIT distance="350" swimtime="00:04:39.83" />
                    <SPLIT distance="400" swimtime="00:05:20.83" />
                    <SPLIT distance="450" swimtime="00:06:01.54" />
                    <SPLIT distance="500" swimtime="00:06:42.36" />
                    <SPLIT distance="550" swimtime="00:07:22.98" />
                    <SPLIT distance="600" swimtime="00:08:03.52" />
                    <SPLIT distance="650" swimtime="00:08:43.78" />
                    <SPLIT distance="700" swimtime="00:09:24.21" />
                    <SPLIT distance="750" swimtime="00:10:03.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="445" swimtime="00:00:31.99" resultid="4438" heatid="5326" lane="6" entrytime="00:00:31.37" entrycourse="LCM" />
                <RESULT eventid="2328" points="460" swimtime="00:01:11.83" resultid="5999" heatid="6418" lane="3" entrytime="00:01:11.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2343" points="547" swimtime="00:01:03.21" resultid="6108" heatid="6421" lane="8" entrytime="00:01:03.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="De Castro Paiva Maciel" birthdate="2008-04-10" gender="M" nation="BRA" license="378333" swrid="5622275" athleteid="4439" externalid="378333">
              <RESULTS>
                <RESULT eventid="1072" points="445" swimtime="00:04:48.10" resultid="4440" heatid="5061" lane="1" entrytime="00:05:26.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="100" swimtime="00:01:07.41" />
                    <SPLIT distance="150" swimtime="00:01:44.07" />
                    <SPLIT distance="200" swimtime="00:02:21.45" />
                    <SPLIT distance="250" swimtime="00:02:58.74" />
                    <SPLIT distance="300" swimtime="00:03:36.43" />
                    <SPLIT distance="350" swimtime="00:04:13.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="455" swimtime="00:00:27.18" resultid="4441" heatid="5124" lane="6" entrytime="00:00:26.88" entrycourse="LCM" />
                <RESULT eventid="1135" points="405" swimtime="00:01:06.83" resultid="4442" heatid="5174" lane="7" entrytime="00:01:05.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="504" swimtime="00:00:58.86" resultid="4443" heatid="5228" lane="2" entrytime="00:00:58.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="410" swimtime="00:00:31.70" resultid="4444" heatid="5281" lane="5" />
                <RESULT eventid="1267" points="485" swimtime="00:00:28.33" resultid="4445" heatid="5335" lane="1" entrytime="00:00:28.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diego" lastname="Brasil Caropreso" birthdate="2009-10-29" gender="M" nation="BRA" license="399502" swrid="5653287" athleteid="4630" externalid="399502">
              <RESULTS>
                <RESULT eventid="1072" points="331" swimtime="00:05:18.04" resultid="4631" heatid="5060" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:09.10" />
                    <SPLIT distance="150" swimtime="00:01:49.55" />
                    <SPLIT distance="200" swimtime="00:02:30.86" />
                    <SPLIT distance="250" swimtime="00:03:13.30" />
                    <SPLIT distance="300" swimtime="00:03:55.45" />
                    <SPLIT distance="350" swimtime="00:04:37.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="387" swimtime="00:00:28.68" resultid="4632" heatid="5123" lane="7" entrytime="00:00:28.15" entrycourse="LCM" />
                <RESULT eventid="1135" points="222" swimtime="00:01:21.64" resultid="4633" heatid="5173" lane="7" entrytime="00:01:17.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="395" swimtime="00:02:18.92" resultid="4634" heatid="5153" lane="4" entrytime="00:02:23.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.15" />
                    <SPLIT distance="100" swimtime="00:01:06.19" />
                    <SPLIT distance="150" swimtime="00:01:42.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="444" swimtime="00:01:01.41" resultid="4635" heatid="5226" lane="3" entrytime="00:01:02.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" status="DNS" swimtime="00:00:00.00" resultid="4636" heatid="5333" lane="1" entrytime="00:00:31.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Lopes Rempel" birthdate="2010-09-25" gender="M" nation="BRA" license="399739" swrid="5653294" athleteid="4606" externalid="399739">
              <RESULTS>
                <RESULT eventid="1104" points="308" swimtime="00:00:30.96" resultid="4607" heatid="5117" lane="7" entrytime="00:00:30.73" entrycourse="LCM" />
                <RESULT eventid="1151" points="259" swimtime="00:02:58.82" resultid="4608" heatid="5192" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.67" />
                    <SPLIT distance="100" swimtime="00:01:21.26" />
                    <SPLIT distance="150" swimtime="00:02:18.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="307" swimtime="00:01:16.48" resultid="4609" heatid="5257" lane="1" entrytime="00:01:17.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="340" swimtime="00:01:07.08" resultid="4610" heatid="5219" lane="4" entrytime="00:01:08.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="311" swimtime="00:00:34.73" resultid="4611" heatid="5284" lane="2" entrytime="00:00:41.30" entrycourse="LCM" />
                <RESULT eventid="1277" points="304" swimtime="00:02:46.41" resultid="4612" heatid="5345" lane="1" entrytime="00:02:51.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                    <SPLIT distance="100" swimtime="00:01:19.48" />
                    <SPLIT distance="150" swimtime="00:02:02.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietra" lastname="Vitoria Paczrowski" birthdate="2009-08-12" gender="F" nation="BRA" license="351253" swrid="5600275" athleteid="4481" externalid="351253" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1096" points="474" swimtime="00:00:30.28" resultid="4482" heatid="5103" lane="4" entrytime="00:00:29.63" entrycourse="LCM" />
                <RESULT eventid="1112" points="444" swimtime="00:02:27.92" resultid="4483" heatid="5144" lane="1" entrytime="00:02:24.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:09.11" />
                    <SPLIT distance="150" swimtime="00:01:48.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="376" swimtime="00:01:19.39" resultid="4484" heatid="5247" lane="8" entrytime="00:01:18.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="462" swimtime="00:01:06.85" resultid="4485" heatid="5207" lane="4" entrytime="00:01:06.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="435" swimtime="00:00:35.43" resultid="4486" heatid="5294" lane="3" entrytime="00:00:36.09" entrycourse="LCM" />
                <RESULT eventid="1305" points="339" swimtime="00:00:41.79" resultid="4487" heatid="5373" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alexandre" lastname="Celli Schneider" birthdate="2011-02-21" gender="M" nation="BRA" license="367055" swrid="5588587" athleteid="4519" externalid="367055">
              <RESULTS>
                <RESULT eventid="1151" points="310" swimtime="00:02:48.34" resultid="4520" heatid="5195" lane="8" entrytime="00:02:42.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:15.41" />
                    <SPLIT distance="150" swimtime="00:02:06.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="377" swimtime="00:01:11.42" resultid="4521" heatid="5257" lane="3" entrytime="00:01:11.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="373" swimtime="00:05:36.66" resultid="4522" heatid="5276" lane="2" entrytime="00:05:40.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:16.02" />
                    <SPLIT distance="150" swimtime="00:01:59.00" />
                    <SPLIT distance="200" swimtime="00:02:41.15" />
                    <SPLIT distance="250" swimtime="00:03:30.99" />
                    <SPLIT distance="300" swimtime="00:04:20.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="377" swimtime="00:00:32.59" resultid="4523" heatid="5285" lane="3" entrytime="00:00:33.74" entrycourse="LCM" />
                <RESULT eventid="1277" points="341" swimtime="00:02:40.13" resultid="4524" heatid="5346" lane="8" entrytime="00:02:37.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                    <SPLIT distance="100" swimtime="00:01:18.24" />
                    <SPLIT distance="150" swimtime="00:02:00.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1293" points="302" swimtime="00:02:44.35" resultid="4525" heatid="5358" lane="7" entrytime="00:03:01.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:20.09" />
                    <SPLIT distance="150" swimtime="00:02:04.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabrizio" lastname="Bulla Lanaro" birthdate="2009-08-28" gender="M" nation="BRA" license="344303" swrid="5559846" athleteid="4453" externalid="344303">
              <RESULTS>
                <RESULT eventid="1104" points="456" swimtime="00:00:27.15" resultid="4454" heatid="5124" lane="7" entrytime="00:00:26.96" entrycourse="LCM" />
                <RESULT eventid="1135" points="492" swimtime="00:01:02.60" resultid="4455" heatid="5174" lane="4" entrytime="00:01:02.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="488" swimtime="00:02:24.76" resultid="4456" heatid="5196" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.50" />
                    <SPLIT distance="150" swimtime="00:01:52.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="465" swimtime="00:01:06.59" resultid="4457" heatid="5260" lane="3" entrytime="00:01:07.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="454" swimtime="00:00:30.63" resultid="4458" heatid="5286" lane="4" entrytime="00:00:31.16" entrycourse="LCM" />
                <RESULT eventid="1267" points="519" swimtime="00:00:27.70" resultid="4459" heatid="5336" lane="5" entrytime="00:00:27.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Breno" lastname="Borges Piekarzievicz" birthdate="2011-11-11" gender="M" nation="BRA" license="403144" swrid="5676295" athleteid="4618" externalid="403144">
              <RESULTS>
                <RESULT eventid="1088" status="SICK" swimtime="00:00:00.00" resultid="4619" heatid="5079" lane="7" entrytime="00:01:45.57" entrycourse="LCM" />
                <RESULT eventid="1104" status="SICK" swimtime="00:00:00.00" resultid="4620" heatid="5115" lane="7" entrytime="00:00:37.40" entrycourse="LCM" />
                <RESULT eventid="1120" status="DNS" swimtime="00:00:00.00" resultid="4621" heatid="5148" lane="3" entrytime="00:03:07.17" entrycourse="LCM" />
                <RESULT eventid="1297" status="DNS" swimtime="00:00:00.00" resultid="4622" heatid="5366" lane="8" entrytime="00:00:51.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Cardim Martins" birthdate="2010-09-01" gender="F" nation="BRA" license="390920" swrid="5600130" athleteid="4644" externalid="390920">
              <RESULTS>
                <RESULT eventid="1064" points="321" swimtime="00:05:43.55" resultid="4645" heatid="5049" lane="1" entrytime="00:05:37.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                    <SPLIT distance="100" swimtime="00:01:18.80" />
                    <SPLIT distance="150" swimtime="00:02:01.87" />
                    <SPLIT distance="200" swimtime="00:02:45.92" />
                    <SPLIT distance="250" swimtime="00:03:30.09" />
                    <SPLIT distance="300" swimtime="00:04:15.63" />
                    <SPLIT distance="350" swimtime="00:04:59.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="346" swimtime="00:02:40.71" resultid="4646" heatid="5138" lane="5" entrytime="00:02:42.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.63" />
                    <SPLIT distance="100" swimtime="00:01:16.25" />
                    <SPLIT distance="150" swimtime="00:01:57.90" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 18:17), Na volta dos 150m (Medley Individual, Peito)." eventid="1143" status="DSQ" swimtime="00:03:13.53" resultid="4647" heatid="5186" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.48" />
                    <SPLIT distance="100" swimtime="00:01:29.46" />
                    <SPLIT distance="150" swimtime="00:02:31.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="304" swimtime="00:01:25.20" resultid="4648" heatid="5242" lane="3" entrytime="00:01:24.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="297" swimtime="00:00:40.25" resultid="4649" heatid="5293" lane="7" entrytime="00:00:39.90" entrycourse="LCM" />
                <RESULT eventid="1275" points="287" swimtime="00:03:06.50" resultid="4650" heatid="5340" lane="3" entrytime="00:03:01.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.96" />
                    <SPLIT distance="100" swimtime="00:01:30.88" />
                    <SPLIT distance="150" swimtime="00:02:19.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otto" lastname="Hedeke" birthdate="2011-03-24" gender="M" nation="BRA" license="372643" swrid="5588738" athleteid="4572" externalid="372643">
              <RESULTS>
                <RESULT eventid="1072" points="333" swimtime="00:05:17.22" resultid="4573" heatid="5057" lane="2" entrytime="00:05:26.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:13.79" />
                    <SPLIT distance="150" swimtime="00:01:54.59" />
                    <SPLIT distance="200" swimtime="00:02:35.73" />
                    <SPLIT distance="250" swimtime="00:03:16.44" />
                    <SPLIT distance="300" swimtime="00:03:57.29" />
                    <SPLIT distance="350" swimtime="00:04:38.04" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 6.5 - Não terminou a prova enquanto estava de costas.&#10;&#10;&#10;&#10;&#10;&#10;&#10;  (Horário: 18:47), Na volta dos 100m (Medley Individual, Costas)" eventid="1151" status="DSQ" swimtime="00:03:02.60" resultid="4574" heatid="5193" lane="6" entrytime="00:03:09.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.67" />
                    <SPLIT distance="100" swimtime="00:01:28.84" />
                    <SPLIT distance="150" swimtime="00:02:23.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="305" swimtime="00:01:09.59" resultid="4575" heatid="5219" lane="7" entrytime="00:01:15.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="328" swimtime="00:10:55.33" resultid="4576" heatid="5298" lane="1" entrytime="00:11:37.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                    <SPLIT distance="100" swimtime="00:01:15.82" />
                    <SPLIT distance="150" swimtime="00:01:57.10" />
                    <SPLIT distance="200" swimtime="00:02:38.20" />
                    <SPLIT distance="250" swimtime="00:03:19.97" />
                    <SPLIT distance="300" swimtime="00:04:00.99" />
                    <SPLIT distance="350" swimtime="00:04:42.90" />
                    <SPLIT distance="400" swimtime="00:05:24.79" />
                    <SPLIT distance="450" swimtime="00:06:06.77" />
                    <SPLIT distance="500" swimtime="00:06:48.91" />
                    <SPLIT distance="550" swimtime="00:07:30.28" />
                    <SPLIT distance="600" swimtime="00:08:13.26" />
                    <SPLIT distance="650" swimtime="00:08:53.86" />
                    <SPLIT distance="700" swimtime="00:09:35.63" />
                    <SPLIT distance="750" swimtime="00:10:16.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="323" swimtime="00:21:08.89" resultid="4577" heatid="5378" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.41" />
                    <SPLIT distance="100" swimtime="00:01:17.84" />
                    <SPLIT distance="150" swimtime="00:01:59.24" />
                    <SPLIT distance="200" swimtime="00:02:42.85" />
                    <SPLIT distance="250" swimtime="00:03:25.01" />
                    <SPLIT distance="300" swimtime="00:04:08.19" />
                    <SPLIT distance="350" swimtime="00:04:49.84" />
                    <SPLIT distance="400" swimtime="00:05:32.11" />
                    <SPLIT distance="450" swimtime="00:06:14.27" />
                    <SPLIT distance="500" swimtime="00:06:56.87" />
                    <SPLIT distance="550" swimtime="00:07:39.62" />
                    <SPLIT distance="600" swimtime="00:08:23.00" />
                    <SPLIT distance="650" swimtime="00:09:06.23" />
                    <SPLIT distance="700" swimtime="00:09:48.39" />
                    <SPLIT distance="750" swimtime="00:10:32.09" />
                    <SPLIT distance="800" swimtime="00:11:15.21" />
                    <SPLIT distance="850" swimtime="00:11:58.00" />
                    <SPLIT distance="900" swimtime="00:12:41.64" />
                    <SPLIT distance="950" swimtime="00:13:24.11" />
                    <SPLIT distance="1000" swimtime="00:14:07.42" />
                    <SPLIT distance="1050" swimtime="00:14:51.20" />
                    <SPLIT distance="1100" swimtime="00:15:33.89" />
                    <SPLIT distance="1150" swimtime="00:16:16.11" />
                    <SPLIT distance="1200" swimtime="00:16:58.88" />
                    <SPLIT distance="1250" swimtime="00:17:41.30" />
                    <SPLIT distance="1300" swimtime="00:18:23.63" />
                    <SPLIT distance="1350" swimtime="00:19:07.49" />
                    <SPLIT distance="1400" swimtime="00:19:50.57" />
                    <SPLIT distance="1450" swimtime="00:20:31.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Anna" lastname="Leticia Durat" birthdate="2008-02-09" gender="F" nation="BRA" license="331636" swrid="5600200" athleteid="4446" externalid="331636">
              <RESULTS>
                <RESULT eventid="1080" points="285" swimtime="00:01:37.35" resultid="4447" heatid="5068" lane="2" entrytime="00:01:30.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="411" swimtime="00:00:31.73" resultid="4448" heatid="5103" lane="1" entrytime="00:00:30.51" entrycourse="LCM" />
                <RESULT eventid="1112" points="302" swimtime="00:02:48.02" resultid="4449" heatid="5143" lane="1" entrytime="00:02:43.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="100" swimtime="00:01:18.67" />
                    <SPLIT distance="150" swimtime="00:02:03.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="386" swimtime="00:01:10.99" resultid="4450" heatid="5207" lane="1" entrytime="00:01:08.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="270" swimtime="00:03:32.62" resultid="4451" heatid="5311" lane="5" entrytime="00:03:16.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.97" />
                    <SPLIT distance="100" swimtime="00:01:37.99" />
                    <SPLIT distance="150" swimtime="00:02:33.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="349" swimtime="00:00:41.38" resultid="4452" heatid="5375" lane="4" entrytime="00:00:40.19" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kethelyn" lastname="Ribeiro Rodrigues" birthdate="2009-04-24" gender="F" nation="BRA" license="367052" swrid="5600244" athleteid="4505" externalid="367052">
              <RESULTS>
                <RESULT eventid="1064" points="372" swimtime="00:05:27.05" resultid="4506" heatid="5052" lane="4" entrytime="00:05:29.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:15.04" />
                    <SPLIT distance="150" swimtime="00:01:57.19" />
                    <SPLIT distance="200" swimtime="00:02:40.29" />
                    <SPLIT distance="250" swimtime="00:03:21.51" />
                    <SPLIT distance="300" swimtime="00:04:03.99" />
                    <SPLIT distance="350" swimtime="00:04:46.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="421" swimtime="00:00:31.49" resultid="4507" heatid="5102" lane="5" entrytime="00:00:31.32" entrycourse="LCM" />
                <RESULT eventid="1112" points="395" swimtime="00:02:33.78" resultid="4508" heatid="5143" lane="3" entrytime="00:02:29.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.81" />
                    <SPLIT distance="100" swimtime="00:01:13.96" />
                    <SPLIT distance="150" swimtime="00:01:53.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="434" swimtime="00:01:08.27" resultid="4509" heatid="5207" lane="2" entrytime="00:01:07.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="307" swimtime="00:00:39.79" resultid="4510" heatid="5289" lane="7" />
                <RESULT eventid="1275" points="277" swimtime="00:03:08.88" resultid="4511" heatid="5339" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                    <SPLIT distance="100" swimtime="00:01:31.33" />
                    <SPLIT distance="150" swimtime="00:02:21.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Pinterich Almeida" birthdate="2005-03-13" gender="M" nation="BRA" license="330749" swrid="5600235" athleteid="4498" externalid="330749">
              <RESULTS>
                <RESULT eventid="1120" points="652" swimtime="00:01:57.62" resultid="4499" heatid="5158" lane="3" entrytime="00:01:56.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.34" />
                    <SPLIT distance="100" swimtime="00:00:57.51" />
                    <SPLIT distance="150" swimtime="00:01:27.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="508" swimtime="00:02:22.82" resultid="4500" heatid="5200" lane="5" entrytime="00:02:23.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                    <SPLIT distance="100" swimtime="00:01:07.92" />
                    <SPLIT distance="150" swimtime="00:01:53.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="568" swimtime="00:01:02.28" resultid="4501" heatid="5263" lane="2" entrytime="00:01:01.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="648" swimtime="00:00:54.13" resultid="4502" heatid="5233" lane="2" entrytime="00:00:53.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="557" swimtime="00:09:09.34" resultid="4503" heatid="5297" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.58" />
                    <SPLIT distance="100" swimtime="00:01:03.15" />
                    <SPLIT distance="150" swimtime="00:01:38.41" />
                    <SPLIT distance="200" swimtime="00:02:13.78" />
                    <SPLIT distance="250" swimtime="00:02:49.55" />
                    <SPLIT distance="300" swimtime="00:03:24.75" />
                    <SPLIT distance="350" swimtime="00:03:59.91" />
                    <SPLIT distance="400" swimtime="00:04:35.38" />
                    <SPLIT distance="450" swimtime="00:05:10.10" />
                    <SPLIT distance="500" swimtime="00:05:45.22" />
                    <SPLIT distance="550" swimtime="00:06:20.07" />
                    <SPLIT distance="600" swimtime="00:06:54.84" />
                    <SPLIT distance="650" swimtime="00:07:29.40" />
                    <SPLIT distance="700" swimtime="00:08:04.06" />
                    <SPLIT distance="750" swimtime="00:08:37.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="539" swimtime="00:00:27.35" resultid="4504" heatid="5337" lane="1" entrytime="00:00:27.31" entrycourse="LCM" />
                <RESULT eventid="2351" swimtime="00:00:00.00" resultid="6124" entrytime="00:00:54.13" />
                <RESULT eventid="2359" points="524" swimtime="00:01:03.97" resultid="6148" heatid="6423" lane="7" entrytime="00:01:02.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Zanardi" birthdate="2008-10-02" gender="F" nation="BRA" license="398572" athleteid="4663" externalid="398572">
              <RESULTS>
                <RESULT eventid="1096" points="318" swimtime="00:00:34.57" resultid="4664" heatid="5101" lane="3" />
                <RESULT eventid="1112" points="315" swimtime="00:02:45.76" resultid="4665" heatid="5142" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.87" />
                    <SPLIT distance="100" swimtime="00:01:16.46" />
                    <SPLIT distance="150" swimtime="00:02:00.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="335" swimtime="00:01:14.45" resultid="4666" heatid="5206" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="245" swimtime="00:00:46.57" resultid="4667" heatid="5373" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Nalle Bejes" birthdate="2010-04-20" gender="F" nation="BRA" license="377323" swrid="5588826" athleteid="4585" externalid="377323">
              <RESULTS>
                <RESULT eventid="1080" points="405" swimtime="00:01:26.62" resultid="4586" heatid="5066" lane="4" entrytime="00:01:27.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="405" swimtime="00:02:32.45" resultid="4587" heatid="5139" lane="1" entrytime="00:02:34.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                    <SPLIT distance="100" swimtime="00:01:13.96" />
                    <SPLIT distance="150" swimtime="00:01:53.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="400" swimtime="00:02:51.15" resultid="4588" heatid="5187" lane="3" entrytime="00:02:57.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                    <SPLIT distance="100" swimtime="00:01:24.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="397" swimtime="00:01:10.30" resultid="4589" heatid="5203" lane="8" entrytime="00:01:10.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="361" swimtime="00:06:13.36" resultid="4590" heatid="5278" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                    <SPLIT distance="100" swimtime="00:01:28.54" />
                    <SPLIT distance="150" swimtime="00:02:17.71" />
                    <SPLIT distance="200" swimtime="00:03:06.78" />
                    <SPLIT distance="300" swimtime="00:04:48.05" />
                    <SPLIT distance="350" swimtime="00:05:31.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="385" swimtime="00:03:08.94" resultid="4591" heatid="5312" lane="6" entrytime="00:03:09.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.30" />
                    <SPLIT distance="100" swimtime="00:01:30.67" />
                    <SPLIT distance="150" swimtime="00:02:21.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Nogueira Silva" birthdate="2011-08-13" gender="M" nation="BRA" license="367150" swrid="5588832" athleteid="4539" externalid="367150">
              <RESULTS>
                <RESULT comment="SW 7.4 - Movimentos das pernas não simultâneos.  (Horário: 11:29)" eventid="1088" status="DSQ" swimtime="00:01:28.10" resultid="4540" heatid="5080" lane="7" entrytime="00:01:31.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="372" swimtime="00:02:21.70" resultid="4541" heatid="5151" lane="8" entrytime="00:02:22.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:08.87" />
                    <SPLIT distance="150" swimtime="00:01:46.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="382" swimtime="00:01:04.53" resultid="4542" heatid="5221" lane="3" entrytime="00:01:04.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="283" swimtime="00:00:39.48" resultid="4543" heatid="5365" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carol" lastname="Nalle Bejes" birthdate="2010-04-20" gender="F" nation="BRA" license="377315" swrid="5588824" athleteid="4578" externalid="377315">
              <RESULTS>
                <RESULT eventid="1080" points="437" swimtime="00:01:24.49" resultid="4579" heatid="5067" lane="6" entrytime="00:01:23.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" points="390" swimtime="00:05:21.93" resultid="4580" heatid="5049" lane="4" entrytime="00:05:14.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.37" />
                    <SPLIT distance="100" swimtime="00:01:13.99" />
                    <SPLIT distance="150" swimtime="00:01:54.43" />
                    <SPLIT distance="200" swimtime="00:02:36.91" />
                    <SPLIT distance="300" swimtime="00:04:01.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="453" swimtime="00:02:26.87" resultid="4581" heatid="5140" lane="4" entrytime="00:02:26.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:10.89" />
                    <SPLIT distance="150" swimtime="00:01:49.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="452" swimtime="00:01:07.35" resultid="4582" heatid="5204" lane="2" entrytime="00:01:07.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="420" swimtime="00:03:03.56" resultid="4583" heatid="5313" lane="5" entrytime="00:02:58.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.98" />
                    <SPLIT distance="100" swimtime="00:01:29.05" />
                    <SPLIT distance="150" swimtime="00:02:20.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="483" swimtime="00:00:37.14" resultid="4584" heatid="5376" lane="8" entrytime="00:00:39.66" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1235" points="506" swimtime="00:03:56.09" resultid="4671" heatid="5307" lane="6" entrytime="00:03:59.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.48" />
                    <SPLIT distance="100" swimtime="00:00:59.27" />
                    <SPLIT distance="150" swimtime="00:01:27.18" />
                    <SPLIT distance="200" swimtime="00:01:58.56" />
                    <SPLIT distance="250" swimtime="00:02:26.84" />
                    <SPLIT distance="300" swimtime="00:02:58.76" />
                    <SPLIT distance="350" swimtime="00:03:25.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4453" number="1" />
                    <RELAYPOSITION athleteid="4488" number="2" />
                    <RELAYPOSITION athleteid="4599" number="3" />
                    <RELAYPOSITION athleteid="4460" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1336" status="DNS" swimtime="00:00:00.00" resultid="4676" heatid="5387" lane="3" entrytime="00:04:25.95">
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4460" number="1" />
                    <RELAYPOSITION athleteid="4599" number="2" />
                    <RELAYPOSITION athleteid="4453" number="3" />
                    <RELAYPOSITION athleteid="4488" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1233" points="400" swimtime="00:04:15.44" resultid="4672" heatid="5306" lane="5" entrytime="00:04:02.75">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                    <SPLIT distance="100" swimtime="00:01:01.67" />
                    <SPLIT distance="150" swimtime="00:01:30.99" />
                    <SPLIT distance="200" swimtime="00:02:03.07" />
                    <SPLIT distance="250" swimtime="00:02:34.51" />
                    <SPLIT distance="300" swimtime="00:03:08.32" />
                    <SPLIT distance="350" swimtime="00:03:39.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4526" number="1" />
                    <RELAYPOSITION athleteid="4651" number="2" />
                    <RELAYPOSITION athleteid="4592" number="3" />
                    <RELAYPOSITION athleteid="4606" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1334" points="362" swimtime="00:04:50.06" resultid="4675" heatid="5386" lane="4" entrytime="00:04:26.48">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.98" />
                    <SPLIT distance="150" swimtime="00:01:55.84" />
                    <SPLIT distance="200" swimtime="00:02:42.73" />
                    <SPLIT distance="250" swimtime="00:03:12.74" />
                    <SPLIT distance="300" swimtime="00:03:49.00" />
                    <SPLIT distance="350" swimtime="00:04:18.39" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4606" number="1" />
                    <RELAYPOSITION athleteid="4658" number="2" />
                    <RELAYPOSITION athleteid="4526" number="3" />
                    <RELAYPOSITION athleteid="4651" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1231" points="398" swimtime="00:04:15.70" resultid="4673" heatid="5305" lane="6" entrytime="00:04:32.37">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:04.64" />
                    <SPLIT distance="150" swimtime="00:01:35.62" />
                    <SPLIT distance="200" swimtime="00:02:08.66" />
                    <SPLIT distance="250" swimtime="00:02:38.54" />
                    <SPLIT distance="300" swimtime="00:03:12.08" />
                    <SPLIT distance="350" swimtime="00:03:41.89" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4558" number="1" />
                    <RELAYPOSITION athleteid="4539" number="2" />
                    <RELAYPOSITION athleteid="4613" number="3" />
                    <RELAYPOSITION athleteid="4519" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1332" points="357" swimtime="00:04:51.44" resultid="4674" heatid="5385" lane="3" entrytime="00:05:01.68">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                    <SPLIT distance="100" swimtime="00:01:13.36" />
                    <SPLIT distance="150" swimtime="00:01:51.40" />
                    <SPLIT distance="200" swimtime="00:02:38.28" />
                    <SPLIT distance="250" swimtime="00:03:09.67" />
                    <SPLIT distance="300" swimtime="00:03:48.18" />
                    <SPLIT distance="350" swimtime="00:04:18.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4519" number="1" />
                    <RELAYPOSITION athleteid="4533" number="2" />
                    <RELAYPOSITION athleteid="4613" number="3" />
                    <RELAYPOSITION athleteid="4558" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1223" points="518" swimtime="00:04:18.89" resultid="4668" heatid="5303" lane="3" entrytime="00:04:16.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                    <SPLIT distance="150" swimtime="00:01:31.72" />
                    <SPLIT distance="200" swimtime="00:02:06.53" />
                    <SPLIT distance="250" swimtime="00:02:38.06" />
                    <SPLIT distance="300" swimtime="00:03:11.02" />
                    <SPLIT distance="350" swimtime="00:03:42.45" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4418" number="1" />
                    <RELAYPOSITION athleteid="4481" number="2" />
                    <RELAYPOSITION athleteid="4467" number="3" />
                    <RELAYPOSITION athleteid="4505" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1221" points="432" swimtime="00:04:35.04" resultid="4669" heatid="5302" lane="5" entrytime="00:04:21.61">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                    <SPLIT distance="100" swimtime="00:01:07.83" />
                    <SPLIT distance="150" swimtime="00:01:39.66" />
                    <SPLIT distance="200" swimtime="00:02:15.28" />
                    <SPLIT distance="250" swimtime="00:02:48.53" />
                    <SPLIT distance="300" swimtime="00:03:25.35" />
                    <SPLIT distance="350" swimtime="00:03:58.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4544" number="1" />
                    <RELAYPOSITION athleteid="4578" number="2" />
                    <RELAYPOSITION athleteid="4637" number="3" />
                    <RELAYPOSITION athleteid="4585" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1322" points="383" swimtime="00:05:17.05" resultid="4670" heatid="5382" lane="5" entrytime="00:05:04.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.44" />
                    <SPLIT distance="100" swimtime="00:01:27.08" />
                    <SPLIT distance="150" swimtime="00:02:05.90" />
                    <SPLIT distance="200" swimtime="00:02:50.91" />
                    <SPLIT distance="250" swimtime="00:03:26.23" />
                    <SPLIT distance="350" swimtime="00:04:40.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4644" number="1" />
                    <RELAYPOSITION athleteid="4578" number="2" />
                    <RELAYPOSITION athleteid="4544" number="3" />
                    <RELAYPOSITION athleteid="4637" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1287" points="368" swimtime="00:05:03.57" resultid="4677" heatid="5354" lane="5" entrytime="00:04:28.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.99" />
                    <SPLIT distance="150" swimtime="00:02:10.78" />
                    <SPLIT distance="200" swimtime="00:03:02.51" />
                    <SPLIT distance="250" swimtime="00:03:31.89" />
                    <SPLIT distance="300" swimtime="00:04:08.29" />
                    <SPLIT distance="350" swimtime="00:04:34.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4663" number="1" />
                    <RELAYPOSITION athleteid="4446" number="2" />
                    <RELAYPOSITION athleteid="4439" number="3" />
                    <RELAYPOSITION athleteid="4474" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1285" points="512" swimtime="00:04:31.81" resultid="4678" heatid="5353" lane="7" entrytime="00:05:04.38">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:06.91" />
                    <SPLIT distance="150" swimtime="00:01:42.09" />
                    <SPLIT distance="200" swimtime="00:02:19.75" />
                    <SPLIT distance="250" swimtime="00:02:51.12" />
                    <SPLIT distance="350" swimtime="00:03:58.37" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4460" number="1" />
                    <RELAYPOSITION athleteid="4599" number="2" />
                    <RELAYPOSITION athleteid="4418" number="3" />
                    <RELAYPOSITION athleteid="4467" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1283" points="407" swimtime="00:04:53.37" resultid="4679" heatid="5352" lane="4" entrytime="00:04:33.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                    <SPLIT distance="100" swimtime="00:01:15.70" />
                    <SPLIT distance="150" swimtime="00:01:55.58" />
                    <SPLIT distance="200" swimtime="00:02:41.04" />
                    <SPLIT distance="250" swimtime="00:03:10.38" />
                    <SPLIT distance="300" swimtime="00:03:46.29" />
                    <SPLIT distance="350" swimtime="00:04:18.24" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4606" number="1" />
                    <RELAYPOSITION athleteid="4578" number="2" />
                    <RELAYPOSITION athleteid="4526" number="3" />
                    <RELAYPOSITION athleteid="4544" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1281" points="358" swimtime="00:05:06.37" resultid="4680" heatid="5351" lane="7" entrytime="00:05:15.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.42" />
                    <SPLIT distance="100" swimtime="00:01:11.85" />
                    <SPLIT distance="150" swimtime="00:01:54.40" />
                    <SPLIT distance="200" swimtime="00:02:41.55" />
                    <SPLIT distance="250" swimtime="00:03:12.69" />
                    <SPLIT distance="300" swimtime="00:03:51.00" />
                    <SPLIT distance="350" swimtime="00:04:25.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4519" number="1" />
                    <RELAYPOSITION athleteid="4565" number="2" />
                    <RELAYPOSITION athleteid="4613" number="3" />
                    <RELAYPOSITION athleteid="4512" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1285" points="440" swimtime="00:04:46.04" resultid="4681" heatid="5353" lane="6" entrytime="00:04:35.37">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:18.14" />
                    <SPLIT distance="150" swimtime="00:01:53.12" />
                    <SPLIT distance="200" swimtime="00:02:35.76" />
                    <SPLIT distance="250" swimtime="00:03:04.10" />
                    <SPLIT distance="300" swimtime="00:03:37.82" />
                    <SPLIT distance="350" swimtime="00:04:10.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4481" number="1" />
                    <RELAYPOSITION athleteid="4488" number="2" />
                    <RELAYPOSITION athleteid="4453" number="3" />
                    <RELAYPOSITION athleteid="4505" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="SANTA MÔNICA &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1283" points="318" swimtime="00:05:18.66" resultid="4682" heatid="5352" lane="7" entrytime="00:04:55.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                    <SPLIT distance="150" swimtime="00:02:09.07" />
                    <SPLIT distance="200" swimtime="00:02:55.11" />
                    <SPLIT distance="250" swimtime="00:03:30.60" />
                    <SPLIT distance="300" swimtime="00:04:09.32" />
                    <SPLIT distance="350" swimtime="00:04:41.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4585" number="1" />
                    <RELAYPOSITION athleteid="4658" number="2" />
                    <RELAYPOSITION athleteid="4592" number="3" />
                    <RELAYPOSITION athleteid="4637" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="10443" nation="BRA" region="SC" clubid="4228" swrid="93763" name="Associação Joinvilense De Natação" shortname="Joinville Natação">
          <ATHLETES>
            <ATHLETE firstname="Guilherme" lastname="Furlan" birthdate="2006-06-16" gender="M" nation="BRA" license="369512" swrid="5682812" athleteid="4229" externalid="369512">
              <RESULTS>
                <RESULT eventid="1104" points="529" status="EXH" swimtime="00:00:25.84" resultid="4230" heatid="5129" lane="7" entrytime="00:00:25.34" entrycourse="LCM" />
                <RESULT eventid="1167" points="609" status="EXH" swimtime="00:00:55.27" resultid="4231" heatid="5232" lane="6" entrytime="00:00:55.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.04" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="11303" nation="BRA" region="PR" clubid="2874" swrid="93760" name="Associação De Talentos Da Natação" shortname="Atn/Curitiba">
          <ATHLETES>
            <ATHLETE firstname="Murilo" lastname="Iglesias Prado" birthdate="2010-06-15" gender="M" nation="BRA" license="408052" swrid="5723025" athleteid="3015" externalid="408052">
              <RESULTS>
                <RESULT eventid="1104" points="339" swimtime="00:00:29.98" resultid="3016" heatid="5117" lane="2" entrytime="00:00:30.45" entrycourse="LCM" />
                <RESULT eventid="1120" points="247" swimtime="00:02:42.54" resultid="3017" heatid="5149" lane="6" entrytime="00:02:37.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.90" />
                    <SPLIT distance="100" swimtime="00:01:16.22" />
                    <SPLIT distance="150" swimtime="00:02:00.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="336" swimtime="00:01:07.34" resultid="3018" heatid="5220" lane="5" entrytime="00:01:07.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="282" swimtime="00:00:35.88" resultid="3019" heatid="5284" lane="6" entrytime="00:00:38.27" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fabiana" lastname="Zaleski Dallazem" birthdate="2009-05-16" gender="F" nation="BRA" license="344287" swrid="5600279" athleteid="2875" externalid="344287" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1143" points="495" swimtime="00:02:39.34" resultid="2876" heatid="5190" lane="3" entrytime="00:02:41.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                    <SPLIT distance="100" swimtime="00:01:13.50" />
                    <SPLIT distance="150" swimtime="00:02:03.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="570" swimtime="00:01:09.13" resultid="2877" heatid="5247" lane="3" entrytime="00:01:10.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="579" swimtime="00:00:32.22" resultid="2878" heatid="5295" lane="2" entrytime="00:00:32.75" entrycourse="LCM" />
                <RESULT eventid="1275" points="486" swimtime="00:02:36.59" resultid="2879" heatid="5343" lane="3" entrytime="00:02:33.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="100" swimtime="00:01:15.95" />
                    <SPLIT distance="150" swimtime="00:01:57.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2391" points="568" swimtime="00:01:09.21" resultid="6128" heatid="6424" lane="5" entrytime="00:01:09.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Camila" lastname="Duarte De Almeida" birthdate="2009-11-26" gender="F" nation="BRA" license="378819" swrid="5600152" athleteid="2946" externalid="378819">
              <RESULTS>
                <RESULT eventid="1096" points="485" swimtime="00:00:30.05" resultid="2947" heatid="5103" lane="3" entrytime="00:00:30.06" entrycourse="LCM" />
                <RESULT eventid="1112" points="415" swimtime="00:02:31.29" resultid="2948" heatid="5143" lane="2" entrytime="00:02:30.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:10.99" />
                    <SPLIT distance="150" swimtime="00:01:50.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="472" swimtime="00:01:06.40" resultid="2949" heatid="5207" lane="5" entrytime="00:01:06.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="371" swimtime="00:00:33.98" resultid="2950" heatid="5325" lane="6" entrytime="00:00:34.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Kerppers Kreia" birthdate="2006-12-01" gender="M" nation="BRA" license="366815" swrid="5600195" athleteid="2897" externalid="366815">
              <RESULTS>
                <RESULT eventid="1104" points="461" swimtime="00:00:27.06" resultid="2898" heatid="5128" lane="2" entrytime="00:00:27.25" entrycourse="LCM" />
                <RESULT eventid="1120" points="482" swimtime="00:02:10.04" resultid="2899" heatid="5158" lane="8" entrytime="00:02:11.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.26" />
                    <SPLIT distance="100" swimtime="00:01:01.95" />
                    <SPLIT distance="150" swimtime="00:01:35.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="524" swimtime="00:00:58.10" resultid="2900" heatid="5231" lane="4" entrytime="00:00:58.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="403" swimtime="00:00:30.14" resultid="2901" heatid="5330" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Rosa Pech" birthdate="2010-10-26" gender="M" nation="BRA" license="413378" swrid="5755377" athleteid="3020" externalid="413378">
              <RESULTS>
                <RESULT eventid="1088" points="190" swimtime="00:01:38.87" resultid="3021" heatid="5079" lane="2" entrytime="00:01:44.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="189" swimtime="00:00:36.38" resultid="3022" heatid="5115" lane="5" entrytime="00:00:35.73" entrycourse="LCM" />
                <RESULT eventid="1167" points="193" swimtime="00:01:21.03" resultid="3023" heatid="5217" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada.  (Horário: 16:47)" eventid="1297" status="DSQ" swimtime="00:00:44.62" resultid="3024" heatid="5365" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Yuji Yamazato" birthdate="2008-10-01" gender="M" nation="BRA" license="392664" swrid="5622313" athleteid="2985" externalid="392664">
              <RESULTS>
                <RESULT eventid="1104" points="390" swimtime="00:00:28.61" resultid="2986" heatid="5122" lane="3" entrytime="00:00:28.69" entrycourse="LCM" />
                <RESULT comment="SW 10.2 - Não completou a distância total da prova.  (Horário: 18:01)" eventid="1135" status="DSQ" swimtime="00:00:00.00" resultid="2987" heatid="5173" lane="1" entrytime="00:01:24.30" entrycourse="LCM" />
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 9:50)" eventid="1167" status="DSQ" swimtime="00:01:03.97" resultid="2988" heatid="5226" lane="1" entrytime="00:01:03.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="376" swimtime="00:00:30.83" resultid="2989" heatid="5333" lane="6" entrytime="00:00:31.01" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Riccieri" lastname="Rodrigues Muzolon" birthdate="2010-11-08" gender="M" nation="BRA" license="385439" swrid="5588887" athleteid="2951" externalid="385439">
              <RESULTS>
                <RESULT eventid="1088" points="264" swimtime="00:01:28.64" resultid="2952" heatid="5081" lane="7" entrytime="00:01:28.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="359" swimtime="00:00:29.40" resultid="2953" heatid="5118" lane="2" entrytime="00:00:29.60" entrycourse="LCM" />
                <RESULT eventid="1120" points="287" swimtime="00:02:34.55" resultid="2954" heatid="5149" lane="7" entrytime="00:02:37.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.82" />
                    <SPLIT distance="100" swimtime="00:01:10.78" />
                    <SPLIT distance="150" swimtime="00:01:51.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="285" swimtime="00:01:18.35" resultid="2955" heatid="5256" lane="5" entrytime="00:01:19.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="292" swimtime="00:00:35.49" resultid="2956" heatid="5285" lane="8" entrytime="00:00:36.34" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Garcia Fraga" birthdate="2003-10-07" gender="M" nation="BRA" license="283467" swrid="5717265" athleteid="2889" externalid="283467" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1251" points="444" swimtime="00:02:44.41" resultid="2890" heatid="5319" lane="1" entrytime="00:02:44.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                    <SPLIT distance="100" swimtime="00:01:15.33" />
                    <SPLIT distance="150" swimtime="00:01:58.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="422" swimtime="00:02:29.15" resultid="2891" heatid="5347" lane="8" entrytime="00:02:27.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                    <SPLIT distance="100" swimtime="00:01:12.55" />
                    <SPLIT distance="150" swimtime="00:01:51.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Garcia De Fraga" birthdate="2009-03-24" gender="M" nation="BRA" license="342147" swrid="5600172" athleteid="2880" externalid="342147" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1151" points="599" swimtime="00:02:15.18" resultid="2881" heatid="5198" lane="3" entrytime="00:02:16.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.21" />
                    <SPLIT distance="100" swimtime="00:01:02.11" />
                    <SPLIT distance="150" swimtime="00:01:43.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="628" swimtime="00:01:00.25" resultid="2882" heatid="5261" lane="5" entrytime="00:01:01.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.97" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 6.3 - A cabeça não rompeu a superfície da água no ou antes do marco de 15m após o início ou a virada.  (Horário: 17:47)" eventid="1213" status="DSQ" swimtime="00:00:28.21" resultid="2883" heatid="5287" lane="2" entrytime="00:00:29.91" entrycourse="LCM" />
                <RESULT eventid="1277" points="596" swimtime="00:02:12.97" resultid="2884" heatid="5348" lane="6" entrytime="00:02:13.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.95" />
                    <SPLIT distance="100" swimtime="00:01:04.85" />
                    <SPLIT distance="150" swimtime="00:01:38.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2359" points="630" swimtime="00:01:00.18" resultid="6144" heatid="6423" lane="6" entrytime="00:01:00.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mauricio" lastname="Furtado Niwa" birthdate="1978-05-30" gender="M" nation="BRA" license="398757" swrid="5653291" athleteid="2909" externalid="398757">
              <RESULTS>
                <RESULT eventid="1135" points="486" swimtime="00:01:02.87" resultid="2910" heatid="5177" lane="3" entrytime="00:01:01.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="517" swimtime="00:00:58.37" resultid="2911" heatid="5232" lane="8" entrytime="00:00:58.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="517" swimtime="00:00:27.73" resultid="2912" heatid="5336" lane="6" entrytime="00:00:27.68" entrycourse="LCM" />
                <RESULT eventid="1293" points="382" swimtime="00:02:32.02" resultid="2913" heatid="5359" lane="6" entrytime="00:02:31.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.60" />
                    <SPLIT distance="100" swimtime="00:01:12.56" />
                    <SPLIT distance="150" swimtime="00:01:54.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Neves Vianna" birthdate="2007-12-30" gender="F" nation="BRA" license="391106" swrid="5600223" athleteid="2968" externalid="391106">
              <RESULTS>
                <RESULT eventid="1096" points="293" swimtime="00:00:35.53" resultid="2969" heatid="5105" lane="4" entrytime="00:00:36.00" entrycourse="LCM" />
                <RESULT eventid="1112" points="239" swimtime="00:03:01.69" resultid="2970" heatid="5145" lane="5" entrytime="00:02:58.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.62" />
                    <SPLIT distance="100" swimtime="00:01:26.38" />
                    <SPLIT distance="150" swimtime="00:02:14.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="241" swimtime="00:01:32.09" resultid="2971" heatid="5248" lane="7" entrytime="00:01:32.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="244" swimtime="00:00:42.96" resultid="2972" heatid="5292" lane="2" entrytime="00:00:43.30" entrycourse="LCM" />
                <RESULT eventid="1259" points="164" swimtime="00:00:44.61" resultid="2973" heatid="5323" lane="8" entrytime="00:00:48.13" entrycourse="LCM" />
                <RESULT eventid="1275" points="212" swimtime="00:03:26.36" resultid="2974" heatid="5340" lane="1" entrytime="00:03:20.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.80" />
                    <SPLIT distance="100" swimtime="00:01:40.16" />
                    <SPLIT distance="150" swimtime="00:02:34.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Kerniski Demantova" birthdate="1982-05-25" gender="M" nation="BRA" license="398222" swrid="5653293" athleteid="2902" externalid="398222">
              <RESULTS>
                <RESULT eventid="1072" points="392" swimtime="00:05:00.49" resultid="2903" heatid="5064" lane="1" entrytime="00:04:59.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                    <SPLIT distance="100" swimtime="00:01:08.53" />
                    <SPLIT distance="150" swimtime="00:01:45.57" />
                    <SPLIT distance="200" swimtime="00:02:24.45" />
                    <SPLIT distance="250" swimtime="00:03:02.72" />
                    <SPLIT distance="300" swimtime="00:03:42.80" />
                    <SPLIT distance="350" swimtime="00:04:21.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="342" swimtime="00:10:46.44" resultid="2904" heatid="5299" lane="1" entrytime="00:10:20.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.26" />
                    <SPLIT distance="100" swimtime="00:01:13.59" />
                    <SPLIT distance="150" swimtime="00:01:53.44" />
                    <SPLIT distance="200" swimtime="00:02:33.72" />
                    <SPLIT distance="250" swimtime="00:03:14.33" />
                    <SPLIT distance="300" swimtime="00:03:54.69" />
                    <SPLIT distance="350" swimtime="00:04:35.30" />
                    <SPLIT distance="450" swimtime="00:05:57.26" />
                    <SPLIT distance="500" swimtime="00:06:38.14" />
                    <SPLIT distance="550" swimtime="00:07:19.51" />
                    <SPLIT distance="600" swimtime="00:08:00.90" />
                    <SPLIT distance="650" swimtime="00:08:42.54" />
                    <SPLIT distance="700" swimtime="00:09:24.37" />
                    <SPLIT distance="750" swimtime="00:10:06.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="354" swimtime="00:20:30.16" resultid="2905" heatid="5379" lane="6" entrytime="00:20:14.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.05" />
                    <SPLIT distance="100" swimtime="00:01:15.10" />
                    <SPLIT distance="150" swimtime="00:01:55.53" />
                    <SPLIT distance="250" swimtime="00:03:16.52" />
                    <SPLIT distance="300" swimtime="00:03:56.97" />
                    <SPLIT distance="350" swimtime="00:04:37.83" />
                    <SPLIT distance="400" swimtime="00:05:18.59" />
                    <SPLIT distance="450" swimtime="00:05:59.64" />
                    <SPLIT distance="500" swimtime="00:06:40.27" />
                    <SPLIT distance="550" swimtime="00:07:21.21" />
                    <SPLIT distance="600" swimtime="00:08:01.80" />
                    <SPLIT distance="650" swimtime="00:08:42.93" />
                    <SPLIT distance="700" swimtime="00:09:24.38" />
                    <SPLIT distance="750" swimtime="00:10:05.81" />
                    <SPLIT distance="800" swimtime="00:10:47.32" />
                    <SPLIT distance="850" swimtime="00:11:29.02" />
                    <SPLIT distance="900" swimtime="00:12:10.76" />
                    <SPLIT distance="950" swimtime="00:12:52.54" />
                    <SPLIT distance="1000" swimtime="00:13:33.59" />
                    <SPLIT distance="1050" swimtime="00:14:15.23" />
                    <SPLIT distance="1100" swimtime="00:14:57.27" />
                    <SPLIT distance="1150" swimtime="00:15:38.79" />
                    <SPLIT distance="1200" swimtime="00:16:20.26" />
                    <SPLIT distance="1250" swimtime="00:17:02.02" />
                    <SPLIT distance="1300" swimtime="00:17:43.75" />
                    <SPLIT distance="1350" swimtime="00:18:26.61" />
                    <SPLIT distance="1400" swimtime="00:19:09.20" />
                    <SPLIT distance="1450" swimtime="00:19:50.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Zaleski Dallazem" birthdate="2009-05-16" gender="M" nation="BRA" license="344286" swrid="5600280" athleteid="2914" externalid="344286" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1088" points="427" swimtime="00:01:15.53" resultid="2915" heatid="5084" lane="3" entrytime="00:01:15.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="371" swimtime="00:01:08.80" resultid="2916" heatid="5173" lane="6" entrytime="00:01:12.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="476" swimtime="00:00:59.98" resultid="2917" heatid="5227" lane="2" entrytime="00:01:00.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="421" swimtime="00:02:47.38" resultid="2918" heatid="5318" lane="2" entrytime="00:02:49.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="100" swimtime="00:01:21.02" />
                    <SPLIT distance="150" swimtime="00:02:04.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="422" swimtime="00:00:34.59" resultid="2919" heatid="5369" lane="3" entrytime="00:00:34.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Fonseca Vendramin" birthdate="2008-09-28" gender="F" nation="BRA" license="393918" swrid="5622282" athleteid="2990" externalid="393918">
              <RESULTS>
                <RESULT eventid="1096" points="419" swimtime="00:00:31.55" resultid="2991" heatid="5102" lane="6" entrytime="00:00:31.84" entrycourse="LCM" />
                <RESULT eventid="1159" points="395" swimtime="00:01:10.46" resultid="2992" heatid="5206" lane="4" entrytime="00:01:10.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="304" swimtime="00:00:36.31" resultid="2993" heatid="5324" lane="6" entrytime="00:00:36.37" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Muller" birthdate="2009-10-10" gender="F" nation="BRA" license="376952" swrid="5600221" athleteid="2941" externalid="376952">
              <RESULTS>
                <RESULT eventid="1080" points="531" swimtime="00:01:19.17" resultid="2942" heatid="5069" lane="7" entrytime="00:01:20.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="387" swimtime="00:02:52.97" resultid="2943" heatid="5189" lane="5" entrytime="00:02:50.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.18" />
                    <SPLIT distance="100" swimtime="00:01:26.77" />
                    <SPLIT distance="150" swimtime="00:02:12.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="448" swimtime="00:02:59.63" resultid="2944" heatid="5313" lane="2" entrytime="00:02:59.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.37" />
                    <SPLIT distance="100" swimtime="00:01:24.71" />
                    <SPLIT distance="150" swimtime="00:02:12.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="514" swimtime="00:00:36.39" resultid="2945" heatid="5377" lane="6" entrytime="00:00:36.62" entrycourse="LCM" />
                <RESULT eventid="2312" points="521" swimtime="00:01:19.67" resultid="5943" heatid="6416" lane="2" entrytime="00:01:19.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Arthur Ribeiro" birthdate="2010-02-05" gender="M" nation="BRA" license="408025" swrid="5723020" athleteid="3009" externalid="408025">
              <RESULTS>
                <RESULT eventid="1088" points="301" swimtime="00:01:24.79" resultid="3010" heatid="5081" lane="3" entrytime="00:01:26.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="310" swimtime="00:00:30.87" resultid="3011" heatid="5117" lane="5" entrytime="00:00:30.23" entrycourse="LCM" />
                <RESULT eventid="1167" points="311" swimtime="00:01:09.15" resultid="3012" heatid="5220" lane="7" entrytime="00:01:08.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="281" swimtime="00:03:11.40" resultid="3013" heatid="5315" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.72" />
                    <SPLIT distance="100" swimtime="00:01:34.26" />
                    <SPLIT distance="150" swimtime="00:02:25.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="320" swimtime="00:00:37.92" resultid="3014" heatid="5367" lane="3" entrytime="00:00:38.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Angelo" lastname="De Queiroz Neto" birthdate="2003-10-31" gender="M" nation="BRA" license="342814" swrid="5600149" athleteid="2892" externalid="342814" level="AERC">
              <RESULTS>
                <RESULT eventid="1135" points="426" swimtime="00:01:05.71" resultid="2893" heatid="5176" lane="4" entrytime="00:01:07.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" status="DNS" swimtime="00:00:00.00" resultid="2894" heatid="5262" lane="7" />
                <RESULT eventid="1213" points="347" swimtime="00:00:33.49" resultid="2895" heatid="5282" lane="3" />
                <RESULT eventid="1267" points="441" swimtime="00:00:29.25" resultid="2896" heatid="5334" lane="1" entrytime="00:00:29.73" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Castellano Purkot" birthdate="2010-01-25" gender="M" nation="BRA" license="392484" swrid="5622268" athleteid="2980" externalid="392484">
              <RESULTS>
                <RESULT eventid="1088" points="243" swimtime="00:01:31.07" resultid="2981" heatid="5080" lane="8" entrytime="00:01:32.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="314" swimtime="00:00:30.75" resultid="2982" heatid="5117" lane="6" entrytime="00:00:30.44" entrycourse="LCM" />
                <RESULT eventid="1167" points="307" swimtime="00:01:09.46" resultid="2983" heatid="5220" lane="8" entrytime="00:01:08.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="275" swimtime="00:00:39.86" resultid="2984" heatid="5367" lane="8" entrytime="00:00:40.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Freitas Szucs" birthdate="2011-10-02" gender="M" nation="BRA" license="377272" swrid="5588708" athleteid="2926" externalid="377272">
              <RESULTS>
                <RESULT eventid="1104" points="241" swimtime="00:00:33.59" resultid="2927" heatid="5116" lane="1" entrytime="00:00:33.90" entrycourse="LCM" />
                <RESULT eventid="1167" points="235" swimtime="00:01:15.91" resultid="2928" heatid="5219" lane="1" entrytime="00:01:16.00" entrycourse="LCM" />
                <RESULT eventid="1267" points="193" swimtime="00:00:38.51" resultid="2929" heatid="5331" lane="8" entrytime="00:00:39.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcos" lastname="Demchuk" birthdate="2011-06-15" gender="M" nation="BRA" license="388540" swrid="5602530" athleteid="2957" externalid="388540">
              <RESULTS>
                <RESULT eventid="1104" points="316" swimtime="00:00:30.68" resultid="2958" heatid="5117" lane="1" entrytime="00:00:30.85" entrycourse="LCM" />
                <RESULT eventid="1151" points="221" swimtime="00:03:08.55" resultid="2959" heatid="5192" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.18" />
                    <SPLIT distance="100" swimtime="00:01:30.31" />
                    <SPLIT distance="150" swimtime="00:02:27.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="310" swimtime="00:01:09.22" resultid="2960" heatid="5219" lane="5" entrytime="00:01:09.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="192" swimtime="00:00:38.55" resultid="2961" heatid="5329" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelo" lastname="Correia Bonfim" birthdate="2009-06-21" gender="M" nation="BRA" license="391663" swrid="5622271" athleteid="2975" externalid="391663">
              <RESULTS>
                <RESULT eventid="1104" points="408" swimtime="00:00:28.18" resultid="2976" heatid="5123" lane="2" entrytime="00:00:28.01" entrycourse="LCM" />
                <RESULT eventid="1120" points="371" swimtime="00:02:21.85" resultid="2977" heatid="5153" lane="5" entrytime="00:02:24.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                    <SPLIT distance="100" swimtime="00:01:06.64" />
                    <SPLIT distance="150" swimtime="00:01:43.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="432" swimtime="00:01:01.98" resultid="2978" heatid="5226" lane="5" entrytime="00:01:01.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="340" swimtime="00:00:31.90" resultid="2979" heatid="5332" lane="4" entrytime="00:00:31.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Sofia Silva" birthdate="2007-05-28" gender="F" nation="BRA" license="390921" swrid="5600260" athleteid="2962" externalid="390921">
              <RESULTS>
                <RESULT eventid="1080" points="234" swimtime="00:01:44.03" resultid="2963" heatid="5070" lane="2" entrytime="00:01:43.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="226" swimtime="00:03:26.85" resultid="2964" heatid="5191" lane="1" entrytime="00:03:23.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.43" />
                    <SPLIT distance="100" swimtime="00:01:39.11" />
                    <SPLIT distance="150" swimtime="00:02:38.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="239" swimtime="00:01:23.23" resultid="2965" heatid="5209" lane="1" entrytime="00:01:24.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="155" swimtime="00:00:45.47" resultid="2966" heatid="5322" lane="1" />
                <RESULT eventid="1243" points="216" swimtime="00:03:48.97" resultid="2967" heatid="5311" lane="8" entrytime="00:03:42.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.68" />
                    <SPLIT distance="100" swimtime="00:01:47.68" />
                    <SPLIT distance="150" swimtime="00:02:47.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="James" lastname="Roberto Zoschke" birthdate="1976-02-08" gender="M" nation="BRA" license="312251" swrid="5688617" athleteid="2906" externalid="312251">
              <RESULTS>
                <RESULT comment="SW 7.4 - Movimentos das pernas não simultâneos.  (Horário: 11:47)" eventid="1088" status="DSQ" swimtime="00:01:15.04" resultid="2907" heatid="5087" lane="1" entrytime="00:01:14.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="470" swimtime="00:00:33.36" resultid="2908" heatid="5370" lane="2" entrytime="00:00:33.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Bortoleto" birthdate="2008-09-05" gender="M" nation="BRA" license="406709" swrid="5717249" athleteid="2994" externalid="406709">
              <RESULTS>
                <RESULT eventid="1104" points="452" swimtime="00:00:27.24" resultid="2995" heatid="5124" lane="8" entrytime="00:00:27.35" entrycourse="LCM" />
                <RESULT eventid="1120" points="423" swimtime="00:02:15.85" resultid="2996" heatid="5155" lane="1" entrytime="00:02:15.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.78" />
                    <SPLIT distance="100" swimtime="00:01:05.95" />
                    <SPLIT distance="150" swimtime="00:01:41.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="474" swimtime="00:01:00.08" resultid="2997" heatid="5227" lane="5" entrytime="00:00:59.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="378" swimtime="00:00:30.78" resultid="2998" heatid="5333" lane="3" entrytime="00:00:30.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Navarro Silva" birthdate="2011-01-10" gender="F" nation="BRA" license="406711" swrid="5717284" athleteid="2999" externalid="406711">
              <RESULTS>
                <RESULT eventid="1096" points="366" swimtime="00:00:32.98" resultid="3000" heatid="5097" lane="6" entrytime="00:00:34.90" entrycourse="LCM" />
                <RESULT eventid="1175" points="299" swimtime="00:01:25.71" resultid="3001" heatid="5242" lane="7" entrytime="00:01:27.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="288" swimtime="00:00:40.65" resultid="3002" heatid="5289" lane="6" />
                <RESULT eventid="1275" points="267" swimtime="00:03:11.01" resultid="3003" heatid="5340" lane="7" entrytime="00:03:06.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.79" />
                    <SPLIT distance="100" swimtime="00:01:32.69" />
                    <SPLIT distance="150" swimtime="00:02:22.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Ocanha" birthdate="2005-06-21" gender="M" nation="BRA" license="313769" swrid="5600231" athleteid="2885" externalid="313769" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1088" points="528" swimtime="00:01:10.35" resultid="2886" heatid="5087" lane="2" entrytime="00:01:11.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="580" swimtime="00:00:25.07" resultid="2887" heatid="5129" lane="4" entrytime="00:00:24.52" entrycourse="LCM" />
                <RESULT eventid="1297" points="609" swimtime="00:00:30.60" resultid="2888" heatid="5371" lane="2" entrytime="00:00:31.07" entrycourse="LCM" />
                <RESULT eventid="2320" swimtime="00:00:00.00" resultid="5961" entrytime="00:01:10.35" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jhon" lastname="Caleb Dos Santos" birthdate="2010-03-02" gender="M" nation="BRA" license="359020" swrid="5588574" athleteid="2930" externalid="359020">
              <RESULTS>
                <RESULT eventid="1151" points="520" swimtime="00:02:21.71" resultid="2931" heatid="5195" lane="4" entrytime="00:02:23.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                    <SPLIT distance="100" swimtime="00:01:05.86" />
                    <SPLIT distance="150" swimtime="00:01:49.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="521" swimtime="00:01:04.11" resultid="2932" heatid="5258" lane="4" entrytime="00:01:04.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="432" swimtime="00:05:20.69" resultid="2933" heatid="5277" lane="8" entrytime="00:05:16.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.73" />
                    <SPLIT distance="100" swimtime="00:01:10.45" />
                    <SPLIT distance="150" swimtime="00:01:50.99" />
                    <SPLIT distance="200" swimtime="00:02:31.22" />
                    <SPLIT distance="250" swimtime="00:03:19.43" />
                    <SPLIT distance="300" swimtime="00:04:07.27" />
                    <SPLIT distance="350" swimtime="00:04:44.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1293" points="435" swimtime="00:02:25.55" resultid="2934" heatid="5360" lane="8" entrytime="00:02:25.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                    <SPLIT distance="100" swimtime="00:01:10.10" />
                    <SPLIT distance="150" swimtime="00:01:48.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2359" swimtime="00:00:00.00" resultid="6449" entrytime="00:01:04.11" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Inacio Carneiro" birthdate="2009-09-09" gender="M" nation="BRA" license="408023" swrid="5723026" athleteid="3004" externalid="408023">
              <RESULTS>
                <RESULT eventid="1104" points="372" swimtime="00:00:29.07" resultid="3005" heatid="5122" lane="7" entrytime="00:00:29.17" entrycourse="LCM" />
                <RESULT eventid="1120" points="282" swimtime="00:02:35.49" resultid="3006" heatid="5153" lane="7" entrytime="00:02:36.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.05" />
                    <SPLIT distance="100" swimtime="00:01:14.55" />
                    <SPLIT distance="150" swimtime="00:01:56.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="313" swimtime="00:01:09.00" resultid="3007" heatid="5225" lane="7" entrytime="00:01:07.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="174" swimtime="00:00:42.12" resultid="3008" heatid="5284" lane="8" entrytime="00:00:44.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Faria Del Valle" birthdate="2009-08-28" gender="M" nation="BRA" license="376328" swrid="5600155" athleteid="2935" externalid="376328">
              <RESULTS>
                <RESULT eventid="1104" points="531" swimtime="00:00:25.81" resultid="2936" heatid="5126" lane="1" entrytime="00:00:25.37" entrycourse="LCM" />
                <RESULT eventid="1167" points="510" swimtime="00:00:58.62" resultid="2937" heatid="5229" lane="1" entrytime="00:00:57.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="444" swimtime="00:00:30.85" resultid="2938" heatid="5287" lane="8" entrytime="00:00:31.05" entrycourse="LCM" />
                <RESULT eventid="1267" points="500" swimtime="00:00:28.05" resultid="2939" heatid="5335" lane="3" entrytime="00:00:28.13" entrycourse="LCM" />
                <RESULT eventid="1297" points="478" swimtime="00:00:33.18" resultid="2940" heatid="5370" lane="8" entrytime="00:00:34.15" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Araujo Do Rego Barros" birthdate="2009-04-30" gender="M" nation="BRA" license="376325" swrid="5377739" athleteid="2920" externalid="376325">
              <RESULTS>
                <RESULT eventid="1104" points="363" swimtime="00:00:29.31" resultid="2921" heatid="5123" lane="1" entrytime="00:00:28.24" entrycourse="LCM" />
                <RESULT eventid="1135" points="368" swimtime="00:01:09.00" resultid="2922" heatid="5173" lane="5" entrytime="00:01:09.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="411" swimtime="00:01:02.99" resultid="2923" heatid="5225" lane="3" entrytime="00:01:04.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="378" swimtime="00:00:30.78" resultid="2924" heatid="5333" lane="2" entrytime="00:00:31.19" entrycourse="LCM" />
                <RESULT eventid="1293" points="350" swimtime="00:02:36.48" resultid="2925" heatid="5358" lane="4" entrytime="00:02:43.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:11.34" />
                    <SPLIT distance="150" swimtime="00:01:53.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="20" agetotalmax="-1" agetotalmin="-1" gender="M" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1241" points="492" swimtime="00:03:58.43" resultid="3027" heatid="5310" lane="7" entrytime="00:04:01.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.72" />
                    <SPLIT distance="100" swimtime="00:00:58.10" />
                    <SPLIT distance="150" swimtime="00:01:26.64" />
                    <SPLIT distance="200" swimtime="00:01:58.58" />
                    <SPLIT distance="250" swimtime="00:02:27.52" />
                    <SPLIT distance="300" swimtime="00:02:59.88" />
                    <SPLIT distance="350" swimtime="00:03:28.36" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2889" number="1" />
                    <RELAYPOSITION athleteid="2892" number="2" />
                    <RELAYPOSITION athleteid="2906" number="3" />
                    <RELAYPOSITION athleteid="2909" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1342" points="435" swimtime="00:04:32.85" resultid="3030" heatid="5390" lane="5" entrytime="00:04:29.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                    <SPLIT distance="100" swimtime="00:01:06.13" />
                    <SPLIT distance="150" swimtime="00:01:44.42" />
                    <SPLIT distance="200" swimtime="00:02:29.56" />
                    <SPLIT distance="250" swimtime="00:02:59.17" />
                    <SPLIT distance="300" swimtime="00:03:32.03" />
                    <SPLIT distance="350" swimtime="00:04:00.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2889" number="1" />
                    <RELAYPOSITION athleteid="2902" number="2" />
                    <RELAYPOSITION athleteid="2909" number="3" />
                    <RELAYPOSITION athleteid="2892" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1235" points="508" swimtime="00:03:55.87" resultid="3028" heatid="5307" lane="3" entrytime="00:03:58.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.63" />
                    <SPLIT distance="100" swimtime="00:00:58.10" />
                    <SPLIT distance="150" swimtime="00:01:27.19" />
                    <SPLIT distance="200" swimtime="00:01:58.25" />
                    <SPLIT distance="250" swimtime="00:02:27.61" />
                    <SPLIT distance="300" swimtime="00:03:00.72" />
                    <SPLIT distance="350" swimtime="00:03:26.13" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2935" number="1" />
                    <RELAYPOSITION athleteid="2914" number="2" />
                    <RELAYPOSITION athleteid="2975" number="3" />
                    <RELAYPOSITION athleteid="2880" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1336" points="469" swimtime="00:04:26.09" resultid="3032" heatid="5387" lane="6" entrytime="00:04:32.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.61" />
                    <SPLIT distance="100" swimtime="00:01:00.47" />
                    <SPLIT distance="150" swimtime="00:01:36.37" />
                    <SPLIT distance="200" swimtime="00:02:15.39" />
                    <SPLIT distance="250" swimtime="00:02:46.58" />
                    <SPLIT distance="300" swimtime="00:03:23.80" />
                    <SPLIT distance="350" swimtime="00:03:52.84" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2880" number="1" />
                    <RELAYPOSITION athleteid="2914" number="2" />
                    <RELAYPOSITION athleteid="2920" number="3" />
                    <RELAYPOSITION athleteid="2975" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1233" points="346" swimtime="00:04:28.03" resultid="3029" heatid="5306" lane="6" entrytime="00:04:20.49">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.94" />
                    <SPLIT distance="100" swimtime="00:01:09.60" />
                    <SPLIT distance="150" swimtime="00:01:40.38" />
                    <SPLIT distance="200" swimtime="00:02:15.04" />
                    <SPLIT distance="250" swimtime="00:02:46.16" />
                    <SPLIT distance="300" swimtime="00:03:20.49" />
                    <SPLIT distance="350" swimtime="00:03:52.20" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2980" number="1" />
                    <RELAYPOSITION athleteid="2951" number="2" />
                    <RELAYPOSITION athleteid="3015" number="3" />
                    <RELAYPOSITION athleteid="3009" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1334" points="363" swimtime="00:04:49.74" resultid="3031" heatid="5386" lane="6" entrytime="00:04:46.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="100" swimtime="00:01:17.40" />
                    <SPLIT distance="150" swimtime="00:01:56.84" />
                    <SPLIT distance="200" swimtime="00:02:41.01" />
                    <SPLIT distance="250" swimtime="00:03:10.26" />
                    <SPLIT distance="300" swimtime="00:03:43.71" />
                    <SPLIT distance="350" swimtime="00:04:15.14" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2951" number="1" />
                    <RELAYPOSITION athleteid="3009" number="2" />
                    <RELAYPOSITION athleteid="2930" number="3" />
                    <RELAYPOSITION athleteid="3015" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1225" points="457" swimtime="00:04:29.86" resultid="3025" heatid="5304" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:05.06" />
                    <SPLIT distance="150" swimtime="00:01:36.75" />
                    <SPLIT distance="200" swimtime="00:02:11.87" />
                    <SPLIT distance="250" swimtime="00:02:44.54" />
                    <SPLIT distance="300" swimtime="00:03:20.58" />
                    <SPLIT distance="350" swimtime="00:03:53.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2875" number="1" />
                    <RELAYPOSITION athleteid="2946" number="2" />
                    <RELAYPOSITION athleteid="2941" number="3" />
                    <RELAYPOSITION athleteid="2990" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1326" points="406" swimtime="00:05:10.92" resultid="3026" heatid="5384" lane="6" entrytime="00:05:11.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                    <SPLIT distance="100" swimtime="00:01:13.60" />
                    <SPLIT distance="150" swimtime="00:01:50.92" />
                    <SPLIT distance="200" swimtime="00:02:33.19" />
                    <SPLIT distance="250" swimtime="00:03:08.50" />
                    <SPLIT distance="350" swimtime="00:04:34.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2875" number="1" />
                    <RELAYPOSITION athleteid="2941" number="2" />
                    <RELAYPOSITION athleteid="2946" number="3" />
                    <RELAYPOSITION athleteid="2990" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="19" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1289" points="298" swimtime="00:05:25.69" resultid="3033" heatid="5355" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.32" />
                    <SPLIT distance="100" swimtime="00:01:32.58" />
                    <SPLIT distance="150" swimtime="00:02:23.51" />
                    <SPLIT distance="200" swimtime="00:03:17.71" />
                    <SPLIT distance="250" swimtime="00:03:48.50" />
                    <SPLIT distance="300" swimtime="00:04:27.01" />
                    <SPLIT distance="350" swimtime="00:04:55.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2968" number="1" />
                    <RELAYPOSITION athleteid="2962" number="2" />
                    <RELAYPOSITION athleteid="2897" number="3" />
                    <RELAYPOSITION athleteid="2885" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="ATN/CURITIBA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1285" points="541" swimtime="00:04:26.93" resultid="3034" heatid="5353" lane="3" entrytime="00:04:34.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.48" />
                    <SPLIT distance="100" swimtime="00:01:11.45" />
                    <SPLIT distance="150" swimtime="00:01:49.73" />
                    <SPLIT distance="200" swimtime="00:02:31.18" />
                    <SPLIT distance="250" swimtime="00:02:58.76" />
                    <SPLIT distance="300" swimtime="00:03:30.83" />
                    <SPLIT distance="350" swimtime="00:03:57.64" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2875" number="1" />
                    <RELAYPOSITION athleteid="2941" number="2" />
                    <RELAYPOSITION athleteid="2880" number="3" />
                    <RELAYPOSITION athleteid="2935" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="4096" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Lorenzo" lastname="Jacobsen Donati" birthdate="2011-07-14" gender="M" nation="BRA" license="391851" swrid="5615735" athleteid="4125" externalid="391851">
              <RESULTS>
                <RESULT eventid="1104" points="428" swimtime="00:00:27.74" resultid="4126" heatid="5120" lane="8" entrytime="00:00:27.51" entrycourse="LCM" />
                <RESULT eventid="1135" points="283" swimtime="00:01:15.28" resultid="4127" heatid="5169" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="365" swimtime="00:02:22.71" resultid="4128" heatid="5149" lane="2" entrytime="00:02:37.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="100" swimtime="00:01:07.31" />
                    <SPLIT distance="150" swimtime="00:01:45.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="435" swimtime="00:01:08.08" resultid="4129" heatid="5257" lane="4" entrytime="00:01:09.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="364" swimtime="00:02:36.63" resultid="4130" heatid="5346" lane="6" entrytime="00:02:32.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.18" />
                    <SPLIT distance="100" swimtime="00:01:16.82" />
                    <SPLIT distance="150" swimtime="00:01:57.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="281" swimtime="00:22:09.78" resultid="4131" heatid="5378" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.84" />
                    <SPLIT distance="100" swimtime="00:01:17.45" />
                    <SPLIT distance="150" swimtime="00:01:59.92" />
                    <SPLIT distance="200" swimtime="00:02:43.51" />
                    <SPLIT distance="250" swimtime="00:03:27.07" />
                    <SPLIT distance="300" swimtime="00:04:10.45" />
                    <SPLIT distance="350" swimtime="00:04:53.93" />
                    <SPLIT distance="400" swimtime="00:05:38.56" />
                    <SPLIT distance="450" swimtime="00:06:22.77" />
                    <SPLIT distance="500" swimtime="00:07:07.47" />
                    <SPLIT distance="550" swimtime="00:07:51.19" />
                    <SPLIT distance="600" swimtime="00:08:36.92" />
                    <SPLIT distance="650" swimtime="00:09:21.36" />
                    <SPLIT distance="700" swimtime="00:10:07.38" />
                    <SPLIT distance="750" swimtime="00:10:51.90" />
                    <SPLIT distance="800" swimtime="00:11:37.64" />
                    <SPLIT distance="850" swimtime="00:12:23.12" />
                    <SPLIT distance="900" swimtime="00:13:08.61" />
                    <SPLIT distance="950" swimtime="00:13:54.31" />
                    <SPLIT distance="1000" swimtime="00:14:39.54" />
                    <SPLIT distance="1050" swimtime="00:15:23.70" />
                    <SPLIT distance="1100" swimtime="00:16:09.49" />
                    <SPLIT distance="1150" swimtime="00:16:54.19" />
                    <SPLIT distance="1200" swimtime="00:17:40.24" />
                    <SPLIT distance="1250" swimtime="00:18:25.76" />
                    <SPLIT distance="1300" swimtime="00:19:11.49" />
                    <SPLIT distance="1350" swimtime="00:19:57.29" />
                    <SPLIT distance="1400" swimtime="00:20:43.28" />
                    <SPLIT distance="1450" swimtime="00:21:26.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rodrigo" lastname="Zanatta Duda" birthdate="2011-09-12" gender="M" nation="BRA" license="406917" swrid="5717307" athleteid="4198" externalid="406917">
              <RESULTS>
                <RESULT eventid="1151" points="233" swimtime="00:03:05.23" resultid="4199" heatid="5193" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                    <SPLIT distance="100" swimtime="00:01:24.80" />
                    <SPLIT distance="150" swimtime="00:02:20.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="287" swimtime="00:01:18.16" resultid="4200" heatid="5256" lane="7" entrytime="00:01:22.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="290" swimtime="00:00:35.55" resultid="4201" heatid="5284" lane="3" entrytime="00:00:37.54" entrycourse="LCM" />
                <RESULT eventid="1277" points="304" swimtime="00:02:46.44" resultid="4202" heatid="5344" lane="3" entrytime="00:03:06.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.32" />
                    <SPLIT distance="100" swimtime="00:01:23.08" />
                    <SPLIT distance="150" swimtime="00:02:05.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="203" swimtime="00:00:44.11" resultid="4203" heatid="5366" lane="6" entrytime="00:00:47.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Braga" birthdate="2010-05-07" gender="M" nation="BRA" license="378345" swrid="5343953" athleteid="4160" externalid="378345">
              <RESULTS>
                <RESULT eventid="1088" points="404" swimtime="00:01:16.93" resultid="4161" heatid="5082" lane="4" entrytime="00:01:13.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="166" swimtime="00:01:29.80" resultid="4162" heatid="5169" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="350" swimtime="00:01:06.49" resultid="4163" heatid="5217" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="217" swimtime="00:00:39.16" resultid="4164" heatid="5283" lane="4" entrytime="00:00:44.45" entrycourse="LCM" />
                <RESULT eventid="1251" points="401" swimtime="00:02:50.08" resultid="4165" heatid="5319" lane="2" entrytime="00:02:43.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                    <SPLIT distance="100" swimtime="00:01:20.80" />
                    <SPLIT distance="150" swimtime="00:02:05.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="428" swimtime="00:00:34.42" resultid="4166" heatid="5368" lane="3" entrytime="00:00:35.86" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Kenji Yamaguchi" birthdate="2011-08-25" gender="M" nation="BRA" license="385708" swrid="5603862" athleteid="4132" externalid="385708">
              <RESULTS>
                <RESULT eventid="1088" points="244" swimtime="00:01:30.90" resultid="4133" heatid="5079" lane="5" entrytime="00:01:33.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="271" swimtime="00:01:16.37" resultid="4134" heatid="5170" lane="7" entrytime="00:01:23.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="285" swimtime="00:06:08.15" resultid="4135" heatid="5275" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.29" />
                    <SPLIT distance="100" swimtime="00:01:17.02" />
                    <SPLIT distance="150" swimtime="00:02:07.45" />
                    <SPLIT distance="200" swimtime="00:02:55.65" />
                    <SPLIT distance="250" swimtime="00:03:47.37" />
                    <SPLIT distance="300" swimtime="00:04:37.88" />
                    <SPLIT distance="350" swimtime="00:05:24.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="253" swimtime="00:00:35.21" resultid="4136" heatid="5331" lane="5" entrytime="00:00:35.41" entrycourse="LCM" />
                <RESULT eventid="1251" points="251" swimtime="00:03:18.66" resultid="4137" heatid="5316" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.56" />
                    <SPLIT distance="100" swimtime="00:01:35.10" />
                    <SPLIT distance="150" swimtime="00:02:27.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1293" points="252" swimtime="00:02:54.68" resultid="4138" heatid="5357" lane="5" entrytime="00:03:18.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                    <SPLIT distance="100" swimtime="00:01:20.17" />
                    <SPLIT distance="150" swimtime="00:02:07.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Sales" birthdate="2011-02-28" gender="F" nation="BRA" license="374103" swrid="5616410" athleteid="4167" externalid="374103">
              <RESULTS>
                <RESULT eventid="1080" points="359" swimtime="00:01:30.17" resultid="4168" heatid="5066" lane="3" entrytime="00:01:29.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="507" swimtime="00:00:29.59" resultid="4169" heatid="5100" lane="3" entrytime="00:00:29.26" entrycourse="LCM" />
                <RESULT eventid="1128" points="443" swimtime="00:01:12.73" resultid="4170" heatid="5160" lane="2" entrytime="00:01:16.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="375" swimtime="00:02:54.85" resultid="4171" heatid="5186" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:24.07" />
                    <SPLIT distance="150" swimtime="00:02:13.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="312" swimtime="00:01:24.49" resultid="4172" heatid="5241" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="462" swimtime="00:01:06.87" resultid="4173" heatid="5202" lane="4" entrytime="00:01:11.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2328" points="367" swimtime="00:01:17.48" resultid="6001" heatid="6418" lane="2" entrytime="00:01:12.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eloah" lastname="Juvedi Trindade" birthdate="2011-03-05" gender="F" nation="BRA" license="396829" swrid="5641768" athleteid="4174" externalid="396829">
              <RESULTS>
                <RESULT eventid="1080" points="272" swimtime="00:01:38.92" resultid="4175" heatid="5065" lane="6" entrytime="00:01:50.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="319" swimtime="00:00:34.55" resultid="4176" heatid="5096" lane="2" entrytime="00:00:38.02" entrycourse="LCM" />
                <RESULT eventid="1143" points="235" swimtime="00:03:24.25" resultid="4177" heatid="5186" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.14" />
                    <SPLIT distance="100" swimtime="00:01:36.17" />
                    <SPLIT distance="150" swimtime="00:02:36.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="239" swimtime="00:01:32.33" resultid="4178" heatid="5241" lane="2" />
                <RESULT eventid="1215" points="258" swimtime="00:00:42.18" resultid="4179" heatid="5291" lane="2" entrytime="00:00:47.07" entrycourse="LCM" />
                <RESULT eventid="1259" points="182" swimtime="00:00:43.07" resultid="4180" heatid="5321" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benicio" lastname="Garcia" birthdate="2011-09-09" gender="M" nation="BRA" license="378347" swrid="5603842" athleteid="4097" externalid="378347">
              <RESULTS>
                <RESULT eventid="1072" points="227" swimtime="00:06:00.52" resultid="4098" heatid="5056" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                    <SPLIT distance="100" swimtime="00:01:19.80" />
                    <SPLIT distance="150" swimtime="00:02:06.20" />
                    <SPLIT distance="200" swimtime="00:02:53.11" />
                    <SPLIT distance="250" swimtime="00:03:41.89" />
                    <SPLIT distance="300" swimtime="00:04:28.23" />
                    <SPLIT distance="350" swimtime="00:05:15.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="272" swimtime="00:00:32.24" resultid="4099" heatid="5115" lane="4" entrytime="00:00:34.48" entrycourse="LCM" />
                <RESULT eventid="1135" points="147" swimtime="00:01:33.63" resultid="4100" heatid="5169" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="285" swimtime="00:01:18.34" resultid="4101" heatid="5256" lane="3" entrytime="00:01:19.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="256" swimtime="00:11:51.23" resultid="4102" heatid="5297" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.64" />
                    <SPLIT distance="100" swimtime="00:01:21.73" />
                    <SPLIT distance="150" swimtime="00:02:06.87" />
                    <SPLIT distance="200" swimtime="00:02:52.11" />
                    <SPLIT distance="250" swimtime="00:03:37.68" />
                    <SPLIT distance="300" swimtime="00:04:23.60" />
                    <SPLIT distance="350" swimtime="00:05:09.79" />
                    <SPLIT distance="400" swimtime="00:05:55.33" />
                    <SPLIT distance="450" swimtime="00:06:40.66" />
                    <SPLIT distance="500" swimtime="00:07:26.35" />
                    <SPLIT distance="550" swimtime="00:08:11.30" />
                    <SPLIT distance="600" swimtime="00:08:56.74" />
                    <SPLIT distance="650" swimtime="00:09:41.97" />
                    <SPLIT distance="700" swimtime="00:10:26.80" />
                    <SPLIT distance="750" swimtime="00:11:09.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="244" swimtime="00:02:58.87" resultid="4103" heatid="5344" lane="5" entrytime="00:03:01.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.84" />
                    <SPLIT distance="100" swimtime="00:01:23.43" />
                    <SPLIT distance="150" swimtime="00:02:12.38" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theodoro" lastname="Marques Serra" birthdate="2009-11-24" gender="M" nation="BRA" license="370661" swrid="5603870" athleteid="4118" externalid="370661">
              <RESULTS>
                <RESULT eventid="1104" points="407" swimtime="00:00:28.20" resultid="4119" heatid="5121" lane="5" entrytime="00:00:30.33" entrycourse="LCM" />
                <RESULT eventid="1120" points="400" swimtime="00:02:18.33" resultid="4120" heatid="5154" lane="3" entrytime="00:02:17.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.30" />
                    <SPLIT distance="100" swimtime="00:01:04.93" />
                    <SPLIT distance="150" swimtime="00:01:41.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="366" swimtime="00:02:39.28" resultid="4121" heatid="5196" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                    <SPLIT distance="100" swimtime="00:01:14.33" />
                    <SPLIT distance="150" swimtime="00:02:03.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="406" swimtime="00:01:09.68" resultid="4122" heatid="5260" lane="2" entrytime="00:01:10.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="387" swimtime="00:10:20.26" resultid="4123" heatid="5296" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.44" />
                    <SPLIT distance="100" swimtime="00:01:11.81" />
                    <SPLIT distance="150" swimtime="00:01:51.63" />
                    <SPLIT distance="200" swimtime="00:02:30.95" />
                    <SPLIT distance="250" swimtime="00:03:10.89" />
                    <SPLIT distance="300" swimtime="00:03:50.56" />
                    <SPLIT distance="350" swimtime="00:04:30.89" />
                    <SPLIT distance="400" swimtime="00:05:09.95" />
                    <SPLIT distance="450" swimtime="00:05:50.27" />
                    <SPLIT distance="500" swimtime="00:06:29.55" />
                    <SPLIT distance="550" swimtime="00:07:09.23" />
                    <SPLIT distance="600" swimtime="00:07:48.19" />
                    <SPLIT distance="650" swimtime="00:08:27.52" />
                    <SPLIT distance="700" swimtime="00:09:05.93" />
                    <SPLIT distance="750" swimtime="00:09:43.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="412" swimtime="00:19:29.99" resultid="4124" heatid="5378" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="100" swimtime="00:01:10.65" />
                    <SPLIT distance="150" swimtime="00:01:50.24" />
                    <SPLIT distance="200" swimtime="00:02:29.87" />
                    <SPLIT distance="250" swimtime="00:03:10.16" />
                    <SPLIT distance="300" swimtime="00:03:49.72" />
                    <SPLIT distance="350" swimtime="00:04:29.95" />
                    <SPLIT distance="400" swimtime="00:05:10.14" />
                    <SPLIT distance="450" swimtime="00:05:50.32" />
                    <SPLIT distance="500" swimtime="00:06:30.33" />
                    <SPLIT distance="550" swimtime="00:07:10.80" />
                    <SPLIT distance="600" swimtime="00:07:50.65" />
                    <SPLIT distance="650" swimtime="00:08:30.49" />
                    <SPLIT distance="700" swimtime="00:09:09.93" />
                    <SPLIT distance="750" swimtime="00:09:49.83" />
                    <SPLIT distance="800" swimtime="00:10:29.51" />
                    <SPLIT distance="850" swimtime="00:11:09.39" />
                    <SPLIT distance="900" swimtime="00:11:48.86" />
                    <SPLIT distance="950" swimtime="00:12:28.28" />
                    <SPLIT distance="1000" swimtime="00:13:07.55" />
                    <SPLIT distance="1050" swimtime="00:13:46.75" />
                    <SPLIT distance="1100" swimtime="00:14:25.90" />
                    <SPLIT distance="1150" swimtime="00:15:04.25" />
                    <SPLIT distance="1200" swimtime="00:15:42.88" />
                    <SPLIT distance="1250" swimtime="00:16:21.82" />
                    <SPLIT distance="1300" swimtime="00:17:00.45" />
                    <SPLIT distance="1350" swimtime="00:17:38.50" />
                    <SPLIT distance="1400" swimtime="00:18:16.52" />
                    <SPLIT distance="1450" swimtime="00:18:53.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Traci Rodrigues" birthdate="2011-03-06" gender="M" nation="BRA" license="406927" swrid="5718893" athleteid="4104" externalid="406927">
              <RESULTS>
                <RESULT eventid="1088" points="174" swimtime="00:01:41.74" resultid="4105" heatid="5079" lane="1" entrytime="00:01:50.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="231" swimtime="00:00:34.06" resultid="4106" heatid="5115" lane="2" entrytime="00:00:36.29" entrycourse="LCM" />
                <RESULT eventid="1120" points="181" swimtime="00:03:00.23" resultid="4107" heatid="5148" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.53" />
                    <SPLIT distance="100" swimtime="00:01:21.75" />
                    <SPLIT distance="150" swimtime="00:02:11.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="237" swimtime="00:01:15.66" resultid="4108" heatid="5218" lane="2" entrytime="00:01:23.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="155" swimtime="00:00:43.78" resultid="4109" heatid="5283" lane="3" entrytime="00:00:46.27" entrycourse="LCM" />
                <RESULT eventid="1297" points="185" swimtime="00:00:45.47" resultid="4110" heatid="5366" lane="3" entrytime="00:00:46.94" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Jennifer" lastname="De Abreu" birthdate="2009-11-07" gender="F" nation="BRA" license="356212" swrid="5600144" athleteid="4153" externalid="356212">
              <RESULTS>
                <RESULT eventid="1096" points="477" swimtime="00:00:30.21" resultid="4154" heatid="5104" lane="1" entrytime="00:00:29.54" entrycourse="LCM" />
                <RESULT eventid="1112" points="531" swimtime="00:02:19.28" resultid="4155" heatid="5144" lane="2" entrytime="00:02:21.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.84" />
                    <SPLIT distance="100" swimtime="00:01:08.31" />
                    <SPLIT distance="150" swimtime="00:01:43.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="426" swimtime="00:02:47.56" resultid="4156" heatid="5190" lane="6" entrytime="00:02:42.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                    <SPLIT distance="100" swimtime="00:01:20.17" />
                    <SPLIT distance="150" swimtime="00:02:12.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="517" swimtime="00:01:04.39" resultid="4157" heatid="5208" lane="1" entrytime="00:01:03.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="392" swimtime="00:00:36.67" resultid="4158" heatid="5290" lane="7" />
                <RESULT eventid="1259" points="463" swimtime="00:00:31.57" resultid="4159" heatid="5325" lane="7" entrytime="00:00:34.95" entrycourse="LCM" />
                <RESULT eventid="2343" swimtime="00:00:00.00" resultid="6110" entrytime="00:01:04.39" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Ferreira Rais" birthdate="2007-07-04" gender="M" nation="BRA" license="398656" swrid="5697227" athleteid="4186" externalid="398656">
              <RESULTS>
                <RESULT eventid="1104" points="431" swimtime="00:00:27.68" resultid="4187" heatid="5127" lane="4" entrytime="00:00:28.28" entrycourse="LCM" />
                <RESULT eventid="1135" points="251" swimtime="00:01:18.36" resultid="4188" heatid="5176" lane="6" entrytime="00:01:22.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="373" swimtime="00:01:05.09" resultid="4189" heatid="5231" lane="2" entrytime="00:01:06.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="290" swimtime="00:00:33.64" resultid="4190" heatid="5332" lane="5" entrytime="00:00:31.81" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Pazinato" birthdate="2011-01-05" gender="M" nation="BRA" license="368149" swrid="5603889" athleteid="4139" externalid="368149">
              <RESULTS>
                <RESULT eventid="1072" points="328" swimtime="00:05:18.95" resultid="4140" heatid="5057" lane="7" entrytime="00:05:47.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:10.91" />
                    <SPLIT distance="150" swimtime="00:01:51.90" />
                    <SPLIT distance="200" swimtime="00:02:34.02" />
                    <SPLIT distance="250" swimtime="00:03:16.39" />
                    <SPLIT distance="300" swimtime="00:03:59.22" />
                    <SPLIT distance="350" swimtime="00:04:41.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="343" swimtime="00:00:29.85" resultid="4141" heatid="5117" lane="8" entrytime="00:00:30.94" entrycourse="LCM" />
                <RESULT eventid="1120" points="317" swimtime="00:02:29.44" resultid="4142" heatid="5149" lane="5" entrytime="00:02:34.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.25" />
                    <SPLIT distance="100" swimtime="00:01:10.46" />
                    <SPLIT distance="150" swimtime="00:01:50.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="306" swimtime="00:01:16.49" resultid="4143" heatid="5256" lane="2" entrytime="00:01:20.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="383" swimtime="00:01:04.50" resultid="4144" heatid="5220" lane="3" entrytime="00:01:07.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="293" swimtime="00:02:48.50" resultid="4145" heatid="5344" lane="4" entrytime="00:02:57.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.87" />
                    <SPLIT distance="100" swimtime="00:01:19.27" />
                    <SPLIT distance="150" swimtime="00:02:04.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Silveira De Almeida" birthdate="2008-07-08" gender="M" nation="BRA" license="368152" swrid="5603912" athleteid="4146" externalid="368152">
              <RESULTS>
                <RESULT eventid="1088" points="349" swimtime="00:01:20.78" resultid="4147" heatid="5083" lane="2" entrytime="00:01:33.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="439" swimtime="00:00:27.51" resultid="4148" heatid="5123" lane="4" entrytime="00:00:27.49" entrycourse="LCM" />
                <RESULT eventid="1135" points="477" swimtime="00:01:03.25" resultid="4149" heatid="5175" lane="2" entrytime="00:01:01.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="357" swimtime="00:01:12.72" resultid="4150" heatid="5259" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="490" swimtime="00:00:28.23" resultid="4151" heatid="5336" lane="1" entrytime="00:00:27.76" entrycourse="LCM" />
                <RESULT eventid="1297" points="380" swimtime="00:00:35.81" resultid="4152" heatid="5363" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Ribeiro Melo" birthdate="2011-07-01" gender="F" nation="BRA" license="390923" swrid="5602577" athleteid="4111" externalid="390923">
              <RESULTS>
                <RESULT eventid="1064" points="368" swimtime="00:05:28.28" resultid="4112" heatid="5049" lane="2" entrytime="00:05:33.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.69" />
                    <SPLIT distance="100" swimtime="00:01:16.71" />
                    <SPLIT distance="150" swimtime="00:01:59.56" />
                    <SPLIT distance="200" swimtime="00:02:41.73" />
                    <SPLIT distance="250" swimtime="00:03:25.30" />
                    <SPLIT distance="300" swimtime="00:04:07.67" />
                    <SPLIT distance="350" swimtime="00:04:50.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="443" swimtime="00:00:30.97" resultid="4113" heatid="5100" lane="1" entrytime="00:00:30.29" entrycourse="LCM" />
                <RESULT eventid="1112" points="430" swimtime="00:02:29.45" resultid="4114" heatid="5139" lane="7" entrytime="00:02:34.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:11.64" />
                    <SPLIT distance="150" swimtime="00:01:50.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="435" swimtime="00:01:08.22" resultid="4115" heatid="5203" lane="5" entrytime="00:01:09.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="201" swimtime="00:00:41.68" resultid="4116" heatid="5322" lane="2" />
                <RESULT eventid="1243" points="272" swimtime="00:03:32.07" resultid="4117" heatid="5311" lane="1" entrytime="00:03:33.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.64" />
                    <SPLIT distance="100" swimtime="00:01:39.27" />
                    <SPLIT distance="150" swimtime="00:02:36.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Camillo Sabim" birthdate="2010-08-02" gender="F" nation="BRA" license="406931" swrid="5723021" athleteid="4211" externalid="406931">
              <RESULTS>
                <RESULT eventid="1080" points="310" swimtime="00:01:34.67" resultid="4212" heatid="5065" lane="4" entrytime="00:01:37.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="335" swimtime="00:00:33.99" resultid="4213" heatid="5097" lane="1" entrytime="00:00:35.39" entrycourse="LCM" />
                <RESULT eventid="1159" points="358" swimtime="00:01:12.79" resultid="4214" heatid="5201" lane="2" entrytime="00:01:22.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="345" swimtime="00:00:41.57" resultid="4215" heatid="5374" lane="4" entrytime="00:00:43.56" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Guilherme Ballatka" birthdate="2007-06-24" gender="M" nation="BRA" license="398616" swrid="5697228" athleteid="4181" externalid="398616">
              <RESULTS>
                <RESULT eventid="1088" points="304" swimtime="00:01:24.52" resultid="4182" heatid="5086" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="478" swimtime="00:00:26.73" resultid="4183" heatid="5128" lane="7" entrytime="00:00:27.41" entrycourse="LCM" />
                <RESULT eventid="1182" points="447" swimtime="00:01:07.46" resultid="4184" heatid="5262" lane="3" entrytime="00:01:10.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="442" swimtime="00:01:01.48" resultid="4185" heatid="5231" lane="3" entrytime="00:01:02.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Bilemjian Leszczynski" birthdate="2011-08-06" gender="M" nation="BRA" license="406925" swrid="5587326" athleteid="4204" externalid="406925">
              <RESULTS>
                <RESULT eventid="1088" points="154" swimtime="00:01:46.01" resultid="4205" heatid="5078" lane="4" />
                <RESULT eventid="1104" points="225" swimtime="00:00:34.36" resultid="4206" heatid="5115" lane="1" />
                <RESULT eventid="1135" points="114" swimtime="00:01:41.81" resultid="4207" heatid="5169" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="216" swimtime="00:01:18.10" resultid="4208" heatid="5217" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="149" swimtime="00:00:41.93" resultid="4209" heatid="5328" lane="3" />
                <RESULT eventid="1297" points="158" swimtime="00:00:47.91" resultid="4210" heatid="5365" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Aline" lastname="Hirano" birthdate="2007-11-13" gender="F" nation="BRA" license="358898" swrid="5622283" athleteid="4191" externalid="358898">
              <RESULTS>
                <RESULT eventid="1064" points="422" swimtime="00:05:13.66" resultid="4192" heatid="5055" lane="7" entrytime="00:05:13.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.61" />
                    <SPLIT distance="100" swimtime="00:01:10.21" />
                    <SPLIT distance="150" swimtime="00:01:48.23" />
                    <SPLIT distance="200" swimtime="00:02:29.06" />
                    <SPLIT distance="250" swimtime="00:03:11.41" />
                    <SPLIT distance="300" swimtime="00:03:54.66" />
                    <SPLIT distance="350" swimtime="00:04:34.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="392" swimtime="00:02:52.31" resultid="4193" heatid="5191" lane="3" entrytime="00:02:54.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                    <SPLIT distance="100" swimtime="00:01:21.85" />
                    <SPLIT distance="150" swimtime="00:02:16.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="397" swimtime="00:01:17.98" resultid="4194" heatid="5248" lane="6" entrytime="00:01:18.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="394" swimtime="00:11:00.83" resultid="4195" heatid="5273" lane="2" entrytime="00:10:54.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                    <SPLIT distance="100" swimtime="00:01:13.16" />
                    <SPLIT distance="150" swimtime="00:01:52.71" />
                    <SPLIT distance="200" swimtime="00:02:33.40" />
                    <SPLIT distance="250" swimtime="00:03:15.38" />
                    <SPLIT distance="300" swimtime="00:03:57.66" />
                    <SPLIT distance="350" swimtime="00:04:39.92" />
                    <SPLIT distance="400" swimtime="00:05:22.70" />
                    <SPLIT distance="450" swimtime="00:06:05.60" />
                    <SPLIT distance="500" swimtime="00:06:48.62" />
                    <SPLIT distance="550" swimtime="00:07:31.86" />
                    <SPLIT distance="600" swimtime="00:08:14.60" />
                    <SPLIT distance="650" swimtime="00:08:57.78" />
                    <SPLIT distance="700" swimtime="00:09:40.47" />
                    <SPLIT distance="750" swimtime="00:10:21.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="374" swimtime="00:06:08.90" resultid="4196" heatid="5278" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                    <SPLIT distance="100" swimtime="00:01:30.72" />
                    <SPLIT distance="150" swimtime="00:02:17.01" />
                    <SPLIT distance="200" swimtime="00:03:02.28" />
                    <SPLIT distance="250" swimtime="00:03:56.75" />
                    <SPLIT distance="300" swimtime="00:04:50.64" />
                    <SPLIT distance="350" swimtime="00:05:30.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1279" points="385" swimtime="00:21:04.54" resultid="4197" heatid="5349" lane="5" entrytime="00:20:52.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.01" />
                    <SPLIT distance="100" swimtime="00:01:12.82" />
                    <SPLIT distance="150" swimtime="00:01:52.51" />
                    <SPLIT distance="200" swimtime="00:02:33.14" />
                    <SPLIT distance="250" swimtime="00:03:14.11" />
                    <SPLIT distance="300" swimtime="00:03:55.90" />
                    <SPLIT distance="350" swimtime="00:04:37.57" />
                    <SPLIT distance="400" swimtime="00:05:19.66" />
                    <SPLIT distance="450" swimtime="00:06:02.55" />
                    <SPLIT distance="500" swimtime="00:06:46.58" />
                    <SPLIT distance="550" swimtime="00:07:26.45" />
                    <SPLIT distance="600" swimtime="00:08:08.42" />
                    <SPLIT distance="650" swimtime="00:08:51.63" />
                    <SPLIT distance="700" swimtime="00:09:35.01" />
                    <SPLIT distance="750" swimtime="00:10:18.05" />
                    <SPLIT distance="800" swimtime="00:11:01.15" />
                    <SPLIT distance="850" swimtime="00:11:44.71" />
                    <SPLIT distance="900" swimtime="00:12:28.76" />
                    <SPLIT distance="950" swimtime="00:13:12.85" />
                    <SPLIT distance="1000" swimtime="00:13:57.71" />
                    <SPLIT distance="1050" swimtime="00:14:38.47" />
                    <SPLIT distance="1100" swimtime="00:15:20.78" />
                    <SPLIT distance="1150" swimtime="00:16:03.56" />
                    <SPLIT distance="1200" swimtime="00:16:47.12" />
                    <SPLIT distance="1250" swimtime="00:17:30.37" />
                    <SPLIT distance="1300" swimtime="00:18:14.07" />
                    <SPLIT distance="1350" swimtime="00:18:57.87" />
                    <SPLIT distance="1400" swimtime="00:19:41.47" />
                    <SPLIT distance="1450" swimtime="00:20:23.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="263" nation="BRA" region="PR" clubid="3456" swrid="75436" name="Clube Curitibano" shortname="Curitibano">
          <ATHLETES>
            <ATHLETE firstname="Vinícius" lastname="Oliveira Cruz" birthdate="2005-07-02" gender="M" nation="BRA" license="298495" swrid="5653299" athleteid="3958" externalid="298495" level="ADTRISC">
              <RESULTS>
                <RESULT eventid="1072" points="691" swimtime="00:04:08.83" resultid="3959" heatid="5064" lane="4" entrytime="00:04:03.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.65" />
                    <SPLIT distance="100" swimtime="00:00:59.26" />
                    <SPLIT distance="150" swimtime="00:01:30.39" />
                    <SPLIT distance="200" swimtime="00:02:01.69" />
                    <SPLIT distance="250" swimtime="00:02:33.40" />
                    <SPLIT distance="300" swimtime="00:03:05.44" />
                    <SPLIT distance="350" swimtime="00:03:37.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="619" swimtime="00:00:24.53" resultid="3960" heatid="5130" lane="3" entrytime="00:00:23.64" entrycourse="LCM" />
                <RESULT eventid="1120" points="732" swimtime="00:01:53.16" resultid="3961" heatid="5158" lane="4" entrytime="00:01:50.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.24" />
                    <SPLIT distance="100" swimtime="00:00:56.79" />
                    <SPLIT distance="150" swimtime="00:01:25.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="722" swimtime="00:00:52.22" resultid="3962" heatid="5233" lane="3" entrytime="00:00:51.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="646" swimtime="00:08:42.78" resultid="3963" heatid="5296" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.36" />
                    <SPLIT distance="100" swimtime="00:00:59.86" />
                    <SPLIT distance="150" swimtime="00:01:31.84" />
                    <SPLIT distance="200" swimtime="00:02:03.72" />
                    <SPLIT distance="250" swimtime="00:02:36.16" />
                    <SPLIT distance="300" swimtime="00:03:08.70" />
                    <SPLIT distance="350" swimtime="00:03:41.67" />
                    <SPLIT distance="400" swimtime="00:04:14.88" />
                    <SPLIT distance="450" swimtime="00:04:48.56" />
                    <SPLIT distance="500" swimtime="00:05:22.19" />
                    <SPLIT distance="550" swimtime="00:05:55.87" />
                    <SPLIT distance="600" swimtime="00:06:29.75" />
                    <SPLIT distance="650" swimtime="00:07:03.55" />
                    <SPLIT distance="700" swimtime="00:07:37.15" />
                    <SPLIT distance="750" swimtime="00:08:10.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2383" points="616" swimtime="00:00:24.57" resultid="5985" heatid="6425" lane="1" entrytime="00:00:24.53" />
                <RESULT eventid="2351" points="714" swimtime="00:00:52.42" resultid="6118" heatid="6422" lane="3" entrytime="00:00:52.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorena" lastname="Mascarenhas" birthdate="2011-08-31" gender="F" nation="BRA" license="370581" swrid="5602558" athleteid="3838" externalid="370581">
              <RESULTS>
                <RESULT eventid="1096" points="398" swimtime="00:00:32.09" resultid="3839" heatid="5098" lane="7" entrytime="00:00:32.98" entrycourse="LCM" />
                <RESULT eventid="1112" points="381" swimtime="00:02:35.60" resultid="3840" heatid="5140" lane="7" entrytime="00:02:28.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.15" />
                    <SPLIT distance="100" swimtime="00:01:14.44" />
                    <SPLIT distance="150" swimtime="00:01:54.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="401" swimtime="00:02:50.94" resultid="3841" heatid="5187" lane="4" entrytime="00:02:49.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.63" />
                    <SPLIT distance="100" swimtime="00:01:22.35" />
                    <SPLIT distance="150" swimtime="00:02:14.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="383" swimtime="00:01:18.91" resultid="3842" heatid="5244" lane="1" entrytime="00:01:16.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="405" swimtime="00:01:09.86" resultid="3843" heatid="5204" lane="7" entrytime="00:01:08.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1275" points="385" swimtime="00:02:49.15" resultid="3844" heatid="5342" lane="4" entrytime="00:02:45.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.07" />
                    <SPLIT distance="100" swimtime="00:01:22.35" />
                    <SPLIT distance="150" swimtime="00:02:06.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Saboia" birthdate="2009-01-25" gender="M" nation="BRA" license="342252" swrid="5600253" athleteid="3602" externalid="342252">
              <RESULTS>
                <RESULT eventid="1088" points="491" swimtime="00:01:12.06" resultid="3603" heatid="5085" lane="8" entrytime="00:01:13.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="442" swimtime="00:02:29.65" resultid="3604" heatid="5197" lane="7" entrytime="00:02:32.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.97" />
                    <SPLIT distance="100" swimtime="00:01:13.38" />
                    <SPLIT distance="150" swimtime="00:01:55.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="481" swimtime="00:02:40.13" resultid="3605" heatid="5319" lane="3" entrytime="00:02:40.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.40" />
                    <SPLIT distance="100" swimtime="00:01:16.89" />
                    <SPLIT distance="150" swimtime="00:01:58.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="456" swimtime="00:00:33.69" resultid="3606" heatid="5370" lane="1" entrytime="00:00:33.71" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Clara Fernandes Pereira" birthdate="2009-11-19" gender="F" nation="BRA" license="344340" swrid="5600137" athleteid="3461" externalid="344340">
              <RESULTS>
                <RESULT eventid="1064" points="550" swimtime="00:04:47.20" resultid="3462" heatid="5053" lane="3" entrytime="00:04:47.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                    <SPLIT distance="100" swimtime="00:01:07.98" />
                    <SPLIT distance="150" swimtime="00:01:43.71" />
                    <SPLIT distance="200" swimtime="00:02:19.80" />
                    <SPLIT distance="250" swimtime="00:02:56.01" />
                    <SPLIT distance="300" swimtime="00:03:32.33" />
                    <SPLIT distance="350" swimtime="00:04:09.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="499" swimtime="00:02:38.92" resultid="3463" heatid="5190" lane="7" entrytime="00:02:43.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.75" />
                    <SPLIT distance="100" swimtime="00:01:17.00" />
                    <SPLIT distance="150" swimtime="00:02:04.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="533" swimtime="00:09:57.75" resultid="3464" heatid="5272" lane="5" entrytime="00:09:48.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                    <SPLIT distance="100" swimtime="00:01:10.00" />
                    <SPLIT distance="150" swimtime="00:01:48.37" />
                    <SPLIT distance="200" swimtime="00:02:26.54" />
                    <SPLIT distance="250" swimtime="00:03:04.46" />
                    <SPLIT distance="300" swimtime="00:03:42.35" />
                    <SPLIT distance="350" swimtime="00:04:20.77" />
                    <SPLIT distance="400" swimtime="00:04:58.54" />
                    <SPLIT distance="450" swimtime="00:05:36.98" />
                    <SPLIT distance="500" swimtime="00:06:14.67" />
                    <SPLIT distance="550" swimtime="00:06:52.53" />
                    <SPLIT distance="600" swimtime="00:07:29.96" />
                    <SPLIT distance="650" swimtime="00:08:07.78" />
                    <SPLIT distance="700" swimtime="00:08:45.00" />
                    <SPLIT distance="750" swimtime="00:09:22.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="3465" heatid="5280" lane="7" entrytime="00:05:42.05" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fernandes" birthdate="2010-03-13" gender="M" nation="BRA" license="339266" swrid="5588695" athleteid="3896" externalid="339266">
              <RESULTS>
                <RESULT eventid="1104" points="510" swimtime="00:00:26.17" resultid="3897" heatid="5120" lane="3" entrytime="00:00:26.65" entrycourse="LCM" />
                <RESULT eventid="1120" points="518" swimtime="00:02:06.93" resultid="3898" heatid="5152" lane="6" entrytime="00:02:10.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.43" />
                    <SPLIT distance="100" swimtime="00:01:02.05" />
                    <SPLIT distance="150" swimtime="00:01:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="432" swimtime="00:01:08.21" resultid="3899" heatid="5258" lane="1" entrytime="00:01:08.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="539" swimtime="00:00:57.58" resultid="3900" heatid="5223" lane="2" entrytime="00:00:58.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="427" swimtime="00:00:31.27" resultid="3901" heatid="5282" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Martynychen" birthdate="2011-12-19" gender="M" nation="BRA" license="366893" swrid="5602557" athleteid="3740" externalid="366893">
              <RESULTS>
                <RESULT eventid="1072" points="421" swimtime="00:04:53.62" resultid="3741" heatid="5058" lane="4" entrytime="00:04:54.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:08.59" />
                    <SPLIT distance="150" swimtime="00:01:45.69" />
                    <SPLIT distance="200" swimtime="00:02:23.42" />
                    <SPLIT distance="250" swimtime="00:03:01.15" />
                    <SPLIT distance="300" swimtime="00:03:39.44" />
                    <SPLIT distance="350" swimtime="00:04:17.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="367" swimtime="00:02:22.34" resultid="3742" heatid="5150" lane="2" entrytime="00:02:27.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="100" swimtime="00:01:08.59" />
                    <SPLIT distance="150" swimtime="00:01:45.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Bussmann" birthdate="2007-01-16" gender="F" nation="BRA" license="313781" swrid="5579983" athleteid="3512" externalid="313781">
              <RESULTS>
                <RESULT eventid="1080" points="558" swimtime="00:01:17.89" resultid="3513" heatid="5070" lane="5" entrytime="00:01:14.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" points="519" swimtime="00:04:52.71" resultid="3514" heatid="5054" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:11.00" />
                    <SPLIT distance="150" swimtime="00:01:48.69" />
                    <SPLIT distance="200" swimtime="00:02:26.49" />
                    <SPLIT distance="250" swimtime="00:03:03.57" />
                    <SPLIT distance="300" swimtime="00:03:40.49" />
                    <SPLIT distance="350" swimtime="00:04:17.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="544" swimtime="00:02:18.18" resultid="3515" heatid="5146" lane="2" entrytime="00:02:17.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                    <SPLIT distance="100" swimtime="00:01:06.95" />
                    <SPLIT distance="150" swimtime="00:01:42.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Fontolan Gomes" birthdate="2008-05-01" gender="M" nation="BRA" license="307667" swrid="5600166" athleteid="3563" externalid="307667">
              <RESULTS>
                <RESULT eventid="1104" points="446" swimtime="00:00:27.36" resultid="3564" heatid="5123" lane="6" entrytime="00:00:27.86" entrycourse="LCM" />
                <RESULT eventid="1135" points="388" swimtime="00:01:07.76" resultid="3565" heatid="5173" lane="3" entrytime="00:01:11.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="434" swimtime="00:01:08.13" resultid="3566" heatid="5260" lane="6" entrytime="00:01:08.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="424" swimtime="00:02:28.97" resultid="3567" heatid="5346" lane="3" entrytime="00:02:30.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:10.83" />
                    <SPLIT distance="150" swimtime="00:01:49.77" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Peret Saboia" birthdate="2009-11-25" gender="F" nation="BRA" license="342238" swrid="5600234" athleteid="3592" externalid="342238">
              <RESULTS>
                <RESULT eventid="1080" points="539" swimtime="00:01:18.79" resultid="3593" heatid="5069" lane="3" entrytime="00:01:18.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="418" swimtime="00:02:48.56" resultid="3594" heatid="5190" lane="8" entrytime="00:02:46.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="100" swimtime="00:01:24.08" />
                    <SPLIT distance="150" swimtime="00:02:11.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="469" swimtime="00:02:56.97" resultid="3595" heatid="5314" lane="7" entrytime="00:02:55.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.54" />
                    <SPLIT distance="100" swimtime="00:01:25.44" />
                    <SPLIT distance="150" swimtime="00:02:12.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="467" swimtime="00:00:37.58" resultid="3596" heatid="5377" lane="1" entrytime="00:00:37.40" entrycourse="LCM" />
                <RESULT eventid="2312" points="521" swimtime="00:01:19.69" resultid="5942" heatid="6416" lane="6" entrytime="00:01:18.79">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabelly" lastname="Sinnott" birthdate="2009-03-14" gender="F" nation="BRA" license="367255" swrid="5600258" athleteid="3523" externalid="367255">
              <RESULTS>
                <RESULT eventid="1064" points="589" swimtime="00:04:40.76" resultid="3524" heatid="5053" lane="4" entrytime="00:04:38.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.83" />
                    <SPLIT distance="100" swimtime="00:01:08.86" />
                    <SPLIT distance="150" swimtime="00:01:43.94" />
                    <SPLIT distance="200" swimtime="00:02:19.40" />
                    <SPLIT distance="250" swimtime="00:02:54.42" />
                    <SPLIT distance="300" swimtime="00:03:29.92" />
                    <SPLIT distance="350" swimtime="00:04:05.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="629" swimtime="00:02:11.70" resultid="3525" heatid="5144" lane="4" entrytime="00:02:10.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                    <SPLIT distance="100" swimtime="00:01:05.31" />
                    <SPLIT distance="150" swimtime="00:01:38.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="3526" heatid="5272" lane="4" entrytime="00:09:47.39" entrycourse="LCM" />
                <RESULT eventid="1279" status="DNS" swimtime="00:00:00.00" resultid="3527" heatid="5350" lane="3" entrytime="00:18:33.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Artigas Pinheiro" birthdate="2011-08-25" gender="M" nation="BRA" license="377040" swrid="5588535" athleteid="3861" externalid="377040">
              <RESULTS>
                <RESULT eventid="1088" points="295" swimtime="00:01:25.40" resultid="3862" heatid="5081" lane="4" entrytime="00:01:24.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="291" swimtime="00:02:51.99" resultid="3863" heatid="5194" lane="1" entrytime="00:02:52.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.52" />
                    <SPLIT distance="150" swimtime="00:02:13.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="327" swimtime="00:10:56.24" resultid="3864" heatid="5297" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.37" />
                    <SPLIT distance="100" swimtime="00:01:16.10" />
                    <SPLIT distance="150" swimtime="00:01:57.50" />
                    <SPLIT distance="200" swimtime="00:02:39.30" />
                    <SPLIT distance="250" swimtime="00:03:21.73" />
                    <SPLIT distance="300" swimtime="00:04:03.06" />
                    <SPLIT distance="350" swimtime="00:04:44.40" />
                    <SPLIT distance="400" swimtime="00:05:26.40" />
                    <SPLIT distance="450" swimtime="00:06:08.44" />
                    <SPLIT distance="500" swimtime="00:06:49.41" />
                    <SPLIT distance="550" swimtime="00:07:31.68" />
                    <SPLIT distance="600" swimtime="00:08:12.91" />
                    <SPLIT distance="650" swimtime="00:08:53.96" />
                    <SPLIT distance="700" swimtime="00:09:36.00" />
                    <SPLIT distance="750" swimtime="00:10:16.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="305" swimtime="00:03:06.34" resultid="3865" heatid="5317" lane="3" entrytime="00:03:04.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.55" />
                    <SPLIT distance="100" swimtime="00:01:29.98" />
                    <SPLIT distance="150" swimtime="00:02:19.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="264" swimtime="00:02:54.31" resultid="3866" heatid="5345" lane="8" entrytime="00:02:53.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.57" />
                    <SPLIT distance="100" swimtime="00:01:26.90" />
                    <SPLIT distance="150" swimtime="00:02:11.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Fontolan Gomes" birthdate="2010-07-02" gender="M" nation="BRA" license="356245" swrid="5588705" athleteid="3633" externalid="356245">
              <RESULTS>
                <RESULT eventid="1088" points="242" swimtime="00:01:31.18" resultid="3634" heatid="5080" lane="6" entrytime="00:01:31.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="384" swimtime="00:02:20.23" resultid="3635" heatid="5151" lane="1" entrytime="00:02:22.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.71" />
                    <SPLIT distance="100" swimtime="00:01:07.68" />
                    <SPLIT distance="150" swimtime="00:01:44.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="375" swimtime="00:01:11.50" resultid="3636" heatid="5257" lane="7" entrytime="00:01:12.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="332" swimtime="00:00:33.98" resultid="3637" heatid="5282" lane="5" />
                <RESULT eventid="1277" points="376" swimtime="00:02:34.99" resultid="3638" heatid="5346" lane="1" entrytime="00:02:35.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.44" />
                    <SPLIT distance="100" swimtime="00:01:14.36" />
                    <SPLIT distance="150" swimtime="00:01:54.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Rocha" birthdate="2011-08-25" gender="F" nation="BRA" license="366904" swrid="5602578" athleteid="3777" externalid="366904">
              <RESULTS>
                <RESULT eventid="1064" points="434" swimtime="00:05:10.75" resultid="3778" heatid="5050" lane="5" entrytime="00:05:08.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                    <SPLIT distance="100" swimtime="00:01:14.10" />
                    <SPLIT distance="150" swimtime="00:01:53.94" />
                    <SPLIT distance="200" swimtime="00:02:33.54" />
                    <SPLIT distance="250" swimtime="00:03:13.34" />
                    <SPLIT distance="300" swimtime="00:03:53.20" />
                    <SPLIT distance="350" swimtime="00:04:32.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="452" swimtime="00:00:30.75" resultid="3779" heatid="5100" lane="8" entrytime="00:00:30.30" entrycourse="LCM" />
                <RESULT eventid="1112" points="490" swimtime="00:02:23.12" resultid="3780" heatid="5141" lane="7" entrytime="00:02:24.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.65" />
                    <SPLIT distance="100" swimtime="00:01:10.21" />
                    <SPLIT distance="150" swimtime="00:01:46.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="480" swimtime="00:01:06.04" resultid="3781" heatid="5204" lane="3" entrytime="00:01:06.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1275" points="380" swimtime="00:02:49.91" resultid="3782" heatid="5342" lane="8" entrytime="00:02:48.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.24" />
                    <SPLIT distance="100" swimtime="00:01:23.17" />
                    <SPLIT distance="150" swimtime="00:02:07.26" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Krupacz" birthdate="2008-04-18" gender="F" nation="BRA" license="329187" swrid="5634611" athleteid="3940" externalid="329187">
              <RESULTS>
                <RESULT eventid="1143" points="435" swimtime="00:02:46.39" resultid="3941" heatid="5189" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                    <SPLIT distance="100" swimtime="00:01:12.15" />
                    <SPLIT distance="150" swimtime="00:02:06.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="592" swimtime="00:01:08.25" resultid="3942" heatid="5247" lane="4" entrytime="00:01:08.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="612" swimtime="00:00:31.62" resultid="3943" heatid="5295" lane="5" entrytime="00:00:31.74" entrycourse="LCM" />
                <RESULT eventid="1275" points="529" swimtime="00:02:32.25" resultid="3944" heatid="5343" lane="5" entrytime="00:02:31.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                    <SPLIT distance="100" swimtime="00:01:13.72" />
                    <SPLIT distance="150" swimtime="00:01:52.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2391" points="563" swimtime="00:01:09.41" resultid="6127" heatid="6424" lane="4" entrytime="00:01:08.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietra" lastname="Ruschel Carvalho" birthdate="2009-03-21" gender="F" nation="BRA" license="324999" swrid="5600250" athleteid="3473" externalid="324999">
              <RESULTS>
                <RESULT eventid="1096" points="632" swimtime="00:00:27.51" resultid="3474" heatid="5104" lane="4" entrytime="00:00:26.96" entrycourse="LCM" />
                <RESULT eventid="1112" points="583" swimtime="00:02:15.01" resultid="3475" heatid="5144" lane="5" entrytime="00:02:11.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                    <SPLIT distance="100" swimtime="00:01:05.21" />
                    <SPLIT distance="150" swimtime="00:01:39.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="613" swimtime="00:01:00.86" resultid="3476" heatid="5208" lane="4" entrytime="00:00:59.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="463" swimtime="00:00:31.57" resultid="3477" heatid="5326" lane="3" entrytime="00:00:31.15" entrycourse="LCM" />
                <RESULT eventid="2375" points="651" swimtime="00:00:27.23" resultid="5968" heatid="5978" lane="4" entrytime="00:00:27.51" />
                <RESULT eventid="2343" points="620" swimtime="00:01:00.63" resultid="6103" heatid="6421" lane="3" entrytime="00:01:00.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.81" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Pedro Pasqual" birthdate="2009-06-17" gender="M" nation="BRA" license="386136" swrid="5600232" athleteid="3976" externalid="386136">
              <RESULTS>
                <RESULT eventid="1104" points="546" swimtime="00:00:25.57" resultid="3977" heatid="5125" lane="3" entrytime="00:00:26.08" entrycourse="LCM" />
                <RESULT eventid="1182" points="634" swimtime="00:01:00.04" resultid="3978" heatid="5261" lane="3" entrytime="00:01:01.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="607" swimtime="00:00:27.80" resultid="3979" heatid="5288" lane="2" entrytime="00:00:28.62" entrycourse="LCM" />
                <RESULT eventid="1277" points="540" swimtime="00:02:17.41" resultid="3980" heatid="5348" lane="7" entrytime="00:02:16.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.95" />
                    <SPLIT distance="100" swimtime="00:01:07.23" />
                    <SPLIT distance="150" swimtime="00:01:43.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2359" points="592" swimtime="00:01:01.44" resultid="6143" heatid="6423" lane="3" entrytime="00:01:00.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gael" lastname="Gluck" birthdate="2011-01-28" gender="M" nation="BRA" license="366891" swrid="5588726" athleteid="3733" externalid="366891">
              <RESULTS>
                <RESULT eventid="1088" points="381" swimtime="00:01:18.43" resultid="3734" heatid="5082" lane="6" entrytime="00:01:18.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="429" swimtime="00:02:15.15" resultid="3735" heatid="5151" lane="4" entrytime="00:02:17.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                    <SPLIT distance="100" swimtime="00:01:04.86" />
                    <SPLIT distance="150" swimtime="00:01:40.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="377" swimtime="00:02:37.79" resultid="3736" heatid="5195" lane="7" entrytime="00:02:37.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                    <SPLIT distance="100" swimtime="00:01:17.19" />
                    <SPLIT distance="150" swimtime="00:02:01.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="379" swimtime="00:05:34.86" resultid="3737" heatid="5274" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:01:20.75" />
                    <SPLIT distance="150" swimtime="00:02:05.70" />
                    <SPLIT distance="200" swimtime="00:02:50.74" />
                    <SPLIT distance="250" swimtime="00:03:36.31" />
                    <SPLIT distance="300" swimtime="00:04:21.09" />
                    <SPLIT distance="350" swimtime="00:04:59.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="379" swimtime="00:02:53.24" resultid="3738" heatid="5318" lane="6" entrytime="00:02:48.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:22.28" />
                    <SPLIT distance="150" swimtime="00:02:08.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="371" swimtime="00:00:36.10" resultid="3739" heatid="5368" lane="1" entrytime="00:00:37.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nina" lastname="Rocha Ribeiro Da Silva" birthdate="2010-09-22" gender="F" nation="BRA" license="367216" swrid="5588884" athleteid="3884" externalid="367216">
              <RESULTS>
                <RESULT eventid="1080" status="DNS" swimtime="00:00:00.00" resultid="3885" heatid="5067" lane="4" entrytime="00:01:20.23" entrycourse="LCM" />
                <RESULT eventid="1143" status="DNS" swimtime="00:00:00.00" resultid="3886" heatid="5187" lane="6" entrytime="00:02:59.05" entrycourse="LCM" />
                <RESULT eventid="1159" status="DNS" swimtime="00:00:00.00" resultid="3887" heatid="5204" lane="8" entrytime="00:01:09.05" entrycourse="LCM" />
                <RESULT eventid="1243" status="SICK" swimtime="00:00:00.00" resultid="3888" heatid="5314" lane="8" entrytime="00:02:57.67" entrycourse="LCM" />
                <RESULT eventid="1305" status="SICK" swimtime="00:00:00.00" resultid="3889" heatid="5376" lane="4" entrytime="00:00:37.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicole" lastname="Rosario Osternack" birthdate="2008-04-11" gender="F" nation="BRA" license="331584" swrid="5600248" athleteid="3466" externalid="331584">
              <RESULTS>
                <RESULT eventid="1080" points="576" swimtime="00:01:17.04" resultid="3467" heatid="5069" lane="5" entrytime="00:01:18.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="557" swimtime="00:00:28.69" resultid="3468" heatid="5104" lane="6" entrytime="00:00:28.85" entrycourse="LCM" />
                <RESULT eventid="1143" points="575" swimtime="00:02:31.65" resultid="3469" heatid="5190" lane="4" entrytime="00:02:33.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                    <SPLIT distance="100" swimtime="00:01:12.04" />
                    <SPLIT distance="150" swimtime="00:01:56.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="500" swimtime="00:01:12.19" resultid="3470" heatid="5247" lane="5" entrytime="00:01:10.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="579" swimtime="00:01:02.02" resultid="3471" heatid="5208" lane="6" entrytime="00:01:02.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="513" swimtime="00:00:30.51" resultid="3472" heatid="5326" lane="5" entrytime="00:00:30.08" entrycourse="LCM" />
                <RESULT eventid="2312" points="537" swimtime="00:01:18.89" resultid="5940" heatid="6416" lane="3" entrytime="00:01:17.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2343" points="551" swimtime="00:01:03.04" resultid="6104" heatid="6421" lane="6" entrytime="00:01:02.02">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2391" points="498" swimtime="00:01:12.29" resultid="6465" heatid="6424" lane="7" entrytime="00:01:12.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Cury" birthdate="2005-09-28" gender="M" nation="BRA" license="329251" swrid="5600270" athleteid="3714" externalid="329251" level="SMELJ">
              <RESULTS>
                <RESULT eventid="1072" points="564" swimtime="00:04:26.29" resultid="3715" heatid="5064" lane="3" entrytime="00:04:31.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.22" />
                    <SPLIT distance="100" swimtime="00:01:03.64" />
                    <SPLIT distance="150" swimtime="00:01:37.83" />
                    <SPLIT distance="200" swimtime="00:02:12.42" />
                    <SPLIT distance="250" swimtime="00:02:47.48" />
                    <SPLIT distance="300" swimtime="00:03:21.82" />
                    <SPLIT distance="350" swimtime="00:03:54.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="596" swimtime="00:00:58.73" resultid="3716" heatid="5178" lane="2" entrytime="00:00:57.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="590" swimtime="00:00:55.85" resultid="3717" heatid="5232" lane="4" entrytime="00:00:54.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="379" swimtime="00:05:35.08" resultid="3718" heatid="5274" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                    <SPLIT distance="100" swimtime="00:01:09.25" />
                    <SPLIT distance="150" swimtime="00:01:55.32" />
                    <SPLIT distance="200" swimtime="00:02:41.83" />
                    <SPLIT distance="250" swimtime="00:03:31.18" />
                    <SPLIT distance="300" swimtime="00:04:21.91" />
                    <SPLIT distance="350" swimtime="00:05:01.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="573" swimtime="00:00:26.81" resultid="3719" heatid="5338" lane="6" entrytime="00:00:26.16" entrycourse="LCM" />
                <RESULT eventid="2335" points="610" swimtime="00:00:58.30" resultid="6015" heatid="6417" lane="8" entrytime="00:00:58.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Braun Prado" birthdate="2008-04-07" gender="M" nation="BRA" license="307663" swrid="5484324" athleteid="3622" externalid="307663">
              <RESULTS>
                <RESULT eventid="1072" points="488" swimtime="00:04:39.41" resultid="3623" heatid="5060" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                    <SPLIT distance="100" swimtime="00:01:03.91" />
                    <SPLIT distance="150" swimtime="00:01:39.00" />
                    <SPLIT distance="200" swimtime="00:02:15.52" />
                    <SPLIT distance="250" swimtime="00:02:51.72" />
                    <SPLIT distance="300" swimtime="00:03:27.93" />
                    <SPLIT distance="350" swimtime="00:04:04.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="493" swimtime="00:02:09.05" resultid="3624" heatid="5155" lane="4" entrytime="00:02:08.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.84" />
                    <SPLIT distance="100" swimtime="00:01:02.57" />
                    <SPLIT distance="150" swimtime="00:01:35.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="569" swimtime="00:01:02.27" resultid="3625" heatid="5261" lane="6" entrytime="00:01:02.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="488" swimtime="00:02:22.10" resultid="3626" heatid="5348" lane="2" entrytime="00:02:16.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                    <SPLIT distance="100" swimtime="00:01:08.14" />
                    <SPLIT distance="150" swimtime="00:01:44.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Henrique Pasqual" birthdate="2005-05-07" gender="M" nation="BRA" license="329284" swrid="5600185" athleteid="3981" externalid="329284">
              <RESULTS>
                <RESULT eventid="1104" points="663" swimtime="00:00:23.97" resultid="3982" heatid="5130" lane="6" entrytime="00:00:23.65" entrycourse="LCM" />
                <RESULT eventid="1135" points="603" swimtime="00:00:58.52" resultid="3983" heatid="5178" lane="7" entrytime="00:00:57.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="669" swimtime="00:00:53.56" resultid="3984" heatid="5233" lane="7" entrytime="00:00:53.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.51" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 6.3 - A cabeça não rompeu a superfície da água no ou antes do marco de 15m após o início ou a virada.  (Horário: 17:38)" eventid="1213" status="DSQ" swimtime="00:00:30.12" resultid="3985" heatid="5283" lane="8" />
                <RESULT eventid="1267" points="614" swimtime="00:00:26.20" resultid="3986" heatid="5338" lane="3" entrytime="00:00:25.31" entrycourse="LCM" />
                <RESULT eventid="2383" points="647" swimtime="00:00:24.17" resultid="5982" heatid="6425" lane="6" entrytime="00:00:23.97" />
                <RESULT eventid="2335" points="589" swimtime="00:00:58.96" resultid="6012" heatid="6417" lane="2" entrytime="00:00:58.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2351" points="656" swimtime="00:00:53.91" resultid="6121" heatid="6422" lane="7" entrytime="00:00:53.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Rocha Silva" birthdate="2007-10-10" gender="M" nation="BRA" license="372280" swrid="5717294" athleteid="3551" externalid="372280">
              <RESULTS>
                <RESULT eventid="1072" points="688" swimtime="00:04:09.26" resultid="3552" heatid="5063" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                    <SPLIT distance="100" swimtime="00:01:00.54" />
                    <SPLIT distance="150" swimtime="00:01:31.91" />
                    <SPLIT distance="200" swimtime="00:02:03.55" />
                    <SPLIT distance="250" swimtime="00:02:35.34" />
                    <SPLIT distance="300" swimtime="00:03:07.35" />
                    <SPLIT distance="350" swimtime="00:03:39.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="683" swimtime="00:00:23.74" resultid="3553" heatid="5130" lane="4" entrytime="00:00:23.42" entrycourse="LCM" />
                <RESULT eventid="1120" points="735" swimtime="00:01:52.98" resultid="3554" heatid="5158" lane="5" entrytime="00:01:52.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.11" />
                    <SPLIT distance="100" swimtime="00:00:56.24" />
                    <SPLIT distance="150" swimtime="00:01:25.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="765" swimtime="00:00:51.22" resultid="3555" heatid="5233" lane="4" entrytime="00:00:49.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="625" swimtime="00:08:48.53" resultid="3556" heatid="5296" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                    <SPLIT distance="100" swimtime="00:01:02.78" />
                    <SPLIT distance="150" swimtime="00:01:36.70" />
                    <SPLIT distance="200" swimtime="00:02:10.55" />
                    <SPLIT distance="250" swimtime="00:02:45.04" />
                    <SPLIT distance="300" swimtime="00:03:18.85" />
                    <SPLIT distance="350" swimtime="00:03:52.90" />
                    <SPLIT distance="400" swimtime="00:04:26.74" />
                    <SPLIT distance="450" swimtime="00:05:00.61" />
                    <SPLIT distance="500" swimtime="00:05:34.37" />
                    <SPLIT distance="550" swimtime="00:06:08.45" />
                    <SPLIT distance="600" swimtime="00:06:42.18" />
                    <SPLIT distance="650" swimtime="00:07:16.56" />
                    <SPLIT distance="700" swimtime="00:07:49.96" />
                    <SPLIT distance="750" swimtime="00:08:19.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2383" points="692" swimtime="00:00:23.64" resultid="5979" heatid="6425" lane="4" entrytime="00:00:23.74" />
                <RESULT eventid="2351" points="799" swimtime="00:00:50.48" resultid="6116" heatid="6422" lane="4" entrytime="00:00:51.22">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:24.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Schiavon" birthdate="2010-05-03" gender="M" nation="BRA" license="356354" swrid="5600256" athleteid="3677" externalid="356354">
              <RESULTS>
                <RESULT eventid="1072" points="507" swimtime="00:04:35.85" resultid="3678" heatid="5059" lane="3" entrytime="00:04:36.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                    <SPLIT distance="100" swimtime="00:01:06.65" />
                    <SPLIT distance="150" swimtime="00:01:42.03" />
                    <SPLIT distance="200" swimtime="00:02:17.81" />
                    <SPLIT distance="250" swimtime="00:02:52.44" />
                    <SPLIT distance="300" swimtime="00:03:27.38" />
                    <SPLIT distance="350" swimtime="00:04:01.90" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.4 - Movimentos das pernas não simultâneos.  (Horário: 18:56), (Medley Individual, Peito)." eventid="1151" status="DSQ" swimtime="00:02:29.50" resultid="3679" heatid="5195" lane="6" entrytime="00:02:30.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.64" />
                    <SPLIT distance="150" swimtime="00:01:54.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="353" swimtime="00:01:12.95" resultid="3680" heatid="5257" lane="5" entrytime="00:01:11.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="487" swimtime="00:09:34.29" resultid="3681" heatid="5300" lane="7" entrytime="00:09:35.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:08.00" />
                    <SPLIT distance="150" swimtime="00:01:43.99" />
                    <SPLIT distance="200" swimtime="00:02:20.40" />
                    <SPLIT distance="250" swimtime="00:02:56.10" />
                    <SPLIT distance="300" swimtime="00:03:32.81" />
                    <SPLIT distance="350" swimtime="00:04:09.12" />
                    <SPLIT distance="400" swimtime="00:04:45.08" />
                    <SPLIT distance="450" swimtime="00:05:21.40" />
                    <SPLIT distance="500" swimtime="00:05:58.28" />
                    <SPLIT distance="550" swimtime="00:06:35.06" />
                    <SPLIT distance="600" swimtime="00:07:11.25" />
                    <SPLIT distance="650" swimtime="00:07:47.59" />
                    <SPLIT distance="700" swimtime="00:08:24.50" />
                    <SPLIT distance="750" swimtime="00:08:59.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="403" swimtime="00:02:31.46" resultid="3682" heatid="5344" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.44" />
                    <SPLIT distance="100" swimtime="00:01:16.54" />
                    <SPLIT distance="150" swimtime="00:01:53.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="483" swimtime="00:18:29.64" resultid="3683" heatid="5380" lane="2" entrytime="00:18:07.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.69" />
                    <SPLIT distance="100" swimtime="00:01:09.16" />
                    <SPLIT distance="150" swimtime="00:01:46.61" />
                    <SPLIT distance="200" swimtime="00:02:24.21" />
                    <SPLIT distance="250" swimtime="00:03:01.64" />
                    <SPLIT distance="300" swimtime="00:03:39.27" />
                    <SPLIT distance="350" swimtime="00:04:16.23" />
                    <SPLIT distance="400" swimtime="00:04:53.72" />
                    <SPLIT distance="450" swimtime="00:05:31.25" />
                    <SPLIT distance="500" swimtime="00:06:08.33" />
                    <SPLIT distance="550" swimtime="00:06:44.72" />
                    <SPLIT distance="600" swimtime="00:07:21.78" />
                    <SPLIT distance="650" swimtime="00:07:58.26" />
                    <SPLIT distance="700" swimtime="00:08:35.29" />
                    <SPLIT distance="750" swimtime="00:09:11.91" />
                    <SPLIT distance="800" swimtime="00:09:48.85" />
                    <SPLIT distance="850" swimtime="00:10:26.09" />
                    <SPLIT distance="900" swimtime="00:11:03.25" />
                    <SPLIT distance="950" swimtime="00:11:40.19" />
                    <SPLIT distance="1000" swimtime="00:12:17.27" />
                    <SPLIT distance="1050" swimtime="00:12:54.75" />
                    <SPLIT distance="1100" swimtime="00:13:32.04" />
                    <SPLIT distance="1150" swimtime="00:14:09.50" />
                    <SPLIT distance="1200" swimtime="00:14:46.88" />
                    <SPLIT distance="1250" swimtime="00:15:24.03" />
                    <SPLIT distance="1300" swimtime="00:16:01.77" />
                    <SPLIT distance="1350" swimtime="00:16:40.02" />
                    <SPLIT distance="1400" swimtime="00:17:18.09" />
                    <SPLIT distance="1450" swimtime="00:17:53.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Brandt De Macedo" birthdate="2010-01-13" gender="M" nation="BRA" license="338925" swrid="5588565" athleteid="3710" externalid="338925">
              <RESULTS>
                <RESULT eventid="1104" points="434" swimtime="00:00:27.60" resultid="3711" heatid="5119" lane="7" entrytime="00:00:28.33" entrycourse="LCM" />
                <RESULT eventid="1135" points="291" swimtime="00:01:14.58" resultid="3712" heatid="5170" lane="2" entrytime="00:01:19.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="459" swimtime="00:02:12.22" resultid="3713" heatid="5152" lane="7" entrytime="00:02:12.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                    <SPLIT distance="100" swimtime="00:01:03.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Galvao" birthdate="2011-03-11" gender="M" nation="BRA" license="381989" swrid="5602541" athleteid="3873" externalid="381989">
              <RESULTS>
                <RESULT eventid="1072" points="329" swimtime="00:05:18.51" resultid="3874" heatid="5057" lane="6" entrytime="00:05:16.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.54" />
                    <SPLIT distance="100" swimtime="00:01:13.57" />
                    <SPLIT distance="150" swimtime="00:01:54.71" />
                    <SPLIT distance="200" swimtime="00:02:36.96" />
                    <SPLIT distance="250" swimtime="00:03:18.85" />
                    <SPLIT distance="300" swimtime="00:04:00.37" />
                    <SPLIT distance="350" swimtime="00:04:40.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="306" swimtime="00:00:31.01" resultid="3875" heatid="5116" lane="4" entrytime="00:00:31.07" entrycourse="LCM" />
                <RESULT eventid="1120" points="268" swimtime="00:02:38.15" resultid="3876" heatid="5150" lane="6" entrytime="00:02:27.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:15.59" />
                    <SPLIT distance="150" swimtime="00:01:58.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="354" swimtime="00:01:06.21" resultid="3877" heatid="5220" lane="6" entrytime="00:01:07.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="215" swimtime="00:03:06.63" resultid="3878" heatid="5344" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.07" />
                    <SPLIT distance="100" swimtime="00:01:32.85" />
                    <SPLIT distance="150" swimtime="00:02:21.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="323" swimtime="00:21:09.31" resultid="3879" heatid="5378" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                    <SPLIT distance="100" swimtime="00:01:17.16" />
                    <SPLIT distance="150" swimtime="00:01:59.48" />
                    <SPLIT distance="200" swimtime="00:02:41.50" />
                    <SPLIT distance="250" swimtime="00:03:24.73" />
                    <SPLIT distance="300" swimtime="00:04:06.80" />
                    <SPLIT distance="350" swimtime="00:04:50.17" />
                    <SPLIT distance="400" swimtime="00:05:31.84" />
                    <SPLIT distance="450" swimtime="00:06:14.57" />
                    <SPLIT distance="500" swimtime="00:06:57.00" />
                    <SPLIT distance="550" swimtime="00:07:40.51" />
                    <SPLIT distance="600" swimtime="00:08:23.33" />
                    <SPLIT distance="650" swimtime="00:09:06.84" />
                    <SPLIT distance="700" swimtime="00:09:49.12" />
                    <SPLIT distance="750" swimtime="00:10:32.51" />
                    <SPLIT distance="800" swimtime="00:11:15.60" />
                    <SPLIT distance="850" swimtime="00:11:58.77" />
                    <SPLIT distance="900" swimtime="00:12:41.43" />
                    <SPLIT distance="950" swimtime="00:13:25.03" />
                    <SPLIT distance="1000" swimtime="00:14:07.86" />
                    <SPLIT distance="1050" swimtime="00:14:51.55" />
                    <SPLIT distance="1100" swimtime="00:15:34.39" />
                    <SPLIT distance="1150" swimtime="00:16:17.41" />
                    <SPLIT distance="1200" swimtime="00:17:00.27" />
                    <SPLIT distance="1250" swimtime="00:17:43.53" />
                    <SPLIT distance="1300" swimtime="00:18:26.89" />
                    <SPLIT distance="1350" swimtime="00:19:09.89" />
                    <SPLIT distance="1400" swimtime="00:19:51.04" />
                    <SPLIT distance="1450" swimtime="00:20:32.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Estela" lastname="Albuquerque" birthdate="2010-11-23" gender="F" nation="BRA" license="356344" swrid="5653285" athleteid="3658" externalid="356344">
              <RESULTS>
                <RESULT eventid="1064" points="464" swimtime="00:05:03.95" resultid="3659" heatid="5051" lane="3" entrytime="00:05:01.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="150" swimtime="00:01:51.24" />
                    <SPLIT distance="250" swimtime="00:03:09.24" />
                    <SPLIT distance="350" swimtime="00:04:26.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="415" swimtime="00:00:31.65" resultid="3660" heatid="5099" lane="3" entrytime="00:00:31.26" entrycourse="LCM" />
                <RESULT eventid="1112" points="498" swimtime="00:02:22.35" resultid="3661" heatid="5141" lane="3" entrytime="00:02:22.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:08.79" />
                    <SPLIT distance="150" swimtime="00:01:46.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="334" swimtime="00:01:22.56" resultid="3662" heatid="5243" lane="3" entrytime="00:01:18.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="454" swimtime="00:01:07.25" resultid="3663" heatid="5204" lane="4" entrytime="00:01:06.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Fontes Bonardi" birthdate="2008-10-26" gender="M" nation="BRA" license="307662" swrid="5600164" athleteid="3491" externalid="307662">
              <RESULTS>
                <RESULT eventid="1088" points="523" swimtime="00:01:10.59" resultid="3492" heatid="5085" lane="7" entrytime="00:01:09.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="651" swimtime="00:02:11.48" resultid="3493" heatid="5198" lane="4" entrytime="00:02:12.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.67" />
                    <SPLIT distance="100" swimtime="00:01:01.56" />
                    <SPLIT distance="150" swimtime="00:01:39.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="615" swimtime="00:00:55.09" resultid="3494" heatid="5224" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="565" swimtime="00:04:53.29" resultid="3495" heatid="5277" lane="5" entrytime="00:04:48.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                    <SPLIT distance="100" swimtime="00:01:05.81" />
                    <SPLIT distance="150" swimtime="00:01:45.57" />
                    <SPLIT distance="250" swimtime="00:03:05.56" />
                    <SPLIT distance="300" swimtime="00:03:46.16" />
                    <SPLIT distance="350" swimtime="00:04:21.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="566" swimtime="00:02:31.62" resultid="3496" heatid="5320" lane="3" entrytime="00:02:27.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                    <SPLIT distance="100" swimtime="00:01:12.80" />
                    <SPLIT distance="150" swimtime="00:01:52.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Lacerda" birthdate="2011-05-09" gender="M" nation="BRA" license="366909" swrid="5602550" athleteid="3801" externalid="366909">
              <RESULTS>
                <RESULT eventid="1088" points="261" swimtime="00:01:28.95" resultid="3802" heatid="5081" lane="2" entrytime="00:01:27.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="340" swimtime="00:02:43.21" resultid="3803" heatid="5194" lane="4" entrytime="00:02:42.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.38" />
                    <SPLIT distance="100" swimtime="00:01:20.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="266" swimtime="00:01:20.17" resultid="3804" heatid="5255" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="335" swimtime="00:05:48.83" resultid="3805" heatid="5276" lane="1" entrytime="00:05:45.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                    <SPLIT distance="100" swimtime="00:01:24.36" />
                    <SPLIT distance="150" swimtime="00:02:10.67" />
                    <SPLIT distance="250" swimtime="00:03:45.28" />
                    <SPLIT distance="300" swimtime="00:04:34.63" />
                    <SPLIT distance="350" swimtime="00:05:12.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="291" swimtime="00:03:09.30" resultid="3806" heatid="5317" lane="7" entrytime="00:03:09.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.55" />
                    <SPLIT distance="100" swimtime="00:01:32.15" />
                    <SPLIT distance="150" swimtime="00:02:22.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucca" lastname="Cruz Tonin" birthdate="2004-03-19" gender="M" nation="BRA" license="270821" swrid="5622272" athleteid="3807" externalid="270821" level="FUNDESPORT">
              <RESULTS>
                <RESULT eventid="1104" points="674" swimtime="00:00:23.84" resultid="3808" heatid="5130" lane="7" entrytime="00:00:24.08" entrycourse="LCM" />
                <RESULT eventid="1135" points="694" swimtime="00:00:55.85" resultid="3809" heatid="5178" lane="3" entrytime="00:00:56.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="758" swimtime="00:00:56.58" resultid="3810" heatid="5263" lane="4" entrytime="00:00:56.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="739" swimtime="00:00:51.83" resultid="3811" heatid="5233" lane="6" entrytime="00:00:51.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="683" swimtime="00:00:26.74" resultid="3812" heatid="5288" lane="4" entrytime="00:00:26.50" entrycourse="LCM" />
                <RESULT eventid="1277" points="708" swimtime="00:02:05.57" resultid="3813" heatid="5348" lane="4" entrytime="00:02:02.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.75" />
                    <SPLIT distance="100" swimtime="00:01:00.27" />
                    <SPLIT distance="150" swimtime="00:01:33.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2383" points="654" swimtime="00:00:24.08" resultid="5980" heatid="6425" lane="5" entrytime="00:00:23.84" />
                <RESULT eventid="2335" points="706" swimtime="00:00:55.52" resultid="6008" heatid="6417" lane="4" entrytime="00:00:55.85">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2351" points="683" swimtime="00:00:53.19" resultid="6117" heatid="6422" lane="5" entrytime="00:00:51.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2359" points="738" swimtime="00:00:57.08" resultid="6141" heatid="6423" lane="4" entrytime="00:00:56.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joshua" lastname="Gomide Capraro" birthdate="2009-01-18" gender="M" nation="BRA" license="339030" swrid="5600177" athleteid="3497" externalid="339030">
              <RESULTS>
                <RESULT eventid="1104" points="597" swimtime="00:00:24.82" resultid="3498" heatid="5126" lane="3" entrytime="00:00:24.57" entrycourse="LCM" />
                <RESULT eventid="1120" points="576" swimtime="00:02:02.55" resultid="3499" heatid="5156" lane="2" entrytime="00:02:02.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.85" />
                    <SPLIT distance="100" swimtime="00:00:59.94" />
                    <SPLIT distance="150" swimtime="00:01:31.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="632" swimtime="00:00:54.58" resultid="3500" heatid="5230" lane="6" entrytime="00:00:55.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="472" swimtime="00:00:28.59" resultid="3501" heatid="5330" lane="3" />
                <RESULT eventid="2383" swimtime="00:00:00.00" resultid="5987" entrytime="00:00:24.82" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Fantin Dias De Andrade" birthdate="2010-11-06" gender="F" nation="BRA" license="339262" swrid="5588684" athleteid="3832" externalid="339262">
              <RESULTS>
                <RESULT eventid="1080" points="288" swimtime="00:01:37.01" resultid="3833" heatid="5066" lane="8" entrytime="00:01:33.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="351" swimtime="00:00:33.44" resultid="3834" heatid="5098" lane="6" entrytime="00:00:32.41" entrycourse="LCM" />
                <RESULT eventid="1128" points="231" swimtime="00:01:30.33" resultid="3835" heatid="5159" lane="3" entrytime="00:01:33.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="323" swimtime="00:03:03.76" resultid="3836" heatid="5187" lane="2" entrytime="00:03:00.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.68" />
                    <SPLIT distance="100" swimtime="00:01:30.04" />
                    <SPLIT distance="150" swimtime="00:02:24.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="258" swimtime="00:01:30.02" resultid="3837" heatid="5242" lane="1" entrytime="00:01:29.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Magalhaes Dos Reis" birthdate="2010-05-05" gender="M" nation="BRA" license="356361" swrid="5600207" athleteid="3690" externalid="356361">
              <RESULTS>
                <RESULT comment="SW 7.1 - A cabeça não rompeu a superfície antes que as mãos se virassem para dentro na parte mais ampla do segundo movimento após o início ou a virada.&#10;&#10;&#10;&#10;&#10;&#10;&#10;  (Horário: 11:34), Na saída." eventid="1088" status="DSQ" swimtime="00:01:20.46" resultid="3691" heatid="5082" lane="2" entrytime="00:01:20.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="428" swimtime="00:00:27.74" resultid="3692" heatid="5119" lane="3" entrytime="00:00:27.69" entrycourse="LCM" />
                <RESULT eventid="1151" points="376" swimtime="00:02:37.91" resultid="3693" heatid="5194" lane="5" entrytime="00:02:43.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.06" />
                    <SPLIT distance="100" swimtime="00:01:16.39" />
                    <SPLIT distance="150" swimtime="00:02:03.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="485" swimtime="00:00:59.61" resultid="3694" heatid="5223" lane="8" entrytime="00:01:00.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="282" swimtime="00:00:39.55" resultid="3695" heatid="5364" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Felipe Paes Feres" birthdate="2008-07-28" gender="M" nation="BRA" license="307676" swrid="5600156" athleteid="3568" externalid="307676">
              <RESULTS>
                <RESULT eventid="1104" points="477" swimtime="00:00:26.75" resultid="3569" heatid="5124" lane="2" entrytime="00:00:26.89" entrycourse="LCM" />
                <RESULT eventid="1151" points="464" swimtime="00:02:27.17" resultid="3570" heatid="5197" lane="2" entrytime="00:02:29.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.12" />
                    <SPLIT distance="100" swimtime="00:01:06.88" />
                    <SPLIT distance="150" swimtime="00:01:52.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="471" swimtime="00:01:06.30" resultid="3571" heatid="5261" lane="8" entrytime="00:01:06.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="408" swimtime="00:05:26.76" resultid="3572" heatid="5274" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.16" />
                    <SPLIT distance="100" swimtime="00:01:10.12" />
                    <SPLIT distance="150" swimtime="00:01:52.94" />
                    <SPLIT distance="200" swimtime="00:02:33.87" />
                    <SPLIT distance="250" swimtime="00:03:21.16" />
                    <SPLIT distance="300" swimtime="00:04:10.73" />
                    <SPLIT distance="350" swimtime="00:04:49.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="460" swimtime="00:02:24.98" resultid="3573" heatid="5347" lane="4" entrytime="00:02:23.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.09" />
                    <SPLIT distance="100" swimtime="00:01:08.60" />
                    <SPLIT distance="150" swimtime="00:01:46.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Zaroni" birthdate="2010-03-03" gender="F" nation="BRA" license="356345" swrid="5600282" athleteid="3528" externalid="356345">
              <RESULTS>
                <RESULT eventid="1080" points="475" swimtime="00:01:22.19" resultid="3529" heatid="5067" lane="3" entrytime="00:01:21.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="410" swimtime="00:02:49.76" resultid="3530" heatid="5188" lane="8" entrytime="00:02:48.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.02" />
                    <SPLIT distance="100" swimtime="00:01:24.46" />
                    <SPLIT distance="150" swimtime="00:02:12.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="468" swimtime="00:01:06.60" resultid="3531" heatid="5205" lane="7" entrytime="00:01:05.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="303" swimtime="00:00:36.35" resultid="3532" heatid="5321" lane="7" />
                <RESULT eventid="1243" points="422" swimtime="00:03:03.34" resultid="3533" heatid="5314" lane="1" entrytime="00:02:56.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.76" />
                    <SPLIT distance="100" swimtime="00:01:29.21" />
                    <SPLIT distance="150" swimtime="00:02:16.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Guimaraes E Souza" birthdate="2008-12-21" gender="M" nation="BRA" license="376972" swrid="5600182" athleteid="3856" externalid="376972">
              <RESULTS>
                <RESULT eventid="1088" points="544" swimtime="00:01:09.64" resultid="3857" heatid="5085" lane="6" entrytime="00:01:09.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="486" swimtime="00:02:24.98" resultid="3858" heatid="5197" lane="4" entrytime="00:02:25.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:11.16" />
                    <SPLIT distance="150" swimtime="00:01:54.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="490" swimtime="00:02:39.12" resultid="3859" heatid="5319" lane="4" entrytime="00:02:39.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:17.52" />
                    <SPLIT distance="150" swimtime="00:02:00.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="549" swimtime="00:00:31.68" resultid="3860" heatid="5370" lane="5" entrytime="00:00:32.22" entrycourse="LCM" />
                <RESULT eventid="2320" points="547" swimtime="00:01:09.55" resultid="5960" heatid="6414" lane="8" entrytime="00:01:09.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Valduga Artigas" birthdate="2009-06-01" gender="M" nation="BRA" license="339569" swrid="5600268" athleteid="3613" externalid="339569">
              <RESULTS>
                <RESULT eventid="1167" points="357" swimtime="00:01:06.01" resultid="3614" heatid="5225" lane="6" entrytime="00:01:05.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="317" swimtime="00:00:32.63" resultid="3615" heatid="5332" lane="3" entrytime="00:00:32.57" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Prosdocimo" birthdate="2010-11-23" gender="F" nation="BRA" license="356251" swrid="5600238" athleteid="3651" externalid="356251">
              <RESULTS>
                <RESULT eventid="1064" points="437" swimtime="00:05:10.05" resultid="3652" heatid="5051" lane="1" entrytime="00:05:05.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:13.35" />
                    <SPLIT distance="150" swimtime="00:01:52.98" />
                    <SPLIT distance="200" swimtime="00:02:32.24" />
                    <SPLIT distance="250" swimtime="00:03:12.73" />
                    <SPLIT distance="300" swimtime="00:03:52.13" />
                    <SPLIT distance="350" swimtime="00:04:32.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="465" swimtime="00:00:30.46" resultid="3653" heatid="5099" lane="4" entrytime="00:00:30.62" entrycourse="LCM" />
                <RESULT eventid="1112" points="482" swimtime="00:02:23.92" resultid="3654" heatid="5141" lane="2" entrytime="00:02:23.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.75" />
                    <SPLIT distance="100" swimtime="00:01:09.39" />
                    <SPLIT distance="150" swimtime="00:01:47.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="402" swimtime="00:01:17.65" resultid="3655" heatid="5244" lane="3" entrytime="00:01:15.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="469" swimtime="00:01:06.54" resultid="3656" heatid="5205" lane="6" entrytime="00:01:05.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1275" points="399" swimtime="00:02:47.17" resultid="3657" heatid="5341" lane="4" entrytime="00:02:48.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.03" />
                    <SPLIT distance="100" swimtime="00:01:22.31" />
                    <SPLIT distance="150" swimtime="00:02:05.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Trevisan" birthdate="2000-11-28" gender="M" nation="BRA" license="346847" swrid="5600266" athleteid="3890" externalid="346847">
              <RESULTS>
                <RESULT eventid="1104" points="614" swimtime="00:00:24.60" resultid="3891" heatid="5130" lane="8" entrytime="00:00:24.39" entrycourse="LCM" />
                <RESULT eventid="1120" points="511" swimtime="00:02:07.56" resultid="3892" heatid="5158" lane="2" entrytime="00:02:03.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.15" />
                    <SPLIT distance="100" swimtime="00:01:01.92" />
                    <SPLIT distance="150" swimtime="00:01:35.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="614" swimtime="00:00:55.12" resultid="3893" heatid="5232" lane="5" entrytime="00:00:54.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="524" swimtime="00:00:29.21" resultid="3894" heatid="5287" lane="3" entrytime="00:00:29.40" entrycourse="LCM" />
                <RESULT eventid="1267" points="556" swimtime="00:00:27.07" resultid="3895" heatid="5338" lane="1" entrytime="00:00:26.77" entrycourse="LCM" />
                <RESULT eventid="2383" points="627" swimtime="00:00:24.42" resultid="5986" heatid="6425" lane="8" entrytime="00:00:24.60" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mariana" lastname="Stoberl" birthdate="2010-07-09" gender="F" nation="BRA" license="356250" swrid="5600265" athleteid="3645" externalid="356250">
              <RESULTS>
                <RESULT eventid="1096" points="521" swimtime="00:00:29.33" resultid="3646" heatid="5100" lane="4" entrytime="00:00:29.08" entrycourse="LCM" />
                <RESULT eventid="1112" points="513" swimtime="00:02:20.97" resultid="3647" heatid="5141" lane="4" entrytime="00:02:17.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.79" />
                    <SPLIT distance="100" swimtime="00:01:08.60" />
                    <SPLIT distance="150" swimtime="00:01:44.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="402" swimtime="00:02:50.87" resultid="3648" heatid="5186" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.30" />
                    <SPLIT distance="100" swimtime="00:01:19.34" />
                    <SPLIT distance="150" swimtime="00:02:12.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="516" swimtime="00:01:04.45" resultid="3649" heatid="5205" lane="4" entrytime="00:01:03.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1275" points="407" swimtime="00:02:46.04" resultid="3650" heatid="5342" lane="5" entrytime="00:02:45.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:21.34" />
                    <SPLIT distance="150" swimtime="00:02:04.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2375" swimtime="00:00:00.00" resultid="6451" entrytime="00:00:29.33" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabela" lastname="Mattioli" birthdate="2011-10-22" gender="F" nation="BRA" license="366896" swrid="5602559" athleteid="3743" externalid="366896">
              <RESULTS>
                <RESULT eventid="1080" points="446" swimtime="00:01:23.91" resultid="3744" heatid="5067" lane="2" entrytime="00:01:23.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" points="450" swimtime="00:05:06.99" resultid="3745" heatid="5051" lane="7" entrytime="00:05:04.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.17" />
                    <SPLIT distance="100" swimtime="00:01:12.66" />
                    <SPLIT distance="150" swimtime="00:01:52.09" />
                    <SPLIT distance="200" swimtime="00:02:32.09" />
                    <SPLIT distance="250" swimtime="00:03:11.68" />
                    <SPLIT distance="300" swimtime="00:03:51.41" />
                    <SPLIT distance="350" swimtime="00:04:30.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="440" swimtime="00:02:45.79" resultid="3746" heatid="5188" lane="7" entrytime="00:02:44.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.16" />
                    <SPLIT distance="100" swimtime="00:01:21.34" />
                    <SPLIT distance="150" swimtime="00:02:08.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="441" swimtime="00:01:07.91" resultid="3747" heatid="5204" lane="6" entrytime="00:01:07.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="428" swimtime="00:03:02.50" resultid="3748" heatid="5313" lane="3" entrytime="00:02:58.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.30" />
                    <SPLIT distance="100" swimtime="00:01:26.99" />
                    <SPLIT distance="150" swimtime="00:02:16.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="428" swimtime="00:00:38.69" resultid="3749" heatid="5375" lane="7" entrytime="00:00:42.95" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo" lastname="Gabriel Nascimento" birthdate="2008-11-14" gender="M" nation="BRA" license="348028" swrid="5600171" athleteid="3909" externalid="348028" level="BIG BUM">
              <RESULTS>
                <RESULT eventid="1104" points="467" swimtime="00:00:26.94" resultid="3910" heatid="5124" lane="5" entrytime="00:00:26.68" entrycourse="LCM" />
                <RESULT eventid="1135" points="474" swimtime="00:01:03.42" resultid="3911" heatid="5174" lane="6" entrytime="00:01:03.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="471" swimtime="00:01:00.20" resultid="3912" heatid="5227" lane="3" entrytime="00:00:59.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="509" swimtime="00:00:27.88" resultid="3913" heatid="5335" lane="4" entrytime="00:00:28.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Sachser Rocha" birthdate="2008-07-09" gender="M" nation="BRA" license="330072" swrid="5600254" athleteid="3574" externalid="330072">
              <RESULTS>
                <RESULT eventid="1104" points="554" swimtime="00:00:25.45" resultid="3575" heatid="5126" lane="8" entrytime="00:00:25.46" entrycourse="LCM" />
                <RESULT eventid="1135" points="584" swimtime="00:00:59.16" resultid="3576" heatid="5175" lane="4" entrytime="00:00:58.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="538" swimtime="00:00:57.59" resultid="3577" heatid="5229" lane="2" entrytime="00:00:57.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="568" swimtime="00:00:26.88" resultid="3578" heatid="5338" lane="7" entrytime="00:00:26.63" entrycourse="LCM" />
                <RESULT eventid="1293" status="DNS" swimtime="00:00:00.00" resultid="3579" heatid="5359" lane="3" entrytime="00:02:28.20" entrycourse="LCM" />
                <RESULT eventid="2335" swimtime="00:00:00.00" resultid="6017" entrytime="00:00:59.16" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Novak Bredt" birthdate="2009-09-08" gender="F" nation="BRA" license="338909" swrid="5622297" athleteid="3534" externalid="338909">
              <RESULTS>
                <RESULT eventid="1080" points="451" swimtime="00:01:23.59" resultid="3535" heatid="5069" lane="1" entrytime="00:01:21.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="450" swimtime="00:02:44.50" resultid="3536" heatid="5190" lane="2" entrytime="00:02:42.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                    <SPLIT distance="100" swimtime="00:01:18.86" />
                    <SPLIT distance="150" swimtime="00:02:06.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="412" swimtime="00:03:04.74" resultid="3537" heatid="5313" lane="4" entrytime="00:02:58.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:26.80" />
                    <SPLIT distance="150" swimtime="00:02:16.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="446" swimtime="00:00:38.16" resultid="3538" heatid="5376" lane="5" entrytime="00:00:38.07" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="De Czarnecki" birthdate="2008-06-24" gender="M" nation="BRA" license="329641" swrid="5600146" athleteid="3485" externalid="329641">
              <RESULTS>
                <RESULT eventid="1072" points="576" swimtime="00:04:24.45" resultid="3486" heatid="5062" lane="2" entrytime="00:04:24.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.02" />
                    <SPLIT distance="100" swimtime="00:01:03.09" />
                    <SPLIT distance="150" swimtime="00:01:35.55" />
                    <SPLIT distance="200" swimtime="00:02:08.82" />
                    <SPLIT distance="250" swimtime="00:02:41.90" />
                    <SPLIT distance="300" swimtime="00:03:15.92" />
                    <SPLIT distance="350" swimtime="00:03:50.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="632" swimtime="00:01:58.81" resultid="3487" heatid="5156" lane="8" entrytime="00:02:08.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.32" />
                    <SPLIT distance="100" swimtime="00:00:58.51" />
                    <SPLIT distance="150" swimtime="00:01:28.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="606" swimtime="00:01:00.97" resultid="3488" heatid="5261" lane="4" entrytime="00:01:00.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="551" swimtime="00:00:28.72" resultid="3489" heatid="5287" lane="5" entrytime="00:00:28.92" entrycourse="LCM" />
                <RESULT eventid="1277" points="569" swimtime="00:02:15.03" resultid="3490" heatid="5348" lane="3" entrytime="00:02:11.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.24" />
                    <SPLIT distance="100" swimtime="00:01:04.52" />
                    <SPLIT distance="150" swimtime="00:01:39.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rene" lastname="Osternack Erbe" birthdate="2011-04-03" gender="M" nation="BRA" license="366907" swrid="5588842" athleteid="3789" externalid="366907">
              <RESULTS>
                <RESULT eventid="1072" points="352" swimtime="00:05:11.61" resultid="3790" heatid="5058" lane="8" entrytime="00:05:10.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.54" />
                    <SPLIT distance="100" swimtime="00:01:15.50" />
                    <SPLIT distance="150" swimtime="00:01:55.83" />
                    <SPLIT distance="200" swimtime="00:02:36.46" />
                    <SPLIT distance="250" swimtime="00:03:15.89" />
                    <SPLIT distance="300" swimtime="00:03:55.84" />
                    <SPLIT distance="350" swimtime="00:04:35.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="217" swimtime="00:01:22.18" resultid="3791" heatid="5170" lane="1" entrytime="00:01:25.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="294" swimtime="00:02:51.26" resultid="3792" heatid="5194" lane="8" entrytime="00:02:53.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.87" />
                    <SPLIT distance="100" swimtime="00:01:21.00" />
                    <SPLIT distance="150" swimtime="00:02:16.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="309" swimtime="00:01:16.32" resultid="3793" heatid="5257" lane="8" entrytime="00:01:18.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="304" swimtime="00:02:46.41" resultid="3794" heatid="5345" lane="2" entrytime="00:02:46.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.93" />
                    <SPLIT distance="100" swimtime="00:01:20.06" />
                    <SPLIT distance="150" swimtime="00:02:03.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Araujo Barros" birthdate="2008-12-26" gender="M" nation="BRA" license="331713" swrid="5367497" athleteid="3820" externalid="331713">
              <RESULTS>
                <RESULT eventid="1072" points="617" swimtime="00:04:18.38" resultid="3821" heatid="5062" lane="5" entrytime="00:04:19.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.90" />
                    <SPLIT distance="100" swimtime="00:01:01.88" />
                    <SPLIT distance="150" swimtime="00:01:35.20" />
                    <SPLIT distance="200" swimtime="00:02:08.22" />
                    <SPLIT distance="250" swimtime="00:02:40.66" />
                    <SPLIT distance="300" swimtime="00:03:13.21" />
                    <SPLIT distance="350" swimtime="00:03:46.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="596" swimtime="00:02:01.20" resultid="3822" heatid="5156" lane="5" entrytime="00:02:00.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.77" />
                    <SPLIT distance="100" swimtime="00:00:57.72" />
                    <SPLIT distance="150" swimtime="00:01:29.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="510" swimtime="00:00:27.87" resultid="3823" heatid="5328" lane="2" />
                <RESULT eventid="1293" points="436" swimtime="00:02:25.42" resultid="3824" heatid="5359" lane="4" entrytime="00:02:26.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.50" />
                    <SPLIT distance="100" swimtime="00:01:07.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Estevao" lastname="Valduga Artigas" birthdate="2009-06-01" gender="M" nation="BRA" license="339556" swrid="5600267" athleteid="3584" externalid="339556">
              <RESULTS>
                <RESULT eventid="1104" points="322" swimtime="00:00:30.48" resultid="3585" heatid="5121" lane="6" entrytime="00:00:31.53" entrycourse="LCM" />
                <RESULT eventid="1182" status="DNS" swimtime="00:00:00.00" resultid="3586" heatid="5260" lane="1" entrytime="00:01:18.18" entrycourse="LCM" />
                <RESULT eventid="1217" status="DNS" swimtime="00:00:00.00" resultid="3587" heatid="5298" lane="7" entrytime="00:10:47.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Ramos Marcon" birthdate="2008-01-12" gender="M" nation="BRA" license="372281" swrid="5600240" athleteid="3880" externalid="372281">
              <RESULTS>
                <RESULT eventid="1104" points="564" swimtime="00:00:25.30" resultid="3881" heatid="5126" lane="6" entrytime="00:00:24.82" entrycourse="LCM" />
                <RESULT eventid="1120" points="506" swimtime="00:02:07.95" resultid="3882" heatid="5156" lane="1" entrytime="00:02:08.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                    <SPLIT distance="100" swimtime="00:01:01.44" />
                    <SPLIT distance="150" swimtime="00:01:33.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="594" swimtime="00:00:55.73" resultid="3883" heatid="5230" lane="2" entrytime="00:00:55.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pablo" lastname="Souza Tavares" birthdate="2006-05-03" gender="M" nation="BRA" license="331982" swrid="5600261" athleteid="3478" externalid="331982" level="SMELJ/ECOI">
              <RESULTS>
                <RESULT eventid="1104" points="620" swimtime="00:00:24.51" resultid="3479" heatid="5127" lane="3" />
                <RESULT eventid="1135" points="650" swimtime="00:00:57.07" resultid="3480" heatid="5176" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="652" swimtime="00:00:59.50" resultid="3481" heatid="5263" lane="5" entrytime="00:00:59.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 10.2 - Não completou a distância total da prova.  (Horário: 17:51)" eventid="1213" status="DSQ" swimtime="00:00:00.00" resultid="3482" heatid="5288" lane="3" entrytime="00:00:28.12" entrycourse="LCM" />
                <RESULT eventid="1267" points="621" swimtime="00:00:26.10" resultid="3483" heatid="5329" lane="4" />
                <RESULT eventid="1277" points="612" swimtime="00:02:11.79" resultid="3484" heatid="5348" lane="5" entrytime="00:02:10.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.25" />
                    <SPLIT distance="100" swimtime="00:01:05.46" />
                    <SPLIT distance="150" swimtime="00:01:38.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2383" points="634" swimtime="00:00:24.34" resultid="5984" heatid="6425" lane="7" entrytime="00:00:24.51" />
                <RESULT eventid="2335" points="650" swimtime="00:00:57.06" resultid="6010" heatid="6417" lane="3" entrytime="00:00:57.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2359" points="644" swimtime="00:00:59.73" resultid="6142" heatid="6423" lane="5" entrytime="00:00:59.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcelo" lastname="Vanhazebrouck" birthdate="2010-01-09" gender="M" nation="BRA" license="339043" swrid="5600269" athleteid="3627" externalid="339043">
              <RESULTS>
                <RESULT eventid="1104" points="429" swimtime="00:00:27.72" resultid="3628" heatid="5119" lane="4" entrytime="00:00:27.57" entrycourse="LCM" />
                <RESULT eventid="1135" points="325" swimtime="00:01:11.90" resultid="3629" heatid="5169" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="354" swimtime="00:02:41.13" resultid="3630" heatid="5195" lane="1" entrytime="00:02:41.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.17" />
                    <SPLIT distance="100" swimtime="00:01:18.39" />
                    <SPLIT distance="150" swimtime="00:02:05.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="423" swimtime="00:01:02.42" resultid="3631" heatid="5223" lane="1" entrytime="00:01:00.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="357" swimtime="00:00:31.37" resultid="3632" heatid="5330" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="David Cella" birthdate="2008-02-17" gender="M" nation="BRA" license="341107" swrid="5634581" athleteid="3934" externalid="341107">
              <RESULTS>
                <RESULT eventid="1104" points="587" swimtime="00:00:24.97" resultid="3935" heatid="5126" lane="4" entrytime="00:00:24.16" entrycourse="LCM" />
                <RESULT eventid="1182" points="497" swimtime="00:01:05.12" resultid="3936" heatid="5261" lane="2" entrytime="00:01:04.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="656" swimtime="00:00:53.91" resultid="3937" heatid="5230" lane="5" entrytime="00:00:53.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="516" swimtime="00:00:27.76" resultid="3938" heatid="5329" lane="2" />
                <RESULT eventid="1297" points="583" swimtime="00:00:31.05" resultid="3939" heatid="5371" lane="3" entrytime="00:00:30.69" entrycourse="LCM" />
                <RESULT eventid="2351" points="631" swimtime="00:00:54.61" resultid="6123" heatid="6422" lane="8" entrytime="00:00:53.91">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Vieira Motta" birthdate="2009-09-19" gender="M" nation="BRA" license="339064" swrid="5600271" athleteid="3616" externalid="339064">
              <RESULTS>
                <RESULT eventid="1072" points="538" swimtime="00:04:30.47" resultid="3617" heatid="5061" lane="5" entrytime="00:04:36.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.68" />
                    <SPLIT distance="100" swimtime="00:01:04.13" />
                    <SPLIT distance="150" swimtime="00:01:38.05" />
                    <SPLIT distance="200" swimtime="00:02:12.09" />
                    <SPLIT distance="250" swimtime="00:02:46.65" />
                    <SPLIT distance="300" swimtime="00:03:21.28" />
                    <SPLIT distance="350" swimtime="00:03:56.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="491" swimtime="00:02:09.21" resultid="3618" heatid="5154" lane="7" entrytime="00:02:19.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                    <SPLIT distance="100" swimtime="00:01:02.50" />
                    <SPLIT distance="150" swimtime="00:01:36.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="500" swimtime="00:01:05.01" resultid="3619" heatid="5261" lane="7" entrytime="00:01:05.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="510" swimtime="00:09:25.67" resultid="3620" heatid="5300" lane="8" entrytime="00:09:36.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:06.40" />
                    <SPLIT distance="150" swimtime="00:01:41.42" />
                    <SPLIT distance="200" swimtime="00:02:16.80" />
                    <SPLIT distance="250" swimtime="00:02:52.28" />
                    <SPLIT distance="300" swimtime="00:03:27.84" />
                    <SPLIT distance="350" swimtime="00:04:03.46" />
                    <SPLIT distance="400" swimtime="00:04:39.78" />
                    <SPLIT distance="450" swimtime="00:05:15.34" />
                    <SPLIT distance="500" swimtime="00:05:51.55" />
                    <SPLIT distance="550" swimtime="00:06:27.94" />
                    <SPLIT distance="600" swimtime="00:07:04.26" />
                    <SPLIT distance="650" swimtime="00:07:40.16" />
                    <SPLIT distance="700" swimtime="00:08:16.34" />
                    <SPLIT distance="750" swimtime="00:08:51.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="507" swimtime="00:18:12.00" resultid="3621" heatid="5380" lane="6" entrytime="00:18:04.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.11" />
                    <SPLIT distance="100" swimtime="00:01:06.25" />
                    <SPLIT distance="150" swimtime="00:01:41.33" />
                    <SPLIT distance="200" swimtime="00:02:17.44" />
                    <SPLIT distance="250" swimtime="00:02:53.30" />
                    <SPLIT distance="300" swimtime="00:03:29.90" />
                    <SPLIT distance="350" swimtime="00:04:06.56" />
                    <SPLIT distance="400" swimtime="00:04:43.39" />
                    <SPLIT distance="450" swimtime="00:05:19.96" />
                    <SPLIT distance="500" swimtime="00:05:56.90" />
                    <SPLIT distance="550" swimtime="00:06:33.44" />
                    <SPLIT distance="600" swimtime="00:07:10.56" />
                    <SPLIT distance="650" swimtime="00:07:47.27" />
                    <SPLIT distance="700" swimtime="00:08:24.50" />
                    <SPLIT distance="750" swimtime="00:09:01.23" />
                    <SPLIT distance="800" swimtime="00:09:38.02" />
                    <SPLIT distance="850" swimtime="00:10:15.13" />
                    <SPLIT distance="900" swimtime="00:10:51.85" />
                    <SPLIT distance="950" swimtime="00:11:28.81" />
                    <SPLIT distance="1000" swimtime="00:12:06.03" />
                    <SPLIT distance="1050" swimtime="00:12:42.67" />
                    <SPLIT distance="1100" swimtime="00:13:19.33" />
                    <SPLIT distance="1150" swimtime="00:13:56.26" />
                    <SPLIT distance="1200" swimtime="00:14:33.11" />
                    <SPLIT distance="1250" swimtime="00:15:09.63" />
                    <SPLIT distance="1300" swimtime="00:15:46.43" />
                    <SPLIT distance="1350" swimtime="00:16:23.38" />
                    <SPLIT distance="1400" swimtime="00:17:00.30" />
                    <SPLIT distance="1450" swimtime="00:17:36.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2359" swimtime="00:00:00.00" resultid="6452" entrytime="00:01:05.01" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafaela" lastname="Yolanda Ferreira" birthdate="2008-03-17" gender="F" nation="BRA" license="358335" swrid="5600276" athleteid="3845" externalid="358335">
              <RESULTS>
                <RESULT eventid="1080" points="511" swimtime="00:01:20.19" resultid="3846" heatid="5069" lane="6" entrytime="00:01:19.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="469" swimtime="00:02:57.01" resultid="3847" heatid="5314" lane="6" entrytime="00:02:54.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.51" />
                    <SPLIT distance="100" swimtime="00:01:24.37" />
                    <SPLIT distance="150" swimtime="00:02:11.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="471" swimtime="00:00:37.47" resultid="3848" heatid="5377" lane="8" entrytime="00:00:37.44" entrycourse="LCM" />
                <RESULT eventid="2312" points="502" swimtime="00:01:20.65" resultid="5945" heatid="6416" lane="1" entrytime="00:01:20.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.09" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Carneiro Silva" birthdate="2011-02-21" gender="F" nation="BRA" license="390924" swrid="5602522" athleteid="3921" externalid="390924">
              <RESULTS>
                <RESULT eventid="1096" points="430" swimtime="00:00:31.27" resultid="3922" heatid="5098" lane="5" entrytime="00:00:31.94" entrycourse="LCM" />
                <RESULT eventid="1143" points="335" swimtime="00:03:01.44" resultid="3923" heatid="5187" lane="1" entrytime="00:03:05.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                    <SPLIT distance="100" swimtime="00:01:24.67" />
                    <SPLIT distance="150" swimtime="00:02:22.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="367" swimtime="00:01:20.01" resultid="3924" heatid="5243" lane="7" entrytime="00:01:20.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="376" swimtime="00:01:11.63" resultid="3925" heatid="5203" lane="7" entrytime="00:01:10.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="377" swimtime="00:00:37.15" resultid="3926" heatid="5294" lane="2" entrytime="00:00:36.15" entrycourse="LCM" />
                <RESULT eventid="1275" points="381" swimtime="00:02:49.72" resultid="3927" heatid="5341" lane="6" entrytime="00:02:51.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="LIV" lastname="Carvalho" birthdate="2011-09-13" gender="F" nation="BRA" license="366899" swrid="5602524" athleteid="3756" externalid="366899">
              <RESULTS>
                <RESULT eventid="1080" points="313" swimtime="00:01:34.38" resultid="3757" heatid="5066" lane="6" entrytime="00:01:29.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" points="366" swimtime="00:05:28.86" resultid="3758" heatid="5049" lane="7" entrytime="00:05:36.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.66" />
                    <SPLIT distance="100" swimtime="00:01:18.34" />
                    <SPLIT distance="150" swimtime="00:02:00.31" />
                    <SPLIT distance="200" swimtime="00:02:43.64" />
                    <SPLIT distance="250" swimtime="00:03:26.20" />
                    <SPLIT distance="300" swimtime="00:04:08.52" />
                    <SPLIT distance="350" swimtime="00:04:49.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="377" swimtime="00:02:36.10" resultid="3759" heatid="5138" lane="4" entrytime="00:02:41.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.12" />
                    <SPLIT distance="100" swimtime="00:01:15.78" />
                    <SPLIT distance="150" swimtime="00:01:55.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="337" swimtime="00:11:35.97" resultid="3760" heatid="5271" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.75" />
                    <SPLIT distance="100" swimtime="00:01:20.27" />
                    <SPLIT distance="150" swimtime="00:02:02.98" />
                    <SPLIT distance="200" swimtime="00:02:46.02" />
                    <SPLIT distance="250" swimtime="00:03:29.47" />
                    <SPLIT distance="300" swimtime="00:04:13.17" />
                    <SPLIT distance="350" swimtime="00:04:57.41" />
                    <SPLIT distance="400" swimtime="00:05:42.04" />
                    <SPLIT distance="450" swimtime="00:06:25.97" />
                    <SPLIT distance="500" swimtime="00:07:10.75" />
                    <SPLIT distance="550" swimtime="00:07:55.91" />
                    <SPLIT distance="600" swimtime="00:08:40.34" />
                    <SPLIT distance="650" swimtime="00:09:24.59" />
                    <SPLIT distance="700" swimtime="00:10:09.54" />
                    <SPLIT distance="750" swimtime="00:10:53.00" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 9:30)" eventid="1243" status="DSQ" swimtime="00:03:14.51" resultid="3761" heatid="5312" lane="2" entrytime="00:03:11.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.17" />
                    <SPLIT distance="100" swimtime="00:01:32.41" />
                    <SPLIT distance="150" swimtime="00:02:23.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="363" swimtime="00:00:40.85" resultid="3762" heatid="5375" lane="1" entrytime="00:00:43.03" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="De Krinski" birthdate="2007-07-20" gender="M" nation="BRA" license="334494" swrid="5600148" athleteid="3964" externalid="334494">
              <RESULTS>
                <RESULT eventid="1104" points="521" swimtime="00:00:25.98" resultid="3965" heatid="5129" lane="1" entrytime="00:00:25.85" entrycourse="LCM" />
                <RESULT eventid="1120" points="536" swimtime="00:02:05.49" resultid="3966" heatid="5157" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                    <SPLIT distance="100" swimtime="00:01:00.74" />
                    <SPLIT distance="150" swimtime="00:01:33.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="534" swimtime="00:01:03.57" resultid="3967" heatid="5263" lane="3" entrytime="00:01:01.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="552" swimtime="00:00:28.70" resultid="3968" heatid="5288" lane="6" entrytime="00:00:28.56" entrycourse="LCM" />
                <RESULT eventid="2359" points="527" swimtime="00:01:03.86" resultid="6149" heatid="6423" lane="1" entrytime="00:01:03.57">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Iglesias Vargas" birthdate="2009-01-11" gender="M" nation="BRA" license="324792" swrid="5600189" athleteid="3539" externalid="324792">
              <RESULTS>
                <RESULT eventid="1072" points="581" swimtime="00:04:23.61" resultid="3540" heatid="5062" lane="3" entrytime="00:04:23.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.47" />
                    <SPLIT distance="100" swimtime="00:01:03.59" />
                    <SPLIT distance="150" swimtime="00:01:36.43" />
                    <SPLIT distance="200" swimtime="00:02:09.57" />
                    <SPLIT distance="250" swimtime="00:02:42.71" />
                    <SPLIT distance="300" swimtime="00:03:16.37" />
                    <SPLIT distance="350" swimtime="00:03:50.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="595" swimtime="00:02:01.27" resultid="3541" heatid="5156" lane="3" entrytime="00:02:02.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                    <SPLIT distance="100" swimtime="00:00:59.09" />
                    <SPLIT distance="150" swimtime="00:01:30.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="572" swimtime="00:00:56.42" resultid="3542" heatid="5229" lane="3" entrytime="00:00:57.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="532" swimtime="00:09:17.89" resultid="3543" heatid="5300" lane="6" entrytime="00:09:11.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.09" />
                    <SPLIT distance="100" swimtime="00:01:04.82" />
                    <SPLIT distance="150" swimtime="00:01:39.81" />
                    <SPLIT distance="200" swimtime="00:02:14.77" />
                    <SPLIT distance="250" swimtime="00:02:50.41" />
                    <SPLIT distance="300" swimtime="00:03:25.92" />
                    <SPLIT distance="350" swimtime="00:04:01.32" />
                    <SPLIT distance="400" swimtime="00:04:36.88" />
                    <SPLIT distance="450" swimtime="00:05:12.06" />
                    <SPLIT distance="500" swimtime="00:05:47.81" />
                    <SPLIT distance="550" swimtime="00:06:23.26" />
                    <SPLIT distance="600" swimtime="00:06:58.64" />
                    <SPLIT distance="650" swimtime="00:07:33.79" />
                    <SPLIT distance="700" swimtime="00:08:09.07" />
                    <SPLIT distance="750" swimtime="00:08:44.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="478" swimtime="00:00:28.47" resultid="3544" heatid="5328" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Olivia" lastname="Jeger" birthdate="2004-12-19" gender="F" nation="BRA" license="325493" swrid="5600193" athleteid="3914" externalid="325493" level="UNIDOMBOSC">
              <RESULTS>
                <RESULT eventid="1064" points="597" swimtime="00:04:39.45" resultid="3915" heatid="5055" lane="3" entrytime="00:04:38.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.18" />
                    <SPLIT distance="100" swimtime="00:01:06.59" />
                    <SPLIT distance="150" swimtime="00:01:41.87" />
                    <SPLIT distance="200" swimtime="00:02:17.36" />
                    <SPLIT distance="250" swimtime="00:02:52.99" />
                    <SPLIT distance="300" swimtime="00:03:28.76" />
                    <SPLIT distance="350" swimtime="00:04:04.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="591" swimtime="00:02:14.47" resultid="3916" heatid="5146" lane="6" entrytime="00:02:14.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.69" />
                    <SPLIT distance="100" swimtime="00:01:05.51" />
                    <SPLIT distance="150" swimtime="00:01:40.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="599" swimtime="00:09:34.94" resultid="3917" heatid="5273" lane="5" entrytime="00:09:34.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                    <SPLIT distance="100" swimtime="00:01:08.04" />
                    <SPLIT distance="150" swimtime="00:01:44.11" />
                    <SPLIT distance="200" swimtime="00:02:20.17" />
                    <SPLIT distance="250" swimtime="00:02:56.76" />
                    <SPLIT distance="300" swimtime="00:03:33.33" />
                    <SPLIT distance="350" swimtime="00:04:10.05" />
                    <SPLIT distance="400" swimtime="00:04:46.61" />
                    <SPLIT distance="450" swimtime="00:05:23.12" />
                    <SPLIT distance="500" swimtime="00:05:59.28" />
                    <SPLIT distance="550" swimtime="00:06:35.51" />
                    <SPLIT distance="600" swimtime="00:07:11.56" />
                    <SPLIT distance="650" swimtime="00:07:47.80" />
                    <SPLIT distance="700" swimtime="00:08:24.06" />
                    <SPLIT distance="750" swimtime="00:08:59.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="574" swimtime="00:05:19.82" resultid="3918" heatid="5280" lane="3" entrytime="00:05:20.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:10.78" />
                    <SPLIT distance="150" swimtime="00:01:54.73" />
                    <SPLIT distance="200" swimtime="00:02:36.32" />
                    <SPLIT distance="250" swimtime="00:03:23.93" />
                    <SPLIT distance="300" swimtime="00:04:09.56" />
                    <SPLIT distance="350" swimtime="00:04:45.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1279" points="595" swimtime="00:18:14.00" resultid="3919" heatid="5350" lane="5" entrytime="00:18:04.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                    <SPLIT distance="100" swimtime="00:01:08.55" />
                    <SPLIT distance="150" swimtime="00:01:44.63" />
                    <SPLIT distance="200" swimtime="00:02:20.91" />
                    <SPLIT distance="250" swimtime="00:02:57.57" />
                    <SPLIT distance="300" swimtime="00:03:34.03" />
                    <SPLIT distance="350" swimtime="00:04:10.93" />
                    <SPLIT distance="400" swimtime="00:04:47.67" />
                    <SPLIT distance="450" swimtime="00:05:24.53" />
                    <SPLIT distance="500" swimtime="00:06:01.58" />
                    <SPLIT distance="550" swimtime="00:06:38.17" />
                    <SPLIT distance="600" swimtime="00:07:14.72" />
                    <SPLIT distance="650" swimtime="00:07:51.54" />
                    <SPLIT distance="700" swimtime="00:08:28.35" />
                    <SPLIT distance="750" swimtime="00:09:04.94" />
                    <SPLIT distance="800" swimtime="00:09:41.67" />
                    <SPLIT distance="850" swimtime="00:10:18.04" />
                    <SPLIT distance="900" swimtime="00:10:54.89" />
                    <SPLIT distance="950" swimtime="00:11:31.40" />
                    <SPLIT distance="1000" swimtime="00:12:08.15" />
                    <SPLIT distance="1050" swimtime="00:12:44.62" />
                    <SPLIT distance="1100" swimtime="00:13:21.41" />
                    <SPLIT distance="1150" swimtime="00:13:58.13" />
                    <SPLIT distance="1200" swimtime="00:14:34.87" />
                    <SPLIT distance="1250" swimtime="00:15:11.82" />
                    <SPLIT distance="1300" swimtime="00:15:48.48" />
                    <SPLIT distance="1350" swimtime="00:16:25.24" />
                    <SPLIT distance="1400" swimtime="00:17:02.08" />
                    <SPLIT distance="1450" swimtime="00:17:38.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1295" points="487" swimtime="00:02:34.76" resultid="3920" heatid="5362" lane="3" entrytime="00:02:31.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.86" />
                    <SPLIT distance="100" swimtime="00:01:12.07" />
                    <SPLIT distance="150" swimtime="00:01:53.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ferreira Motta" birthdate="2008-10-24" gender="M" nation="BRA" license="378068" swrid="5600160" athleteid="3867" externalid="378068">
              <RESULTS>
                <RESULT eventid="1088" points="426" swimtime="00:01:15.58" resultid="3868" heatid="5084" lane="4" entrytime="00:01:14.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="390" swimtime="00:02:35.93" resultid="3869" heatid="5196" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:15.11" />
                    <SPLIT distance="150" swimtime="00:01:59.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="349" swimtime="00:01:13.25" resultid="3870" heatid="5259" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="429" swimtime="00:02:46.35" resultid="3871" heatid="5318" lane="4" entrytime="00:02:44.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.91" />
                    <SPLIT distance="100" swimtime="00:01:20.15" />
                    <SPLIT distance="150" swimtime="00:02:03.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="424" swimtime="00:00:34.54" resultid="3872" heatid="5369" lane="7" entrytime="00:00:35.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Presiazniuk" birthdate="2010-10-14" gender="M" nation="BRA" license="356353" swrid="5600237" athleteid="3671" externalid="356353">
              <RESULTS>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 12:21)" eventid="1104" status="DSQ" swimtime="00:00:27.44" resultid="3672" heatid="5120" lane="1" entrytime="00:00:27.51" entrycourse="LCM" />
                <RESULT eventid="1120" points="490" swimtime="00:02:09.34" resultid="3673" heatid="5152" lane="2" entrytime="00:02:11.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.91" />
                    <SPLIT distance="100" swimtime="00:01:03.13" />
                    <SPLIT distance="150" swimtime="00:01:36.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="416" swimtime="00:01:09.10" resultid="3674" heatid="5258" lane="2" entrytime="00:01:08.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="495" swimtime="00:00:59.20" resultid="3675" heatid="5223" lane="7" entrytime="00:00:59.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="412" swimtime="00:00:31.64" resultid="3676" heatid="5282" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Albuquerque" birthdate="2008-03-14" gender="F" nation="BRA" license="324787" swrid="5315259" athleteid="3457" externalid="324787">
              <RESULTS>
                <RESULT eventid="1080" points="578" swimtime="00:01:16.97" resultid="3458" heatid="5069" lane="4" entrytime="00:01:16.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" status="DNS" swimtime="00:00:00.00" resultid="3459" heatid="5208" lane="3" entrytime="00:01:01.87" entrycourse="LCM" />
                <RESULT eventid="1243" points="494" swimtime="00:02:53.96" resultid="3460" heatid="5314" lane="3" entrytime="00:02:47.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.37" />
                    <SPLIT distance="100" swimtime="00:01:21.62" />
                    <SPLIT distance="150" swimtime="00:02:08.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2312" points="562" swimtime="00:01:17.68" resultid="5939" heatid="6416" lane="5" entrytime="00:01:16.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Fontes Hoshina" birthdate="2008-02-15" gender="M" nation="BRA" license="369445" swrid="5600165" athleteid="3502" externalid="369445">
              <RESULTS>
                <RESULT eventid="1135" points="597" swimtime="00:00:58.71" resultid="3503" heatid="5175" lane="3" entrytime="00:00:58.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="570" swimtime="00:00:56.49" resultid="3504" heatid="5230" lane="7" entrytime="00:00:55.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="538" swimtime="00:00:27.38" resultid="3505" heatid="5337" lane="6" entrytime="00:00:27.10" entrycourse="LCM" />
                <RESULT eventid="2335" points="511" swimtime="00:01:01.83" resultid="6014" heatid="6417" lane="1" entrytime="00:00:58.71">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="Heloisa Souza" birthdate="2007-01-15" gender="F" nation="BRA" license="336615" swrid="5600184" athleteid="3545" externalid="336615">
              <RESULTS>
                <RESULT eventid="1064" points="527" swimtime="00:04:51.31" resultid="3546" heatid="5055" lane="5" entrytime="00:04:34.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.03" />
                    <SPLIT distance="100" swimtime="00:01:09.46" />
                    <SPLIT distance="150" swimtime="00:01:46.34" />
                    <SPLIT distance="200" swimtime="00:02:23.51" />
                    <SPLIT distance="250" swimtime="00:03:01.23" />
                    <SPLIT distance="300" swimtime="00:03:38.47" />
                    <SPLIT distance="350" swimtime="00:04:15.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="556" swimtime="00:02:17.18" resultid="3547" heatid="5146" lane="5" entrytime="00:02:08.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:06.25" />
                    <SPLIT distance="150" swimtime="00:01:42.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="544" swimtime="00:01:03.34" resultid="3548" heatid="5209" lane="4" entrytime="00:00:59.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="551" swimtime="00:09:51.30" resultid="3549" heatid="5273" lane="3" entrytime="00:09:41.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.87" />
                    <SPLIT distance="100" swimtime="00:01:09.93" />
                    <SPLIT distance="150" swimtime="00:01:46.88" />
                    <SPLIT distance="200" swimtime="00:02:23.39" />
                    <SPLIT distance="250" swimtime="00:03:00.74" />
                    <SPLIT distance="300" swimtime="00:03:38.06" />
                    <SPLIT distance="350" swimtime="00:04:15.34" />
                    <SPLIT distance="400" swimtime="00:04:52.77" />
                    <SPLIT distance="450" swimtime="00:05:30.20" />
                    <SPLIT distance="500" swimtime="00:06:07.46" />
                    <SPLIT distance="550" swimtime="00:06:45.04" />
                    <SPLIT distance="600" swimtime="00:07:22.45" />
                    <SPLIT distance="650" swimtime="00:08:00.09" />
                    <SPLIT distance="700" swimtime="00:08:37.41" />
                    <SPLIT distance="750" swimtime="00:09:14.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1279" points="538" swimtime="00:18:51.25" resultid="3550" heatid="5349" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                    <SPLIT distance="100" swimtime="00:01:11.06" />
                    <SPLIT distance="150" swimtime="00:01:48.56" />
                    <SPLIT distance="200" swimtime="00:02:26.18" />
                    <SPLIT distance="250" swimtime="00:03:04.45" />
                    <SPLIT distance="300" swimtime="00:03:42.27" />
                    <SPLIT distance="350" swimtime="00:04:20.30" />
                    <SPLIT distance="400" swimtime="00:04:58.74" />
                    <SPLIT distance="450" swimtime="00:05:36.73" />
                    <SPLIT distance="500" swimtime="00:06:14.31" />
                    <SPLIT distance="550" swimtime="00:06:52.27" />
                    <SPLIT distance="600" swimtime="00:07:30.17" />
                    <SPLIT distance="650" swimtime="00:08:08.50" />
                    <SPLIT distance="700" swimtime="00:08:46.66" />
                    <SPLIT distance="750" swimtime="00:09:24.87" />
                    <SPLIT distance="800" swimtime="00:10:03.15" />
                    <SPLIT distance="850" swimtime="00:10:41.25" />
                    <SPLIT distance="900" swimtime="00:11:19.46" />
                    <SPLIT distance="950" swimtime="00:11:57.51" />
                    <SPLIT distance="1000" swimtime="00:12:35.73" />
                    <SPLIT distance="1050" swimtime="00:13:13.57" />
                    <SPLIT distance="1100" swimtime="00:13:51.45" />
                    <SPLIT distance="1150" swimtime="00:14:28.94" />
                    <SPLIT distance="1200" swimtime="00:15:06.82" />
                    <SPLIT distance="1250" swimtime="00:15:44.52" />
                    <SPLIT distance="1300" swimtime="00:16:22.13" />
                    <SPLIT distance="1350" swimtime="00:16:59.54" />
                    <SPLIT distance="1400" swimtime="00:17:36.91" />
                    <SPLIT distance="1450" swimtime="00:18:14.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2343" points="588" swimtime="00:01:01.69" resultid="6107" heatid="6421" lane="1" entrytime="00:01:03.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Martinez Diniz" birthdate="2008-11-22" gender="M" nation="BRA" license="339400" swrid="5717283" athleteid="3580" externalid="339400">
              <RESULTS>
                <RESULT eventid="1104" points="509" swimtime="00:00:26.18" resultid="3581" heatid="5125" lane="1" entrytime="00:00:26.35" entrycourse="LCM" />
                <RESULT eventid="1120" points="482" swimtime="00:02:10.03" resultid="3582" heatid="5155" lane="2" entrytime="00:02:11.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                    <SPLIT distance="100" swimtime="00:01:04.16" />
                    <SPLIT distance="150" swimtime="00:01:37.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="564" swimtime="00:00:56.70" resultid="3583" heatid="5229" lane="4" entrytime="00:00:56.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophie" lastname="Kraemer Geremia" birthdate="2011-07-20" gender="F" nation="BRA" license="366908" swrid="5588763" athleteid="3795" externalid="366908">
              <RESULTS>
                <RESULT eventid="1064" points="451" swimtime="00:05:06.81" resultid="3796" heatid="5051" lane="2" entrytime="00:05:04.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.45" />
                    <SPLIT distance="100" swimtime="00:01:13.38" />
                    <SPLIT distance="150" swimtime="00:01:53.42" />
                    <SPLIT distance="200" swimtime="00:02:32.73" />
                    <SPLIT distance="250" swimtime="00:03:12.50" />
                    <SPLIT distance="300" swimtime="00:03:51.09" />
                    <SPLIT distance="350" swimtime="00:04:29.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="499" swimtime="00:02:22.21" resultid="3797" heatid="5141" lane="6" entrytime="00:02:22.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                    <SPLIT distance="100" swimtime="00:01:08.99" />
                    <SPLIT distance="150" swimtime="00:01:46.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="442" swimtime="00:01:15.24" resultid="3798" heatid="5244" lane="5" entrytime="00:01:13.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="394" swimtime="00:11:00.90" resultid="3799" heatid="5271" lane="3" entrytime="00:10:28.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.90" />
                    <SPLIT distance="100" swimtime="00:01:17.71" />
                    <SPLIT distance="150" swimtime="00:02:00.04" />
                    <SPLIT distance="200" swimtime="00:02:41.80" />
                    <SPLIT distance="250" swimtime="00:03:24.26" />
                    <SPLIT distance="300" swimtime="00:04:06.28" />
                    <SPLIT distance="350" swimtime="00:04:48.25" />
                    <SPLIT distance="400" swimtime="00:05:30.41" />
                    <SPLIT distance="450" swimtime="00:06:13.00" />
                    <SPLIT distance="500" swimtime="00:06:54.68" />
                    <SPLIT distance="550" swimtime="00:07:36.79" />
                    <SPLIT distance="600" swimtime="00:08:18.20" />
                    <SPLIT distance="650" swimtime="00:08:59.57" />
                    <SPLIT distance="700" swimtime="00:09:40.59" />
                    <SPLIT distance="750" swimtime="00:10:21.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1275" points="434" swimtime="00:02:42.62" resultid="3800" heatid="5343" lane="2" entrytime="00:02:39.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.24" />
                    <SPLIT distance="100" swimtime="00:01:20.20" />
                    <SPLIT distance="150" swimtime="00:02:01.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2391" points="421" swimtime="00:01:16.48" resultid="6135" heatid="6424" lane="8" entrytime="00:01:15.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Fontoura" birthdate="2010-08-26" gender="M" nation="BRA" license="338922" swrid="5600167" athleteid="3703" externalid="338922">
              <RESULTS>
                <RESULT eventid="1072" points="376" swimtime="00:05:04.71" resultid="3704" heatid="5057" lane="4" entrytime="00:05:11.17" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.14" />
                    <SPLIT distance="100" swimtime="00:01:13.20" />
                    <SPLIT distance="150" swimtime="00:01:53.25" />
                    <SPLIT distance="200" swimtime="00:02:33.12" />
                    <SPLIT distance="250" swimtime="00:03:12.69" />
                    <SPLIT distance="300" swimtime="00:03:51.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="379" swimtime="00:00:28.88" resultid="3705" heatid="5118" lane="3" entrytime="00:00:29.09" entrycourse="LCM" />
                <RESULT eventid="1120" points="371" swimtime="00:02:21.90" resultid="3706" heatid="5148" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.96" />
                    <SPLIT distance="100" swimtime="00:01:08.19" />
                    <SPLIT distance="150" swimtime="00:01:45.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="331" swimtime="00:02:44.64" resultid="3707" heatid="5194" lane="6" entrytime="00:02:44.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.82" />
                    <SPLIT distance="100" swimtime="00:01:18.91" />
                    <SPLIT distance="150" swimtime="00:02:10.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="405" swimtime="00:01:03.31" resultid="3708" heatid="5222" lane="8" entrytime="00:01:03.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="314" swimtime="00:00:32.75" resultid="3709" heatid="5330" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giulia" lastname="Salesi Chicon" birthdate="2002-04-16" gender="F" nation="BRA" license="250865" swrid="5600255" athleteid="3902" externalid="250865">
              <RESULTS>
                <RESULT eventid="1064" points="677" swimtime="00:04:27.95" resultid="3903" heatid="5055" lane="4" entrytime="00:04:17.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:03.05" />
                    <SPLIT distance="150" swimtime="00:01:36.44" />
                    <SPLIT distance="200" swimtime="00:02:10.38" />
                    <SPLIT distance="250" swimtime="00:02:44.81" />
                    <SPLIT distance="300" swimtime="00:03:19.35" />
                    <SPLIT distance="350" swimtime="00:03:54.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="727" swimtime="00:02:05.49" resultid="3904" heatid="5146" lane="4" entrytime="00:02:03.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.12" />
                    <SPLIT distance="100" swimtime="00:01:00.32" />
                    <SPLIT distance="150" swimtime="00:01:32.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="609" swimtime="00:02:28.78" resultid="3905" heatid="5191" lane="4" entrytime="00:02:28.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.68" />
                    <SPLIT distance="100" swimtime="00:01:12.26" />
                    <SPLIT distance="150" swimtime="00:01:56.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="690" swimtime="00:09:08.49" resultid="3906" heatid="5273" lane="4" entrytime="00:08:58.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                    <SPLIT distance="100" swimtime="00:01:05.59" />
                    <SPLIT distance="150" swimtime="00:01:40.20" />
                    <SPLIT distance="200" swimtime="00:02:14.74" />
                    <SPLIT distance="250" swimtime="00:02:49.61" />
                    <SPLIT distance="300" swimtime="00:03:24.16" />
                    <SPLIT distance="350" swimtime="00:03:58.99" />
                    <SPLIT distance="400" swimtime="00:04:33.73" />
                    <SPLIT distance="450" swimtime="00:05:08.37" />
                    <SPLIT distance="500" swimtime="00:05:42.96" />
                    <SPLIT distance="550" swimtime="00:06:17.23" />
                    <SPLIT distance="600" swimtime="00:06:51.44" />
                    <SPLIT distance="650" swimtime="00:07:25.82" />
                    <SPLIT distance="700" swimtime="00:08:00.51" />
                    <SPLIT distance="750" swimtime="00:08:34.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="590" swimtime="00:05:16.94" resultid="3907" heatid="5280" lane="4" entrytime="00:05:10.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                    <SPLIT distance="100" swimtime="00:01:11.22" />
                    <SPLIT distance="150" swimtime="00:01:53.48" />
                    <SPLIT distance="200" swimtime="00:02:35.08" />
                    <SPLIT distance="250" swimtime="00:03:21.51" />
                    <SPLIT distance="300" swimtime="00:04:07.39" />
                    <SPLIT distance="350" swimtime="00:04:42.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1279" points="635" swimtime="00:17:50.78" resultid="3908" heatid="5350" lane="4" entrytime="00:17:07.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.74" />
                    <SPLIT distance="100" swimtime="00:01:07.26" />
                    <SPLIT distance="150" swimtime="00:01:42.81" />
                    <SPLIT distance="200" swimtime="00:02:18.09" />
                    <SPLIT distance="250" swimtime="00:02:54.06" />
                    <SPLIT distance="300" swimtime="00:03:29.83" />
                    <SPLIT distance="350" swimtime="00:04:05.69" />
                    <SPLIT distance="400" swimtime="00:04:41.55" />
                    <SPLIT distance="450" swimtime="00:05:17.62" />
                    <SPLIT distance="500" swimtime="00:05:53.34" />
                    <SPLIT distance="550" swimtime="00:06:29.20" />
                    <SPLIT distance="600" swimtime="00:07:04.91" />
                    <SPLIT distance="650" swimtime="00:07:41.08" />
                    <SPLIT distance="700" swimtime="00:08:16.88" />
                    <SPLIT distance="750" swimtime="00:08:52.87" />
                    <SPLIT distance="800" swimtime="00:09:28.97" />
                    <SPLIT distance="850" swimtime="00:10:05.21" />
                    <SPLIT distance="900" swimtime="00:10:41.26" />
                    <SPLIT distance="950" swimtime="00:11:17.12" />
                    <SPLIT distance="1000" swimtime="00:11:52.83" />
                    <SPLIT distance="1050" swimtime="00:12:28.37" />
                    <SPLIT distance="1100" swimtime="00:13:04.09" />
                    <SPLIT distance="1150" swimtime="00:13:39.75" />
                    <SPLIT distance="1200" swimtime="00:14:15.79" />
                    <SPLIT distance="1250" swimtime="00:14:51.58" />
                    <SPLIT distance="1300" swimtime="00:15:27.43" />
                    <SPLIT distance="1350" swimtime="00:16:03.73" />
                    <SPLIT distance="1400" swimtime="00:16:40.01" />
                    <SPLIT distance="1450" swimtime="00:17:15.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ricardo" lastname="De Lima Cavalcanti" birthdate="2009-12-17" gender="M" nation="BRA" license="380965" swrid="5634589" athleteid="3945" externalid="380965">
              <RESULTS>
                <RESULT eventid="1104" points="528" swimtime="00:00:25.86" resultid="3946" heatid="5126" lane="7" entrytime="00:00:25.20" entrycourse="LCM" />
                <RESULT eventid="1135" points="560" swimtime="00:00:59.99" resultid="3947" heatid="5175" lane="7" entrytime="00:01:01.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="544" swimtime="00:00:57.38" resultid="3948" heatid="5229" lane="8" entrytime="00:00:57.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="529" swimtime="00:00:27.52" resultid="3949" heatid="5336" lane="2" entrytime="00:00:27.72" entrycourse="LCM" />
                <RESULT eventid="1293" points="453" swimtime="00:02:23.63" resultid="3950" heatid="5360" lane="1" entrytime="00:02:22.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                    <SPLIT distance="100" swimtime="00:01:07.30" />
                    <SPLIT distance="150" swimtime="00:01:46.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helen" lastname="Barato Bernardi" birthdate="2006-07-27" gender="F" nation="BRA" license="317031" swrid="5717244" athleteid="3951" externalid="317031">
              <RESULTS>
                <RESULT eventid="1080" points="639" swimtime="00:01:14.44" resultid="3952" heatid="5070" lane="4" entrytime="00:01:13.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="491" swimtime="00:00:29.92" resultid="3953" heatid="5106" lane="3" entrytime="00:00:29.32" entrycourse="LCM" />
                <RESULT eventid="1143" points="446" swimtime="00:02:45.06" resultid="3954" heatid="5191" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                    <SPLIT distance="100" swimtime="00:01:21.45" />
                    <SPLIT distance="150" swimtime="00:02:07.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="388" swimtime="00:00:33.47" resultid="3955" heatid="5322" lane="5" />
                <RESULT eventid="1243" points="574" swimtime="00:02:45.50" resultid="3956" heatid="5314" lane="4" entrytime="00:02:41.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.71" />
                    <SPLIT distance="100" swimtime="00:01:20.58" />
                    <SPLIT distance="150" swimtime="00:02:03.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="616" swimtime="00:00:34.27" resultid="3957" heatid="5377" lane="4" entrytime="00:00:33.35" entrycourse="LCM" />
                <RESULT eventid="2312" points="629" swimtime="00:01:14.84" resultid="5938" heatid="6416" lane="4" entrytime="00:01:14.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Muxfeldt" birthdate="2011-05-13" gender="F" nation="BRA" license="366903" swrid="5602563" athleteid="3770" externalid="366903">
              <RESULTS>
                <RESULT eventid="1080" points="421" swimtime="00:01:25.54" resultid="3771" heatid="5067" lane="8" entrytime="00:01:25.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="428" swimtime="00:00:31.31" resultid="3772" heatid="5099" lane="5" entrytime="00:00:30.86" entrycourse="LCM" />
                <RESULT eventid="1112" points="450" swimtime="00:02:27.24" resultid="3773" heatid="5140" lane="5" entrytime="00:02:26.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:01:12.48" />
                    <SPLIT distance="150" swimtime="00:01:51.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="401" swimtime="00:03:06.44" resultid="3774" heatid="5312" lane="4" entrytime="00:03:04.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                    <SPLIT distance="100" swimtime="00:01:30.48" />
                    <SPLIT distance="150" swimtime="00:02:20.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1279" points="398" swimtime="00:20:50.92" resultid="3775" heatid="5349" lane="6" entrytime="00:21:41.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                    <SPLIT distance="100" swimtime="00:01:18.75" />
                    <SPLIT distance="150" swimtime="00:02:01.41" />
                    <SPLIT distance="200" swimtime="00:02:44.03" />
                    <SPLIT distance="250" swimtime="00:03:26.66" />
                    <SPLIT distance="300" swimtime="00:04:09.63" />
                    <SPLIT distance="350" swimtime="00:04:52.02" />
                    <SPLIT distance="400" swimtime="00:05:34.38" />
                    <SPLIT distance="450" swimtime="00:06:18.26" />
                    <SPLIT distance="500" swimtime="00:07:01.07" />
                    <SPLIT distance="550" swimtime="00:07:43.32" />
                    <SPLIT distance="600" swimtime="00:08:25.70" />
                    <SPLIT distance="650" swimtime="00:09:07.42" />
                    <SPLIT distance="700" swimtime="00:09:49.21" />
                    <SPLIT distance="750" swimtime="00:10:30.78" />
                    <SPLIT distance="800" swimtime="00:11:12.90" />
                    <SPLIT distance="850" swimtime="00:11:54.07" />
                    <SPLIT distance="900" swimtime="00:12:35.53" />
                    <SPLIT distance="950" swimtime="00:13:17.21" />
                    <SPLIT distance="1000" swimtime="00:13:58.03" />
                    <SPLIT distance="1050" swimtime="00:14:39.11" />
                    <SPLIT distance="1100" swimtime="00:15:20.84" />
                    <SPLIT distance="1150" swimtime="00:16:02.03" />
                    <SPLIT distance="1200" swimtime="00:16:43.64" />
                    <SPLIT distance="1250" swimtime="00:17:25.09" />
                    <SPLIT distance="1300" swimtime="00:18:07.13" />
                    <SPLIT distance="1350" swimtime="00:18:48.76" />
                    <SPLIT distance="1400" swimtime="00:19:30.55" />
                    <SPLIT distance="1450" swimtime="00:20:12.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="366" swimtime="00:00:40.75" resultid="3776" heatid="5375" lane="3" entrytime="00:00:40.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Cabrera Cirino" birthdate="2011-01-28" gender="M" nation="BRA" license="369531" swrid="5588569" athleteid="3825" externalid="369531">
              <RESULTS>
                <RESULT eventid="1072" points="473" swimtime="00:04:42.35" resultid="3826" heatid="5059" lane="7" entrytime="00:04:45.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.55" />
                    <SPLIT distance="100" swimtime="00:01:04.96" />
                    <SPLIT distance="150" swimtime="00:01:40.79" />
                    <SPLIT distance="200" swimtime="00:02:16.66" />
                    <SPLIT distance="250" swimtime="00:02:52.75" />
                    <SPLIT distance="300" swimtime="00:03:29.72" />
                    <SPLIT distance="350" swimtime="00:04:06.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="451" swimtime="00:00:27.26" resultid="3827" heatid="5120" lane="2" entrytime="00:00:27.00" entrycourse="LCM" />
                <RESULT eventid="1120" points="450" swimtime="00:02:13.01" resultid="3828" heatid="5152" lane="1" entrytime="00:02:12.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.81" />
                    <SPLIT distance="100" swimtime="00:01:03.65" />
                    <SPLIT distance="150" swimtime="00:01:38.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="396" swimtime="00:01:10.21" resultid="3829" heatid="5258" lane="7" entrytime="00:01:08.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="476" swimtime="00:00:59.98" resultid="3830" heatid="5222" lane="4" entrytime="00:01:00.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="437" swimtime="00:02:27.48" resultid="3831" heatid="5347" lane="1" entrytime="00:02:27.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="100" swimtime="00:01:12.28" />
                    <SPLIT distance="150" swimtime="00:01:50.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Vitoria Kuzmann Cercal" birthdate="2009-04-10" gender="F" nation="BRA" license="339082" swrid="5600274" athleteid="3607" externalid="339082">
              <RESULTS>
                <RESULT eventid="1096" points="504" swimtime="00:00:29.66" resultid="3608" heatid="5102" lane="4" entrytime="00:00:30.61" entrycourse="LCM" />
                <RESULT eventid="1128" points="412" swimtime="00:01:14.50" resultid="3609" heatid="5161" lane="6" entrytime="00:01:18.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="426" swimtime="00:01:16.15" resultid="3610" heatid="5247" lane="1" entrytime="00:01:16.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="404" swimtime="00:00:36.32" resultid="3611" heatid="5290" lane="2" />
                <RESULT eventid="1275" status="DNS" swimtime="00:00:00.00" resultid="3612" heatid="5342" lane="2" entrytime="00:02:46.94" entrycourse="LCM" />
                <RESULT eventid="2328" points="373" swimtime="00:01:17.05" resultid="6003" heatid="6418" lane="1" entrytime="00:01:14.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Francisco Saldo" birthdate="2007-01-23" gender="M" nation="BRA" license="313537" swrid="5600169" athleteid="3516" externalid="313537">
              <RESULTS>
                <RESULT eventid="1088" points="482" swimtime="00:01:12.51" resultid="3517" heatid="5087" lane="7" entrytime="00:01:11.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="699" swimtime="00:04:07.95" resultid="3518" heatid="5063" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.18" />
                    <SPLIT distance="100" swimtime="00:01:00.05" />
                    <SPLIT distance="150" swimtime="00:01:32.01" />
                    <SPLIT distance="200" swimtime="00:02:03.81" />
                    <SPLIT distance="250" swimtime="00:02:36.13" />
                    <SPLIT distance="300" swimtime="00:03:07.57" />
                    <SPLIT distance="350" swimtime="00:03:39.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="561" swimtime="00:00:59.94" resultid="3519" heatid="5178" lane="5" entrytime="00:00:56.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="644" swimtime="00:01:58.10" resultid="3520" heatid="5157" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.75" />
                    <SPLIT distance="100" swimtime="00:00:57.80" />
                    <SPLIT distance="150" swimtime="00:01:27.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="617" swimtime="00:04:44.70" resultid="3521" heatid="5277" lane="4" entrytime="00:04:39.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.53" />
                    <SPLIT distance="100" swimtime="00:01:00.71" />
                    <SPLIT distance="150" swimtime="00:01:39.71" />
                    <SPLIT distance="200" swimtime="00:02:18.68" />
                    <SPLIT distance="250" swimtime="00:02:59.37" />
                    <SPLIT distance="300" swimtime="00:03:40.13" />
                    <SPLIT distance="350" swimtime="00:04:12.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1293" points="665" swimtime="00:02:06.38" resultid="3522" heatid="5360" lane="4" entrytime="00:02:02.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.56" />
                    <SPLIT distance="100" swimtime="00:01:00.23" />
                    <SPLIT distance="150" swimtime="00:01:34.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Cristina Ferreira" birthdate="2011-08-24" gender="F" nation="BRA" license="358334" swrid="5588611" athleteid="3849" externalid="358334">
              <RESULTS>
                <RESULT eventid="1064" points="517" swimtime="00:04:53.14" resultid="3850" heatid="5051" lane="4" entrytime="00:04:33.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.17" />
                    <SPLIT distance="100" swimtime="00:01:09.32" />
                    <SPLIT distance="150" swimtime="00:01:46.51" />
                    <SPLIT distance="200" swimtime="00:02:23.57" />
                    <SPLIT distance="250" swimtime="00:03:01.21" />
                    <SPLIT distance="300" swimtime="00:03:38.45" />
                    <SPLIT distance="350" swimtime="00:04:16.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" points="619" swimtime="00:01:05.09" resultid="3851" heatid="5160" lane="4" entrytime="00:01:04.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="533" swimtime="00:02:35.51" resultid="3852" heatid="5188" lane="4" entrytime="00:02:28.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.35" />
                    <SPLIT distance="100" swimtime="00:01:14.90" />
                    <SPLIT distance="150" swimtime="00:02:02.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="535" swimtime="00:05:27.49" resultid="3853" heatid="5280" lane="5" entrytime="00:05:13.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:12.29" />
                    <SPLIT distance="150" swimtime="00:01:56.56" />
                    <SPLIT distance="200" swimtime="00:02:40.60" />
                    <SPLIT distance="250" swimtime="00:03:26.89" />
                    <SPLIT distance="300" swimtime="00:04:12.72" />
                    <SPLIT distance="350" swimtime="00:04:50.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="456" swimtime="00:02:58.66" resultid="3854" heatid="5314" lane="5" entrytime="00:02:45.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.48" />
                    <SPLIT distance="100" swimtime="00:01:25.03" />
                    <SPLIT distance="150" swimtime="00:02:11.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1295" points="503" swimtime="00:02:33.16" resultid="3855" heatid="5362" lane="4" entrytime="00:02:21.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.34" />
                    <SPLIT distance="100" swimtime="00:01:11.96" />
                    <SPLIT distance="150" swimtime="00:01:52.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2328" points="598" swimtime="00:01:05.85" resultid="5997" heatid="6418" lane="4" entrytime="00:01:05.09">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Godino" birthdate="2010-04-27" gender="F" nation="BRA" license="356355" swrid="5600176" athleteid="3684" externalid="356355">
              <RESULTS>
                <RESULT eventid="1064" points="433" swimtime="00:05:11.09" resultid="3685" heatid="5050" lane="2" entrytime="00:05:11.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                    <SPLIT distance="100" swimtime="00:01:13.59" />
                    <SPLIT distance="150" swimtime="00:01:52.85" />
                    <SPLIT distance="200" swimtime="00:02:32.26" />
                    <SPLIT distance="250" swimtime="00:03:11.92" />
                    <SPLIT distance="300" swimtime="00:03:51.79" />
                    <SPLIT distance="350" swimtime="00:04:31.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="443" swimtime="00:02:28.01" resultid="3686" heatid="5140" lane="3" entrytime="00:02:27.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:10.54" />
                    <SPLIT distance="150" swimtime="00:01:49.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="442" swimtime="00:10:36.31" resultid="3687" heatid="5271" lane="2" entrytime="00:10:36.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                    <SPLIT distance="100" swimtime="00:01:14.61" />
                    <SPLIT distance="150" swimtime="00:01:54.05" />
                    <SPLIT distance="200" swimtime="00:02:33.73" />
                    <SPLIT distance="250" swimtime="00:03:14.02" />
                    <SPLIT distance="300" swimtime="00:03:54.48" />
                    <SPLIT distance="350" swimtime="00:04:35.10" />
                    <SPLIT distance="400" swimtime="00:05:15.44" />
                    <SPLIT distance="450" swimtime="00:05:56.13" />
                    <SPLIT distance="500" swimtime="00:06:36.81" />
                    <SPLIT distance="550" swimtime="00:07:17.35" />
                    <SPLIT distance="600" swimtime="00:07:57.68" />
                    <SPLIT distance="650" swimtime="00:08:38.07" />
                    <SPLIT distance="700" swimtime="00:09:18.00" />
                    <SPLIT distance="750" swimtime="00:09:58.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1275" points="335" swimtime="00:02:57.29" resultid="3688" heatid="5341" lane="8" entrytime="00:02:54.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                    <SPLIT distance="100" swimtime="00:01:26.66" />
                    <SPLIT distance="150" swimtime="00:02:12.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1279" points="410" swimtime="00:20:38.09" resultid="3689" heatid="5350" lane="1" entrytime="00:20:37.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                    <SPLIT distance="100" swimtime="00:01:17.49" />
                    <SPLIT distance="150" swimtime="00:01:58.60" />
                    <SPLIT distance="200" swimtime="00:02:39.81" />
                    <SPLIT distance="250" swimtime="00:03:21.70" />
                    <SPLIT distance="300" swimtime="00:04:03.34" />
                    <SPLIT distance="350" swimtime="00:04:45.60" />
                    <SPLIT distance="400" swimtime="00:05:27.65" />
                    <SPLIT distance="450" swimtime="00:06:09.65" />
                    <SPLIT distance="500" swimtime="00:06:51.56" />
                    <SPLIT distance="550" swimtime="00:07:33.50" />
                    <SPLIT distance="600" swimtime="00:08:15.10" />
                    <SPLIT distance="650" swimtime="00:08:57.46" />
                    <SPLIT distance="700" swimtime="00:09:39.20" />
                    <SPLIT distance="750" swimtime="00:10:21.32" />
                    <SPLIT distance="800" swimtime="00:11:02.86" />
                    <SPLIT distance="850" swimtime="00:11:44.80" />
                    <SPLIT distance="900" swimtime="00:12:26.47" />
                    <SPLIT distance="950" swimtime="00:13:08.42" />
                    <SPLIT distance="1000" swimtime="00:13:50.23" />
                    <SPLIT distance="1050" swimtime="00:14:31.57" />
                    <SPLIT distance="1100" swimtime="00:15:13.04" />
                    <SPLIT distance="1150" swimtime="00:15:54.48" />
                    <SPLIT distance="1200" swimtime="00:16:35.62" />
                    <SPLIT distance="1250" swimtime="00:17:16.86" />
                    <SPLIT distance="1300" swimtime="00:17:57.89" />
                    <SPLIT distance="1350" swimtime="00:18:38.52" />
                    <SPLIT distance="1400" swimtime="00:19:19.16" />
                    <SPLIT distance="1450" swimtime="00:19:59.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marina" lastname="De Albuquerque" birthdate="2010-06-08" gender="F" nation="BRA" license="356249" swrid="5600145" athleteid="3639" externalid="356249">
              <RESULTS>
                <RESULT eventid="1096" points="373" swimtime="00:00:32.78" resultid="3640" heatid="5099" lane="8" entrytime="00:00:31.83" entrycourse="LCM" />
                <RESULT eventid="1175" points="392" swimtime="00:01:18.30" resultid="3641" heatid="5244" lane="2" entrytime="00:01:16.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="380" swimtime="00:01:11.35" resultid="3642" heatid="5203" lane="2" entrytime="00:01:10.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="424" swimtime="00:00:35.73" resultid="3643" heatid="5294" lane="5" entrytime="00:00:35.45" entrycourse="LCM" />
                <RESULT eventid="1275" points="399" swimtime="00:02:47.19" resultid="3644" heatid="5343" lane="1" entrytime="00:02:44.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.95" />
                    <SPLIT distance="100" swimtime="00:01:21.94" />
                    <SPLIT distance="150" swimtime="00:02:04.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Kremer De Aguiar" birthdate="2009-12-22" gender="F" nation="BRA" license="338987" swrid="5600196" athleteid="3597" externalid="338987">
              <RESULTS>
                <RESULT eventid="1080" points="448" swimtime="00:01:23.80" resultid="3598" heatid="5068" lane="4" entrytime="00:01:23.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="449" swimtime="00:02:44.69" resultid="3599" heatid="5190" lane="1" entrytime="00:02:45.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.42" />
                    <SPLIT distance="100" swimtime="00:01:19.50" />
                    <SPLIT distance="150" swimtime="00:02:07.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="422" swimtime="00:03:03.35" resultid="3600" heatid="5313" lane="1" entrytime="00:03:02.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.43" />
                    <SPLIT distance="100" swimtime="00:01:26.75" />
                    <SPLIT distance="150" swimtime="00:02:15.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="482" swimtime="00:00:37.18" resultid="3601" heatid="5376" lane="1" entrytime="00:00:39.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Leao" birthdate="2011-09-18" gender="M" nation="BRA" license="366880" swrid="5602553" athleteid="3720" externalid="366880">
              <RESULTS>
                <RESULT eventid="1072" points="392" swimtime="00:05:00.60" resultid="3721" heatid="5059" lane="8" entrytime="00:04:52.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:11.51" />
                    <SPLIT distance="150" swimtime="00:01:49.74" />
                    <SPLIT distance="200" swimtime="00:02:28.32" />
                    <SPLIT distance="250" swimtime="00:03:07.61" />
                    <SPLIT distance="300" swimtime="00:03:45.96" />
                    <SPLIT distance="350" swimtime="00:04:24.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="367" swimtime="00:02:22.41" resultid="3722" heatid="5151" lane="6" entrytime="00:02:19.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.28" />
                    <SPLIT distance="100" swimtime="00:01:08.99" />
                    <SPLIT distance="150" swimtime="00:01:46.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="296" swimtime="00:01:17.40" resultid="3723" heatid="5256" lane="1" entrytime="00:01:23.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="412" swimtime="00:10:07.36" resultid="3724" heatid="5299" lane="2" entrytime="00:10:03.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                    <SPLIT distance="100" swimtime="00:01:10.81" />
                    <SPLIT distance="150" swimtime="00:01:49.82" />
                    <SPLIT distance="200" swimtime="00:02:28.20" />
                    <SPLIT distance="250" swimtime="00:03:07.54" />
                    <SPLIT distance="300" swimtime="00:03:46.02" />
                    <SPLIT distance="350" swimtime="00:04:24.70" />
                    <SPLIT distance="400" swimtime="00:05:02.92" />
                    <SPLIT distance="450" swimtime="00:05:41.65" />
                    <SPLIT distance="500" swimtime="00:06:20.14" />
                    <SPLIT distance="550" swimtime="00:06:58.98" />
                    <SPLIT distance="600" swimtime="00:07:36.96" />
                    <SPLIT distance="650" swimtime="00:08:15.74" />
                    <SPLIT distance="700" swimtime="00:08:53.38" />
                    <SPLIT distance="750" swimtime="00:09:31.65" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 6.4 - Não estava de costas ao sair da parede após a virada.&#10;&#10;&#10;&#10;&#10;&#10;&#10;  (Horário: 11:12), Após a volta dos 150m." eventid="1277" status="DSQ" swimtime="00:02:49.53" resultid="3725" heatid="5344" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.20" />
                    <SPLIT distance="150" swimtime="00:02:08.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="406" swimtime="00:19:35.34" resultid="3726" heatid="5380" lane="8" entrytime="00:19:22.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                    <SPLIT distance="100" swimtime="00:01:13.16" />
                    <SPLIT distance="150" swimtime="00:01:53.08" />
                    <SPLIT distance="200" swimtime="00:02:31.97" />
                    <SPLIT distance="250" swimtime="00:03:11.66" />
                    <SPLIT distance="300" swimtime="00:03:51.42" />
                    <SPLIT distance="350" swimtime="00:04:31.86" />
                    <SPLIT distance="400" swimtime="00:05:10.36" />
                    <SPLIT distance="450" swimtime="00:05:50.53" />
                    <SPLIT distance="500" swimtime="00:06:29.70" />
                    <SPLIT distance="550" swimtime="00:07:10.60" />
                    <SPLIT distance="600" swimtime="00:07:49.28" />
                    <SPLIT distance="650" swimtime="00:08:29.51" />
                    <SPLIT distance="700" swimtime="00:09:08.30" />
                    <SPLIT distance="750" swimtime="00:09:48.53" />
                    <SPLIT distance="800" swimtime="00:10:26.68" />
                    <SPLIT distance="850" swimtime="00:11:07.59" />
                    <SPLIT distance="900" swimtime="00:11:46.57" />
                    <SPLIT distance="950" swimtime="00:12:26.31" />
                    <SPLIT distance="1000" swimtime="00:13:05.07" />
                    <SPLIT distance="1050" swimtime="00:13:44.90" />
                    <SPLIT distance="1100" swimtime="00:14:23.63" />
                    <SPLIT distance="1150" swimtime="00:15:04.19" />
                    <SPLIT distance="1200" swimtime="00:15:43.36" />
                    <SPLIT distance="1250" swimtime="00:16:23.72" />
                    <SPLIT distance="1300" swimtime="00:17:02.54" />
                    <SPLIT distance="1350" swimtime="00:17:42.12" />
                    <SPLIT distance="1400" swimtime="00:18:20.09" />
                    <SPLIT distance="1450" swimtime="00:18:59.16" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolau" lastname="Neto" birthdate="2011-03-22" gender="M" nation="BRA" license="366906" swrid="5602565" athleteid="3783" externalid="366906">
              <RESULTS>
                <RESULT eventid="1088" points="361" swimtime="00:01:19.81" resultid="3784" heatid="5082" lane="7" entrytime="00:01:21.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="410" swimtime="00:00:28.13" resultid="3785" heatid="5119" lane="2" entrytime="00:00:27.86" entrycourse="LCM" />
                <RESULT eventid="1167" points="447" swimtime="00:01:01.28" resultid="3786" heatid="5222" lane="3" entrytime="00:01:01.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="332" swimtime="00:03:01.08" resultid="3787" heatid="5318" lane="8" entrytime="00:02:58.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.75" />
                    <SPLIT distance="100" swimtime="00:01:25.02" />
                    <SPLIT distance="150" swimtime="00:02:13.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="382" swimtime="00:00:35.75" resultid="3788" heatid="5367" lane="7" entrytime="00:00:40.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Pereira Galle" birthdate="2011-08-02" gender="F" nation="BRA" license="369465" swrid="5627330" athleteid="3928" externalid="369465">
              <RESULTS>
                <RESULT eventid="1080" points="391" swimtime="00:01:27.64" resultid="3929" heatid="5067" lane="1" entrytime="00:01:24.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" points="397" swimtime="00:05:20.07" resultid="3930" heatid="5050" lane="1" entrytime="00:05:12.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:13.47" />
                    <SPLIT distance="150" swimtime="00:01:53.25" />
                    <SPLIT distance="200" swimtime="00:02:33.49" />
                    <SPLIT distance="250" swimtime="00:03:15.04" />
                    <SPLIT distance="300" swimtime="00:03:56.87" />
                    <SPLIT distance="350" swimtime="00:04:38.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="434" swimtime="00:02:28.99" resultid="3931" heatid="5140" lane="6" entrytime="00:02:27.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.53" />
                    <SPLIT distance="100" swimtime="00:01:12.36" />
                    <SPLIT distance="150" swimtime="00:01:51.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="365" swimtime="00:03:12.33" resultid="3932" heatid="5312" lane="3" entrytime="00:03:07.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.59" />
                    <SPLIT distance="100" swimtime="00:01:30.66" />
                    <SPLIT distance="150" swimtime="00:02:21.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="406" swimtime="00:00:39.36" resultid="3933" heatid="5376" lane="7" entrytime="00:00:38.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Clivatti" birthdate="2010-05-24" gender="M" nation="BRA" license="368007" swrid="5600139" athleteid="3814" externalid="368007">
              <RESULTS>
                <RESULT eventid="1072" points="477" swimtime="00:04:41.61" resultid="3815" heatid="5059" lane="5" entrytime="00:04:30.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.50" />
                    <SPLIT distance="100" swimtime="00:01:04.75" />
                    <SPLIT distance="150" swimtime="00:01:40.35" />
                    <SPLIT distance="200" swimtime="00:02:16.56" />
                    <SPLIT distance="250" swimtime="00:02:52.32" />
                    <SPLIT distance="300" swimtime="00:03:28.82" />
                    <SPLIT distance="350" swimtime="00:04:05.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="495" swimtime="00:00:26.42" resultid="3816" heatid="5120" lane="6" entrytime="00:00:26.69" entrycourse="LCM" />
                <RESULT eventid="1120" points="525" swimtime="00:02:06.38" resultid="3817" heatid="5152" lane="5" entrytime="00:02:05.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.73" />
                    <SPLIT distance="100" swimtime="00:01:02.52" />
                    <SPLIT distance="150" swimtime="00:01:35.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="520" swimtime="00:00:58.24" resultid="3818" heatid="5223" lane="5" entrytime="00:00:57.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="318" swimtime="00:00:34.49" resultid="3819" heatid="5283" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Correa Nascimento" birthdate="2009-01-19" gender="M" nation="BRA" license="342235" swrid="5600140" athleteid="3588" externalid="342235">
              <RESULTS>
                <RESULT eventid="1072" points="471" swimtime="00:04:42.66" resultid="3589" heatid="5062" lane="8" entrytime="00:04:36.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.45" />
                    <SPLIT distance="100" swimtime="00:01:05.03" />
                    <SPLIT distance="150" swimtime="00:01:40.26" />
                    <SPLIT distance="200" swimtime="00:02:16.77" />
                    <SPLIT distance="250" swimtime="00:02:53.46" />
                    <SPLIT distance="300" swimtime="00:03:30.86" />
                    <SPLIT distance="350" swimtime="00:04:07.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="472" swimtime="00:02:10.97" resultid="3590" heatid="5155" lane="3" entrytime="00:02:09.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:03.78" />
                    <SPLIT distance="150" swimtime="00:01:37.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="536" swimtime="00:00:57.67" resultid="3591" heatid="5229" lane="6" entrytime="00:00:57.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luis" lastname="Gustavo Souza" birthdate="2011-08-24" gender="M" nation="BRA" license="366901" swrid="5588733" athleteid="3763" externalid="366901">
              <RESULTS>
                <RESULT eventid="1072" points="366" swimtime="00:05:07.60" resultid="3764" heatid="5058" lane="1" entrytime="00:05:07.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.43" />
                    <SPLIT distance="100" swimtime="00:01:15.79" />
                    <SPLIT distance="150" swimtime="00:01:55.59" />
                    <SPLIT distance="200" swimtime="00:02:35.75" />
                    <SPLIT distance="250" swimtime="00:03:14.86" />
                    <SPLIT distance="300" swimtime="00:03:54.40" />
                    <SPLIT distance="350" swimtime="00:04:32.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="331" swimtime="00:01:11.45" resultid="3765" heatid="5170" lane="4" entrytime="00:01:13.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="299" swimtime="00:02:50.36" resultid="3766" heatid="5194" lane="7" entrytime="00:02:48.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                    <SPLIT distance="100" swimtime="00:01:21.94" />
                    <SPLIT distance="150" swimtime="00:02:14.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="256" swimtime="00:01:21.22" resultid="3767" heatid="5256" lane="8" entrytime="00:01:23.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="341" swimtime="00:05:46.82" resultid="3768" heatid="5275" lane="4" entrytime="00:05:56.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.72" />
                    <SPLIT distance="100" swimtime="00:01:17.25" />
                    <SPLIT distance="150" swimtime="00:02:03.78" />
                    <SPLIT distance="200" swimtime="00:02:47.88" />
                    <SPLIT distance="250" swimtime="00:03:39.56" />
                    <SPLIT distance="300" swimtime="00:04:32.29" />
                    <SPLIT distance="350" swimtime="00:05:10.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="294" swimtime="00:00:33.49" resultid="3769" heatid="5331" lane="2" entrytime="00:00:36.02" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Moreira Segadaes" birthdate="2008-05-15" gender="M" nation="BRA" license="331574" swrid="5600220" athleteid="3506" externalid="331574">
              <RESULTS>
                <RESULT eventid="1088" points="590" swimtime="00:01:07.80" resultid="3507" heatid="5085" lane="4" entrytime="00:01:08.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="501" swimtime="00:02:23.53" resultid="3508" heatid="5198" lane="7" entrytime="00:02:22.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.28" />
                    <SPLIT distance="100" swimtime="00:01:08.08" />
                    <SPLIT distance="150" swimtime="00:01:49.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="583" swimtime="00:00:56.08" resultid="3509" heatid="5224" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="535" swimtime="00:02:34.48" resultid="3510" heatid="5320" lane="6" entrytime="00:02:29.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.98" />
                    <SPLIT distance="100" swimtime="00:01:12.77" />
                    <SPLIT distance="150" swimtime="00:01:54.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="592" swimtime="00:00:30.89" resultid="3511" heatid="5371" lane="7" entrytime="00:00:31.14" entrycourse="LCM" />
                <RESULT eventid="2320" points="579" swimtime="00:01:08.21" resultid="5956" heatid="6414" lane="6" entrytime="00:01:07.80">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="Pellanda" birthdate="2010-11-12" gender="M" nation="BRA" license="356352" swrid="5600233" athleteid="3664" externalid="356352">
              <RESULTS>
                <RESULT eventid="1072" points="564" swimtime="00:04:26.30" resultid="3665" heatid="5059" lane="4" entrytime="00:04:21.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.80" />
                    <SPLIT distance="100" swimtime="00:01:02.56" />
                    <SPLIT distance="150" swimtime="00:01:35.51" />
                    <SPLIT distance="200" swimtime="00:02:08.73" />
                    <SPLIT distance="250" swimtime="00:02:42.23" />
                    <SPLIT distance="300" swimtime="00:03:17.03" />
                    <SPLIT distance="350" swimtime="00:03:51.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="486" swimtime="00:00:26.59" resultid="3666" heatid="5119" lane="6" entrytime="00:00:27.73" entrycourse="LCM" />
                <RESULT eventid="1120" points="539" swimtime="00:02:05.28" resultid="3667" heatid="5152" lane="4" entrytime="00:02:03.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                    <SPLIT distance="100" swimtime="00:01:02.20" />
                    <SPLIT distance="150" swimtime="00:01:33.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="543" swimtime="00:00:57.42" resultid="3668" heatid="5223" lane="6" entrytime="00:00:58.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="582" swimtime="00:09:01.45" resultid="3669" heatid="5300" lane="4" entrytime="00:08:57.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.34" />
                    <SPLIT distance="100" swimtime="00:01:03.30" />
                    <SPLIT distance="150" swimtime="00:01:37.81" />
                    <SPLIT distance="200" swimtime="00:02:12.35" />
                    <SPLIT distance="250" swimtime="00:02:46.96" />
                    <SPLIT distance="300" swimtime="00:03:21.96" />
                    <SPLIT distance="350" swimtime="00:03:56.67" />
                    <SPLIT distance="400" swimtime="00:04:31.49" />
                    <SPLIT distance="450" swimtime="00:05:05.31" />
                    <SPLIT distance="500" swimtime="00:05:39.96" />
                    <SPLIT distance="550" swimtime="00:06:14.59" />
                    <SPLIT distance="600" swimtime="00:06:49.33" />
                    <SPLIT distance="650" swimtime="00:07:23.60" />
                    <SPLIT distance="700" swimtime="00:07:58.14" />
                    <SPLIT distance="750" swimtime="00:08:31.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="312" swimtime="00:00:32.82" resultid="3670" heatid="5327" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Coelho" birthdate="2011-11-11" gender="M" nation="BRA" license="366889" swrid="5602527" athleteid="3727" externalid="366889">
              <RESULTS>
                <RESULT eventid="1072" points="423" swimtime="00:04:53.05" resultid="3728" heatid="5058" lane="3" entrytime="00:04:57.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                    <SPLIT distance="100" swimtime="00:01:09.49" />
                    <SPLIT distance="150" swimtime="00:01:46.64" />
                    <SPLIT distance="200" swimtime="00:02:24.12" />
                    <SPLIT distance="250" swimtime="00:03:01.48" />
                    <SPLIT distance="300" swimtime="00:03:38.97" />
                    <SPLIT distance="350" swimtime="00:04:16.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="315" swimtime="00:01:12.66" resultid="3729" heatid="5171" lane="7" entrytime="00:01:12.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="388" swimtime="00:02:19.79" resultid="3730" heatid="5151" lane="7" entrytime="00:02:22.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                    <SPLIT distance="150" swimtime="00:01:43.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="356" swimtime="00:00:31.42" resultid="3731" heatid="5332" lane="7" entrytime="00:00:33.16" entrycourse="LCM" />
                <RESULT eventid="1293" points="304" swimtime="00:02:44.03" resultid="3732" heatid="5358" lane="3" entrytime="00:02:45.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                    <SPLIT distance="100" swimtime="00:01:17.74" />
                    <SPLIT distance="150" swimtime="00:02:01.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Emili Da Silva Gomes Xavier" birthdate="2010-09-08" gender="F" nation="BRA" license="372519" swrid="5717260" athleteid="3969" externalid="372519">
              <RESULTS>
                <RESULT eventid="1064" points="451" swimtime="00:05:06.82" resultid="3970" heatid="5049" lane="3" entrytime="00:05:29.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.23" />
                    <SPLIT distance="100" swimtime="00:01:12.11" />
                    <SPLIT distance="150" swimtime="00:01:52.40" />
                    <SPLIT distance="200" swimtime="00:02:32.44" />
                    <SPLIT distance="250" swimtime="00:03:12.42" />
                    <SPLIT distance="300" swimtime="00:03:52.25" />
                    <SPLIT distance="350" swimtime="00:04:30.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="521" swimtime="00:00:29.33" resultid="3971" heatid="5099" lane="6" entrytime="00:00:31.30" entrycourse="LCM" />
                <RESULT eventid="1112" points="496" swimtime="00:02:22.48" resultid="3972" heatid="5139" lane="4" entrytime="00:02:30.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.07" />
                    <SPLIT distance="100" swimtime="00:01:09.60" />
                    <SPLIT distance="150" swimtime="00:01:46.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="391" swimtime="00:02:52.43" resultid="3973" heatid="5187" lane="5" entrytime="00:02:56.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                    <SPLIT distance="100" swimtime="00:01:26.55" />
                    <SPLIT distance="150" swimtime="00:02:17.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="506" swimtime="00:01:04.87" resultid="3974" heatid="5205" lane="1" entrytime="00:01:06.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1275" points="339" swimtime="00:02:56.51" resultid="3975" heatid="5341" lane="7" entrytime="00:02:53.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                    <SPLIT distance="100" swimtime="00:01:27.03" />
                    <SPLIT distance="150" swimtime="00:02:12.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2375" swimtime="00:00:00.00" resultid="6455" entrytime="00:00:29.33" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Kirchgassner" birthdate="2007-02-10" gender="M" nation="BRA" license="313535" swrid="5600230" athleteid="3557" externalid="313535">
              <RESULTS>
                <RESULT eventid="1088" points="595" swimtime="00:01:07.59" resultid="3558" heatid="5087" lane="4" entrytime="00:01:05.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="534" swimtime="00:00:25.76" resultid="3559" heatid="5127" lane="6" />
                <RESULT eventid="1151" points="577" swimtime="00:02:16.89" resultid="3560" heatid="5200" lane="4" entrytime="00:02:13.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                    <SPLIT distance="100" swimtime="00:01:05.60" />
                    <SPLIT distance="150" swimtime="00:01:45.29" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.1 - Mais de uma pernada de borboleta antes da primeira pernada de peito após o início ou a virada.  (Horário: 10:06), Após a saida." eventid="1251" status="DSQ" swimtime="00:02:24.40" resultid="3561" heatid="5320" lane="4" entrytime="00:02:21.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                    <SPLIT distance="100" swimtime="00:01:09.46" />
                    <SPLIT distance="150" swimtime="00:01:47.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="556" swimtime="00:00:31.54" resultid="3562" heatid="5371" lane="1" entrytime="00:00:31.14" entrycourse="LCM" />
                <RESULT eventid="2320" points="613" swimtime="00:01:06.93" resultid="5955" heatid="6414" lane="3" entrytime="00:01:07.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Germer Munhoz" birthdate="2010-04-23" gender="F" nation="BRA" license="356632" swrid="5588722" athleteid="3696" externalid="356632">
              <RESULTS>
                <RESULT eventid="1064" points="490" swimtime="00:04:58.45" resultid="3697" heatid="5051" lane="5" entrytime="00:04:54.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:10.48" />
                    <SPLIT distance="150" swimtime="00:01:48.58" />
                    <SPLIT distance="200" swimtime="00:02:26.63" />
                    <SPLIT distance="250" swimtime="00:03:05.32" />
                    <SPLIT distance="300" swimtime="00:03:43.52" />
                    <SPLIT distance="350" swimtime="00:04:22.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" points="458" swimtime="00:01:11.96" resultid="3698" heatid="5160" lane="5" entrytime="00:01:12.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="454" swimtime="00:02:44.09" resultid="3699" heatid="5188" lane="2" entrytime="00:02:44.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                    <SPLIT distance="100" swimtime="00:01:17.76" />
                    <SPLIT distance="150" swimtime="00:02:07.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="473" swimtime="00:10:22.02" resultid="3700" heatid="5271" lane="4" entrytime="00:10:13.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                    <SPLIT distance="100" swimtime="00:01:11.18" />
                    <SPLIT distance="150" swimtime="00:01:50.21" />
                    <SPLIT distance="200" swimtime="00:02:29.37" />
                    <SPLIT distance="250" swimtime="00:03:08.68" />
                    <SPLIT distance="300" swimtime="00:03:47.27" />
                    <SPLIT distance="350" swimtime="00:04:26.92" />
                    <SPLIT distance="400" swimtime="00:05:06.46" />
                    <SPLIT distance="450" swimtime="00:05:46.18" />
                    <SPLIT distance="500" swimtime="00:06:25.57" />
                    <SPLIT distance="550" swimtime="00:07:05.60" />
                    <SPLIT distance="600" swimtime="00:07:45.61" />
                    <SPLIT distance="650" swimtime="00:08:24.98" />
                    <SPLIT distance="700" swimtime="00:09:04.37" />
                    <SPLIT distance="750" swimtime="00:09:44.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="429" swimtime="00:00:32.38" resultid="3701" heatid="5321" lane="2" />
                <RESULT eventid="1295" points="394" swimtime="00:02:46.15" resultid="3702" heatid="5362" lane="2" entrytime="00:02:49.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:18.00" />
                    <SPLIT distance="150" swimtime="00:02:03.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2328" points="433" swimtime="00:01:13.32" resultid="6000" heatid="6418" lane="6" entrytime="00:01:11.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Fontana" birthdate="2011-12-29" gender="M" nation="BRA" license="366897" swrid="5602539" athleteid="3750" externalid="366897">
              <RESULTS>
                <RESULT eventid="1088" points="217" swimtime="00:01:34.65" resultid="3751" heatid="5079" lane="6" entrytime="00:01:43.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="209" swimtime="00:03:12.02" resultid="3752" heatid="5193" lane="7" entrytime="00:03:16.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:33.30" />
                    <SPLIT distance="150" swimtime="00:02:27.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="197" swimtime="00:01:28.66" resultid="3753" heatid="5255" lane="4" entrytime="00:01:28.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="180" swimtime="00:03:42.16" resultid="3754" heatid="5316" lane="7" entrytime="00:03:40.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.16" />
                    <SPLIT distance="100" swimtime="00:01:44.40" />
                    <SPLIT distance="150" swimtime="00:02:43.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="211" swimtime="00:00:43.56" resultid="3755" heatid="5366" lane="7" entrytime="00:00:48.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1237" points="648" swimtime="00:03:37.48" resultid="3995" heatid="5308" lane="4" entrytime="00:03:42.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.67" />
                    <SPLIT distance="100" swimtime="00:00:53.65" />
                    <SPLIT distance="150" swimtime="00:01:20.06" />
                    <SPLIT distance="200" swimtime="00:01:48.78" />
                    <SPLIT distance="250" swimtime="00:02:14.66" />
                    <SPLIT distance="300" swimtime="00:02:42.96" />
                    <SPLIT distance="350" swimtime="00:03:08.35" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3485" number="1" />
                    <RELAYPOSITION athleteid="3491" number="2" />
                    <RELAYPOSITION athleteid="3502" number="3" />
                    <RELAYPOSITION athleteid="3934" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1338" points="557" swimtime="00:04:11.22" resultid="4004" heatid="5388" lane="4" entrytime="00:04:06.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.09" />
                    <SPLIT distance="100" swimtime="00:01:06.84" />
                    <SPLIT distance="150" swimtime="00:01:39.39" />
                    <SPLIT distance="200" swimtime="00:02:15.26" />
                    <SPLIT distance="250" swimtime="00:02:43.71" />
                    <SPLIT distance="300" swimtime="00:03:16.83" />
                    <SPLIT distance="350" swimtime="00:03:42.16" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3568" number="1" />
                    <RELAYPOSITION athleteid="3506" number="2" />
                    <RELAYPOSITION athleteid="3491" number="3" />
                    <RELAYPOSITION athleteid="3934" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="19" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1239" points="654" swimtime="00:03:36.81" resultid="3996" heatid="5309" lane="3" entrytime="00:03:24.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.46" />
                    <SPLIT distance="100" swimtime="00:00:52.43" />
                    <SPLIT distance="150" swimtime="00:01:17.97" />
                    <SPLIT distance="200" swimtime="00:01:46.12" />
                    <SPLIT distance="250" swimtime="00:02:12.59" />
                    <SPLIT distance="300" swimtime="00:02:41.83" />
                    <SPLIT distance="350" swimtime="00:03:07.88" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3478" number="1" />
                    <RELAYPOSITION athleteid="3981" number="2" />
                    <RELAYPOSITION athleteid="3714" number="3" />
                    <RELAYPOSITION athleteid="3557" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1340" points="644" swimtime="00:03:59.40" resultid="4001" heatid="5389" lane="3" entrytime="00:03:47.98">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                    <SPLIT distance="100" swimtime="00:01:00.58" />
                    <SPLIT distance="150" swimtime="00:01:32.44" />
                    <SPLIT distance="200" swimtime="00:02:08.07" />
                    <SPLIT distance="250" swimtime="00:02:36.75" />
                    <SPLIT distance="300" swimtime="00:03:07.61" />
                    <SPLIT distance="350" swimtime="00:03:32.22" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3478" number="1" />
                    <RELAYPOSITION athleteid="3557" number="2" />
                    <RELAYPOSITION athleteid="3981" number="3" />
                    <RELAYPOSITION athleteid="3551" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1235" points="608" swimtime="00:03:42.15" resultid="3997" heatid="5307" lane="4" entrytime="00:03:49.59">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.57" />
                    <SPLIT distance="100" swimtime="00:00:55.72" />
                    <SPLIT distance="150" swimtime="00:01:22.37" />
                    <SPLIT distance="200" swimtime="00:01:51.60" />
                    <SPLIT distance="250" swimtime="00:02:18.95" />
                    <SPLIT distance="300" swimtime="00:02:48.36" />
                    <SPLIT distance="350" swimtime="00:03:14.08" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3976" number="1" />
                    <RELAYPOSITION athleteid="3945" number="2" />
                    <RELAYPOSITION athleteid="3539" number="3" />
                    <RELAYPOSITION athleteid="3497" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1336" points="572" swimtime="00:04:09.08" resultid="4005" heatid="5387" lane="4" entrytime="00:04:15.46">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.70" />
                    <SPLIT distance="100" swimtime="00:01:01.07" />
                    <SPLIT distance="150" swimtime="00:01:35.42" />
                    <SPLIT distance="200" swimtime="00:02:13.95" />
                    <SPLIT distance="250" swimtime="00:02:42.58" />
                    <SPLIT distance="300" swimtime="00:03:14.68" />
                    <SPLIT distance="350" swimtime="00:03:40.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3976" number="1" />
                    <RELAYPOSITION athleteid="3602" number="2" />
                    <RELAYPOSITION athleteid="3945" number="3" />
                    <RELAYPOSITION athleteid="3497" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1233" points="528" swimtime="00:03:52.77" resultid="3998" heatid="5306" lane="4" entrytime="00:03:58.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                    <SPLIT distance="100" swimtime="00:00:58.24" />
                    <SPLIT distance="150" swimtime="00:01:25.90" />
                    <SPLIT distance="200" swimtime="00:01:56.41" />
                    <SPLIT distance="250" swimtime="00:02:24.30" />
                    <SPLIT distance="300" swimtime="00:02:55.00" />
                    <SPLIT distance="350" swimtime="00:03:22.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3671" number="1" />
                    <RELAYPOSITION athleteid="3896" number="2" />
                    <RELAYPOSITION athleteid="3664" number="3" />
                    <RELAYPOSITION athleteid="3814" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1334" points="411" swimtime="00:04:37.95" resultid="4003" heatid="5386" lane="5" entrytime="00:04:38.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.89" />
                    <SPLIT distance="150" swimtime="00:01:46.81" />
                    <SPLIT distance="200" swimtime="00:02:28.26" />
                    <SPLIT distance="250" swimtime="00:03:00.73" />
                    <SPLIT distance="300" swimtime="00:03:39.65" />
                    <SPLIT distance="350" swimtime="00:04:07.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3671" number="1" />
                    <RELAYPOSITION athleteid="3690" number="2" />
                    <RELAYPOSITION athleteid="3627" number="3" />
                    <RELAYPOSITION athleteid="3896" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1231" points="440" swimtime="00:04:07.43" resultid="3999" heatid="5305" lane="4" entrytime="00:04:04.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.18" />
                    <SPLIT distance="100" swimtime="00:00:58.96" />
                    <SPLIT distance="150" swimtime="00:01:28.64" />
                    <SPLIT distance="200" swimtime="00:02:00.99" />
                    <SPLIT distance="250" swimtime="00:02:31.59" />
                    <SPLIT distance="300" swimtime="00:03:05.29" />
                    <SPLIT distance="350" swimtime="00:03:34.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3825" number="1" />
                    <RELAYPOSITION athleteid="3783" number="2" />
                    <RELAYPOSITION athleteid="3727" number="3" />
                    <RELAYPOSITION athleteid="3733" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1332" points="398" swimtime="00:04:40.95" resultid="4002" heatid="5385" lane="5" entrytime="00:04:54.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.62" />
                    <SPLIT distance="100" swimtime="00:01:09.26" />
                    <SPLIT distance="150" swimtime="00:01:46.43" />
                    <SPLIT distance="200" swimtime="00:02:27.80" />
                    <SPLIT distance="250" swimtime="00:03:01.65" />
                    <SPLIT distance="300" swimtime="00:03:38.54" />
                    <SPLIT distance="350" swimtime="00:04:08.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3825" number="1" />
                    <RELAYPOSITION athleteid="3733" number="2" />
                    <RELAYPOSITION athleteid="3727" number="3" />
                    <RELAYPOSITION athleteid="3783" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="20" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1342" status="WDR" swimtime="00:00:00.00" resultid="4000" heatid="5390" lane="8" entrytime="00:03:57.97" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="19" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1239" points="658" swimtime="00:03:36.35" resultid="4016" heatid="5309" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.81" />
                    <SPLIT distance="100" swimtime="00:00:57.44" />
                    <SPLIT distance="150" swimtime="00:01:24.53" />
                    <SPLIT distance="200" swimtime="00:01:53.82" />
                    <SPLIT distance="250" swimtime="00:02:18.45" />
                    <SPLIT distance="300" swimtime="00:02:45.84" />
                    <SPLIT distance="350" swimtime="00:03:10.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3516" number="1" />
                    <RELAYPOSITION athleteid="3964" number="2" />
                    <RELAYPOSITION athleteid="3958" number="3" />
                    <RELAYPOSITION athleteid="3551" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1340" status="WDR" swimtime="00:00:00.00" resultid="4019" heatid="5389" lane="2" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1233" points="453" swimtime="00:04:05.04" resultid="4017" heatid="5306" lane="3" entrytime="00:04:04.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.82" />
                    <SPLIT distance="150" swimtime="00:01:29.71" />
                    <SPLIT distance="200" swimtime="00:02:02.75" />
                    <SPLIT distance="250" swimtime="00:02:32.50" />
                    <SPLIT distance="300" swimtime="00:03:03.93" />
                    <SPLIT distance="350" swimtime="00:03:32.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3690" number="1" />
                    <RELAYPOSITION athleteid="3703" number="2" />
                    <RELAYPOSITION athleteid="3677" number="3" />
                    <RELAYPOSITION athleteid="3627" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1334" points="377" swimtime="00:04:46.20" resultid="4021" heatid="5386" lane="2" entrytime="00:04:48.18">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.36" />
                    <SPLIT distance="100" swimtime="00:01:12.34" />
                    <SPLIT distance="150" swimtime="00:01:49.93" />
                    <SPLIT distance="200" swimtime="00:02:33.05" />
                    <SPLIT distance="250" swimtime="00:03:08.66" />
                    <SPLIT distance="300" swimtime="00:03:48.09" />
                    <SPLIT distance="350" swimtime="00:04:15.95" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3633" number="1" />
                    <RELAYPOSITION athleteid="3677" number="2" />
                    <RELAYPOSITION athleteid="3703" number="3" />
                    <RELAYPOSITION athleteid="3814" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1231" points="353" swimtime="00:04:26.24" resultid="4018" heatid="5305" lane="5" entrytime="00:04:17.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="100" swimtime="00:01:04.69" />
                    <SPLIT distance="150" swimtime="00:01:36.71" />
                    <SPLIT distance="200" swimtime="00:02:11.60" />
                    <SPLIT distance="250" swimtime="00:02:44.07" />
                    <SPLIT distance="300" swimtime="00:03:19.63" />
                    <SPLIT distance="350" swimtime="00:03:51.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3720" number="1" />
                    <RELAYPOSITION athleteid="3801" number="2" />
                    <RELAYPOSITION athleteid="3763" number="3" />
                    <RELAYPOSITION athleteid="3873" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1332" points="318" swimtime="00:05:02.92" resultid="4020" heatid="5385" lane="6" entrytime="00:05:06.31">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                    <SPLIT distance="100" swimtime="00:01:17.60" />
                    <SPLIT distance="150" swimtime="00:01:58.87" />
                    <SPLIT distance="200" swimtime="00:02:44.55" />
                    <SPLIT distance="250" swimtime="00:03:18.24" />
                    <SPLIT distance="300" swimtime="00:03:57.00" />
                    <SPLIT distance="350" swimtime="00:04:28.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3789" number="1" />
                    <RELAYPOSITION athleteid="3861" number="2" />
                    <RELAYPOSITION athleteid="3763" number="3" />
                    <RELAYPOSITION athleteid="3720" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1223" points="538" swimtime="00:04:15.58" resultid="3987" heatid="5303" lane="2" entrytime="00:04:12.44">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.53" />
                    <SPLIT distance="100" swimtime="00:01:02.32" />
                    <SPLIT distance="150" swimtime="00:01:33.11" />
                    <SPLIT distance="200" swimtime="00:02:06.58" />
                    <SPLIT distance="250" swimtime="00:02:37.84" />
                    <SPLIT distance="300" swimtime="00:03:10.78" />
                    <SPLIT distance="350" swimtime="00:03:42.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3473" number="1" />
                    <RELAYPOSITION athleteid="3607" number="2" />
                    <RELAYPOSITION athleteid="3461" number="3" />
                    <RELAYPOSITION athleteid="3592" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1324" points="445" swimtime="00:05:01.58" resultid="3992" heatid="5383" lane="3" entrytime="00:04:52.51">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.40" />
                    <SPLIT distance="100" swimtime="00:01:17.54" />
                    <SPLIT distance="150" swimtime="00:01:55.63" />
                    <SPLIT distance="200" swimtime="00:02:38.49" />
                    <SPLIT distance="250" swimtime="00:03:13.41" />
                    <SPLIT distance="300" swimtime="00:03:55.77" />
                    <SPLIT distance="350" swimtime="00:04:27.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3473" number="1" />
                    <RELAYPOSITION athleteid="3592" number="2" />
                    <RELAYPOSITION athleteid="3534" number="3" />
                    <RELAYPOSITION athleteid="3597" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1221" points="496" swimtime="00:04:22.65" resultid="3988" heatid="5302" lane="4" entrytime="00:04:19.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:04.76" />
                    <SPLIT distance="150" swimtime="00:01:35.63" />
                    <SPLIT distance="200" swimtime="00:02:10.08" />
                    <SPLIT distance="250" swimtime="00:02:41.24" />
                    <SPLIT distance="300" swimtime="00:03:16.31" />
                    <SPLIT distance="350" swimtime="00:03:47.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3696" number="1" />
                    <RELAYPOSITION athleteid="3969" number="2" />
                    <RELAYPOSITION athleteid="3651" number="3" />
                    <RELAYPOSITION athleteid="3645" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1322" points="457" swimtime="00:04:58.95" resultid="3993" heatid="5382" lane="4" entrytime="00:04:57.86">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                    <SPLIT distance="100" swimtime="00:01:15.98" />
                    <SPLIT distance="150" swimtime="00:01:56.56" />
                    <SPLIT distance="200" swimtime="00:02:40.91" />
                    <SPLIT distance="250" swimtime="00:03:15.63" />
                    <SPLIT distance="300" swimtime="00:03:53.84" />
                    <SPLIT distance="350" swimtime="00:04:24.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3651" number="1" />
                    <RELAYPOSITION athleteid="3528" number="2" />
                    <RELAYPOSITION athleteid="3696" number="3" />
                    <RELAYPOSITION athleteid="3645" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1219" points="508" swimtime="00:04:20.61" resultid="3989" heatid="5301" lane="4" entrytime="00:04:29.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                    <SPLIT distance="100" swimtime="00:01:05.12" />
                    <SPLIT distance="150" swimtime="00:01:37.14" />
                    <SPLIT distance="200" swimtime="00:02:11.58" />
                    <SPLIT distance="250" swimtime="00:02:43.26" />
                    <SPLIT distance="300" swimtime="00:03:17.92" />
                    <SPLIT distance="350" swimtime="00:03:47.93" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3777" number="1" />
                    <RELAYPOSITION athleteid="3795" number="2" />
                    <RELAYPOSITION athleteid="3743" number="3" />
                    <RELAYPOSITION athleteid="3849" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1320" points="488" swimtime="00:04:52.46" resultid="3994" heatid="5381" lane="4" entrytime="00:04:59.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.74" />
                    <SPLIT distance="100" swimtime="00:01:16.40" />
                    <SPLIT distance="150" swimtime="00:01:55.75" />
                    <SPLIT distance="200" swimtime="00:02:41.55" />
                    <SPLIT distance="250" swimtime="00:03:12.41" />
                    <SPLIT distance="300" swimtime="00:03:48.78" />
                    <SPLIT distance="350" swimtime="00:04:19.02" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3795" number="1" />
                    <RELAYPOSITION athleteid="3743" number="2" />
                    <RELAYPOSITION athleteid="3849" number="3" />
                    <RELAYPOSITION athleteid="3777" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1225" points="541" swimtime="00:04:15.19" resultid="3990" heatid="5304" lane="5" entrytime="00:04:10.66">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                    <SPLIT distance="100" swimtime="00:01:02.87" />
                    <SPLIT distance="150" swimtime="00:01:32.92" />
                    <SPLIT distance="200" swimtime="00:02:06.90" />
                    <SPLIT distance="250" swimtime="00:02:37.68" />
                    <SPLIT distance="300" swimtime="00:03:12.36" />
                    <SPLIT distance="350" swimtime="00:03:42.19" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3457" number="1" />
                    <RELAYPOSITION athleteid="3845" number="2" />
                    <RELAYPOSITION athleteid="3940" number="3" />
                    <RELAYPOSITION athleteid="3466" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1326" status="WDR" swimtime="00:00:00.00" resultid="3991" heatid="5384" lane="5" entrytime="00:04:42.72" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1221" points="442" swimtime="00:04:32.90" resultid="4012" heatid="5302" lane="3" entrytime="00:04:34.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                    <SPLIT distance="100" swimtime="00:01:06.66" />
                    <SPLIT distance="150" swimtime="00:01:38.91" />
                    <SPLIT distance="200" swimtime="00:02:13.49" />
                    <SPLIT distance="250" swimtime="00:02:46.10" />
                    <SPLIT distance="300" swimtime="00:03:21.81" />
                    <SPLIT distance="350" swimtime="00:03:55.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3658" number="1" />
                    <RELAYPOSITION athleteid="3528" number="2" />
                    <RELAYPOSITION athleteid="3684" number="3" />
                    <RELAYPOSITION athleteid="3639" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1322" points="385" swimtime="00:05:16.46" resultid="4014" heatid="5382" lane="3" entrytime="00:05:16.01">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                    <SPLIT distance="100" swimtime="00:01:17.20" />
                    <SPLIT distance="150" swimtime="00:01:59.03" />
                    <SPLIT distance="200" swimtime="00:02:44.47" />
                    <SPLIT distance="250" swimtime="00:03:24.92" />
                    <SPLIT distance="300" swimtime="00:04:11.12" />
                    <SPLIT distance="350" swimtime="00:04:42.25" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3639" number="1" />
                    <RELAYPOSITION athleteid="3969" number="2" />
                    <RELAYPOSITION athleteid="3684" number="3" />
                    <RELAYPOSITION athleteid="3658" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1219" points="429" swimtime="00:04:35.60" resultid="4013" heatid="5301" lane="5" entrytime="00:04:37.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                    <SPLIT distance="100" swimtime="00:01:09.32" />
                    <SPLIT distance="150" swimtime="00:01:41.65" />
                    <SPLIT distance="200" swimtime="00:02:17.44" />
                    <SPLIT distance="250" swimtime="00:02:50.93" />
                    <SPLIT distance="300" swimtime="00:03:28.39" />
                    <SPLIT distance="350" swimtime="00:04:00.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3838" number="1" />
                    <RELAYPOSITION athleteid="3770" number="2" />
                    <RELAYPOSITION athleteid="3921" number="3" />
                    <RELAYPOSITION athleteid="3928" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1320" points="372" swimtime="00:05:20.12" resultid="4015" heatid="5381" lane="5" entrytime="00:05:27.14">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.14" />
                    <SPLIT distance="100" swimtime="00:01:18.17" />
                    <SPLIT distance="150" swimtime="00:02:00.86" />
                    <SPLIT distance="200" swimtime="00:02:46.08" />
                    <SPLIT distance="250" swimtime="00:03:23.85" />
                    <SPLIT distance="300" swimtime="00:04:10.07" />
                    <SPLIT distance="350" swimtime="00:04:43.28" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3921" number="1" />
                    <RELAYPOSITION athleteid="3770" number="2" />
                    <RELAYPOSITION athleteid="3928" number="3" />
                    <RELAYPOSITION athleteid="3838" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1287" points="567" swimtime="00:04:22.88" resultid="4006" heatid="5354" lane="4" entrytime="00:04:22.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.07" />
                    <SPLIT distance="100" swimtime="00:01:10.52" />
                    <SPLIT distance="150" swimtime="00:01:48.45" />
                    <SPLIT distance="200" swimtime="00:02:30.07" />
                    <SPLIT distance="250" swimtime="00:02:56.80" />
                    <SPLIT distance="300" swimtime="00:03:29.12" />
                    <SPLIT distance="350" swimtime="00:03:54.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3940" number="1" />
                    <RELAYPOSITION athleteid="3457" number="2" />
                    <RELAYPOSITION athleteid="3574" number="3" />
                    <RELAYPOSITION athleteid="3934" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="19" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1289" points="561" swimtime="00:04:23.70" resultid="4007" heatid="5355" lane="3" entrytime="00:04:11.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.34" />
                    <SPLIT distance="100" swimtime="00:01:03.16" />
                    <SPLIT distance="150" swimtime="00:01:40.31" />
                    <SPLIT distance="200" swimtime="00:02:21.02" />
                    <SPLIT distance="250" swimtime="00:02:48.89" />
                    <SPLIT distance="300" swimtime="00:03:21.00" />
                    <SPLIT distance="350" swimtime="00:03:51.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3478" number="1" />
                    <RELAYPOSITION athleteid="3951" number="2" />
                    <RELAYPOSITION athleteid="3981" number="3" />
                    <RELAYPOSITION athleteid="3545" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="20" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1291" points="519" swimtime="00:04:30.61" resultid="4008" heatid="5356" lane="5" entrytime="00:04:10.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.35" />
                    <SPLIT distance="100" swimtime="00:01:01.17" />
                    <SPLIT distance="150" swimtime="00:01:40.92" />
                    <SPLIT distance="200" swimtime="00:02:25.28" />
                    <SPLIT distance="250" swimtime="00:02:58.87" />
                    <SPLIT distance="300" swimtime="00:03:35.15" />
                    <SPLIT distance="350" swimtime="00:04:01.57" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3807" number="1" />
                    <RELAYPOSITION athleteid="3902" number="2" />
                    <RELAYPOSITION athleteid="3914" number="3" />
                    <RELAYPOSITION athleteid="3890" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1285" points="540" swimtime="00:04:27.15" resultid="4009" heatid="5353" lane="4" entrytime="00:04:29.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                    <SPLIT distance="100" swimtime="00:01:03.13" />
                    <SPLIT distance="150" swimtime="00:01:41.97" />
                    <SPLIT distance="200" swimtime="00:02:23.47" />
                    <SPLIT distance="250" swimtime="00:02:51.96" />
                    <SPLIT distance="300" swimtime="00:03:24.43" />
                    <SPLIT distance="350" swimtime="00:03:54.07" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3976" number="1" />
                    <RELAYPOSITION athleteid="3592" number="2" />
                    <RELAYPOSITION athleteid="3945" number="3" />
                    <RELAYPOSITION athleteid="3473" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1283" points="444" swimtime="00:04:45.11" resultid="4010" heatid="5352" lane="5" entrytime="00:04:42.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="100" swimtime="00:01:07.98" />
                    <SPLIT distance="150" swimtime="00:01:49.30" />
                    <SPLIT distance="200" swimtime="00:02:33.14" />
                    <SPLIT distance="250" swimtime="00:03:06.29" />
                    <SPLIT distance="300" swimtime="00:03:46.02" />
                    <SPLIT distance="350" swimtime="00:04:13.98" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3896" number="1" />
                    <RELAYPOSITION athleteid="3528" number="2" />
                    <RELAYPOSITION athleteid="3696" number="3" />
                    <RELAYPOSITION athleteid="3814" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1281" points="478" swimtime="00:04:38.24" resultid="4011" heatid="5351" lane="4" entrytime="00:04:53.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                    <SPLIT distance="100" swimtime="00:01:09.55" />
                    <SPLIT distance="150" swimtime="00:01:47.71" />
                    <SPLIT distance="200" swimtime="00:02:28.24" />
                    <SPLIT distance="250" swimtime="00:02:59.42" />
                    <SPLIT distance="300" swimtime="00:03:34.43" />
                    <SPLIT distance="350" swimtime="00:04:05.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3825" number="1" />
                    <RELAYPOSITION athleteid="3733" number="2" />
                    <RELAYPOSITION athleteid="3849" number="3" />
                    <RELAYPOSITION athleteid="3777" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1287" points="545" swimtime="00:04:26.31" resultid="4022" heatid="5354" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                    <SPLIT distance="100" swimtime="00:01:03.04" />
                    <SPLIT distance="150" swimtime="00:01:41.91" />
                    <SPLIT distance="200" swimtime="00:02:23.90" />
                    <SPLIT distance="250" swimtime="00:02:55.74" />
                    <SPLIT distance="300" swimtime="00:03:31.01" />
                    <SPLIT distance="350" swimtime="00:03:56.97" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3485" number="1" />
                    <RELAYPOSITION athleteid="3845" number="2" />
                    <RELAYPOSITION athleteid="3466" number="3" />
                    <RELAYPOSITION athleteid="3502" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1285" points="480" swimtime="00:04:37.81" resultid="4023" heatid="5353" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                    <SPLIT distance="100" swimtime="00:01:05.47" />
                    <SPLIT distance="150" swimtime="00:01:43.30" />
                    <SPLIT distance="200" swimtime="00:02:27.13" />
                    <SPLIT distance="250" swimtime="00:02:56.58" />
                    <SPLIT distance="300" swimtime="00:03:31.73" />
                    <SPLIT distance="350" swimtime="00:04:03.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3616" number="1" />
                    <RELAYPOSITION athleteid="3534" number="2" />
                    <RELAYPOSITION athleteid="3539" number="3" />
                    <RELAYPOSITION athleteid="3597" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1283" points="403" swimtime="00:04:54.49" resultid="4024" heatid="5352" lane="6" entrytime="00:04:53.37">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:08.16" />
                    <SPLIT distance="150" swimtime="00:01:49.65" />
                    <SPLIT distance="200" swimtime="00:02:36.11" />
                    <SPLIT distance="250" swimtime="00:03:09.40" />
                    <SPLIT distance="300" swimtime="00:03:49.31" />
                    <SPLIT distance="350" swimtime="00:04:20.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3671" number="1" />
                    <RELAYPOSITION athleteid="3969" number="2" />
                    <RELAYPOSITION athleteid="3690" number="3" />
                    <RELAYPOSITION athleteid="3645" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="CURITIBANO &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1281" points="408" swimtime="00:04:53.24" resultid="4025" heatid="5351" lane="6" entrytime="00:05:07.33">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.59" />
                    <SPLIT distance="150" swimtime="00:01:55.51" />
                    <SPLIT distance="200" swimtime="00:02:39.95" />
                    <SPLIT distance="250" swimtime="00:03:13.98" />
                    <SPLIT distance="300" swimtime="00:03:51.40" />
                    <SPLIT distance="350" swimtime="00:04:20.49" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3795" number="1" />
                    <RELAYPOSITION athleteid="3743" number="2" />
                    <RELAYPOSITION athleteid="3727" number="3" />
                    <RELAYPOSITION athleteid="3783" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="16830" nation="BRA" region="PR" clubid="2863" swrid="94883" name="Arenna Carvalho Ltda" shortname="Arenna Carvalho">
          <ATHLETES>
            <ATHLETE firstname="Nicolle" lastname="Akemi Wajima" birthdate="2008-02-01" gender="F" nation="BRA" license="399346" swrid="5658056" athleteid="2864" externalid="399346">
              <RESULTS>
                <RESULT eventid="1064" points="414" swimtime="00:05:15.68" resultid="2865" heatid="5053" lane="6" entrytime="00:05:11.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.67" />
                    <SPLIT distance="100" swimtime="00:01:11.29" />
                    <SPLIT distance="150" swimtime="00:01:51.06" />
                    <SPLIT distance="200" swimtime="00:02:31.87" />
                    <SPLIT distance="250" swimtime="00:03:12.85" />
                    <SPLIT distance="300" swimtime="00:03:55.01" />
                    <SPLIT distance="350" swimtime="00:04:36.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="440" swimtime="00:02:28.34" resultid="2866" heatid="5142" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.55" />
                    <SPLIT distance="100" swimtime="00:01:10.63" />
                    <SPLIT distance="150" swimtime="00:01:49.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="404" swimtime="00:10:55.57" resultid="2867" heatid="5272" lane="6" entrytime="00:10:44.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:01:12.52" />
                    <SPLIT distance="150" swimtime="00:01:52.68" />
                    <SPLIT distance="200" swimtime="00:02:34.18" />
                    <SPLIT distance="250" swimtime="00:03:15.65" />
                    <SPLIT distance="300" swimtime="00:03:57.32" />
                    <SPLIT distance="350" swimtime="00:04:38.61" />
                    <SPLIT distance="400" swimtime="00:05:20.61" />
                    <SPLIT distance="450" swimtime="00:06:02.95" />
                    <SPLIT distance="500" swimtime="00:06:44.82" />
                    <SPLIT distance="550" swimtime="00:07:26.44" />
                    <SPLIT distance="600" swimtime="00:08:08.32" />
                    <SPLIT distance="650" swimtime="00:08:50.56" />
                    <SPLIT distance="700" swimtime="00:09:32.78" />
                    <SPLIT distance="750" swimtime="00:10:15.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1279" points="399" swimtime="00:20:49.45" resultid="2868" heatid="5350" lane="7" entrytime="00:20:21.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:13.81" />
                    <SPLIT distance="150" swimtime="00:01:54.41" />
                    <SPLIT distance="200" swimtime="00:02:35.18" />
                    <SPLIT distance="250" swimtime="00:03:16.17" />
                    <SPLIT distance="300" swimtime="00:03:58.05" />
                    <SPLIT distance="350" swimtime="00:04:39.70" />
                    <SPLIT distance="400" swimtime="00:05:21.84" />
                    <SPLIT distance="450" swimtime="00:06:03.50" />
                    <SPLIT distance="500" swimtime="00:06:45.83" />
                    <SPLIT distance="550" swimtime="00:07:27.59" />
                    <SPLIT distance="600" swimtime="00:08:10.27" />
                    <SPLIT distance="650" swimtime="00:08:52.44" />
                    <SPLIT distance="700" swimtime="00:09:35.45" />
                    <SPLIT distance="750" swimtime="00:10:18.02" />
                    <SPLIT distance="800" swimtime="00:10:59.95" />
                    <SPLIT distance="850" swimtime="00:11:42.45" />
                    <SPLIT distance="900" swimtime="00:12:25.90" />
                    <SPLIT distance="950" swimtime="00:13:08.65" />
                    <SPLIT distance="1000" swimtime="00:13:51.25" />
                    <SPLIT distance="1050" swimtime="00:14:33.64" />
                    <SPLIT distance="1100" swimtime="00:15:15.87" />
                    <SPLIT distance="1150" swimtime="00:15:58.52" />
                    <SPLIT distance="1200" swimtime="00:16:40.26" />
                    <SPLIT distance="1250" swimtime="00:17:22.22" />
                    <SPLIT distance="1300" swimtime="00:18:03.84" />
                    <SPLIT distance="1350" swimtime="00:18:47.09" />
                    <SPLIT distance="1400" swimtime="00:19:28.52" />
                    <SPLIT distance="1450" swimtime="00:20:10.29" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietro" lastname="Lobo Mussoi" birthdate="2008-07-05" gender="M" nation="BRA" license="398573" swrid="5658061" athleteid="2869" externalid="398573">
              <RESULTS>
                <RESULT eventid="1104" points="485" swimtime="00:00:26.61" resultid="2870" heatid="5125" lane="8" entrytime="00:00:26.56" entrycourse="LCM" />
                <RESULT eventid="1167" points="486" swimtime="00:00:59.59" resultid="2871" heatid="5226" lane="2" entrytime="00:01:03.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="418" swimtime="00:00:31.48" resultid="2872" heatid="5285" lane="5" entrytime="00:00:33.05" entrycourse="LCM" />
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 10:33)" eventid="1267" status="DSQ" swimtime="00:00:28.53" resultid="2873" heatid="5334" lane="5" entrytime="00:00:29.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13068" nation="BRA" region="PR" clubid="4232" swrid="93787" name="Sociedade Morgenau" shortname="Morgenau">
          <ATHLETES>
            <ATHLETE firstname="Luana" lastname="Yoshie Kimura" birthdate="2010-07-08" gender="F" nation="BRA" license="391142" swrid="5600277" athleteid="4261" externalid="391142">
              <RESULTS>
                <RESULT eventid="1080" points="520" swimtime="00:01:19.72" resultid="4262" heatid="5067" lane="5" entrytime="00:01:20.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="408" swimtime="00:02:49.99" resultid="4263" heatid="5188" lane="1" entrytime="00:02:47.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                    <SPLIT distance="100" swimtime="00:01:24.99" />
                    <SPLIT distance="150" swimtime="00:02:11.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="385" swimtime="00:06:05.28" resultid="4264" heatid="5278" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.79" />
                    <SPLIT distance="100" swimtime="00:01:28.72" />
                    <SPLIT distance="150" swimtime="00:02:18.68" />
                    <SPLIT distance="200" swimtime="00:03:07.36" />
                    <SPLIT distance="250" swimtime="00:03:54.41" />
                    <SPLIT distance="300" swimtime="00:04:42.74" />
                    <SPLIT distance="350" swimtime="00:05:25.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="412" swimtime="00:03:04.76" resultid="4265" heatid="5313" lane="7" entrytime="00:03:00.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.28" />
                    <SPLIT distance="100" swimtime="00:01:28.65" />
                    <SPLIT distance="150" swimtime="00:02:17.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="528" swimtime="00:00:36.06" resultid="4266" heatid="5377" lane="7" entrytime="00:00:37.03" entrycourse="LCM" />
                <RESULT eventid="2312" points="499" swimtime="00:01:20.84" resultid="5944" heatid="6416" lane="7" entrytime="00:01:19.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabryel" lastname="Denk" birthdate="2011-05-09" gender="M" nation="BRA" license="391138" swrid="5602531" athleteid="4342" externalid="391138">
              <RESULTS>
                <RESULT eventid="1072" points="388" swimtime="00:05:01.60" resultid="4343" heatid="5058" lane="7" entrytime="00:05:01.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.55" />
                    <SPLIT distance="100" swimtime="00:01:09.97" />
                    <SPLIT distance="150" swimtime="00:01:48.57" />
                    <SPLIT distance="200" swimtime="00:02:27.60" />
                    <SPLIT distance="250" swimtime="00:03:06.42" />
                    <SPLIT distance="300" swimtime="00:03:45.79" />
                    <SPLIT distance="350" swimtime="00:04:24.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="346" swimtime="00:02:25.18" resultid="4344" heatid="5150" lane="8" entrytime="00:02:29.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.33" />
                    <SPLIT distance="100" swimtime="00:01:09.36" />
                    <SPLIT distance="150" swimtime="00:01:47.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="299" swimtime="00:01:17.10" resultid="4345" heatid="5256" lane="4" entrytime="00:01:19.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="279" swimtime="00:00:36.01" resultid="4346" heatid="5284" lane="5" entrytime="00:00:37.15" entrycourse="LCM" />
                <RESULT eventid="1217" points="372" swimtime="00:10:28.22" resultid="4347" heatid="5298" lane="4" entrytime="00:10:26.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.14" />
                    <SPLIT distance="100" swimtime="00:01:10.55" />
                    <SPLIT distance="150" swimtime="00:01:49.79" />
                    <SPLIT distance="200" swimtime="00:02:29.63" />
                    <SPLIT distance="250" swimtime="00:03:09.74" />
                    <SPLIT distance="300" swimtime="00:03:49.61" />
                    <SPLIT distance="350" swimtime="00:04:29.58" />
                    <SPLIT distance="400" swimtime="00:05:10.20" />
                    <SPLIT distance="450" swimtime="00:05:50.75" />
                    <SPLIT distance="500" swimtime="00:06:31.14" />
                    <SPLIT distance="550" swimtime="00:07:11.94" />
                    <SPLIT distance="600" swimtime="00:07:52.04" />
                    <SPLIT distance="650" swimtime="00:08:32.10" />
                    <SPLIT distance="700" swimtime="00:09:12.39" />
                    <SPLIT distance="750" swimtime="00:09:51.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="394" swimtime="00:19:47.66" resultid="4348" heatid="5379" lane="3" entrytime="00:19:50.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="100" swimtime="00:01:12.31" />
                    <SPLIT distance="150" swimtime="00:01:51.78" />
                    <SPLIT distance="200" swimtime="00:02:31.66" />
                    <SPLIT distance="250" swimtime="00:03:11.36" />
                    <SPLIT distance="300" swimtime="00:03:51.67" />
                    <SPLIT distance="350" swimtime="00:04:31.32" />
                    <SPLIT distance="400" swimtime="00:05:11.17" />
                    <SPLIT distance="450" swimtime="00:05:51.61" />
                    <SPLIT distance="500" swimtime="00:06:32.25" />
                    <SPLIT distance="550" swimtime="00:07:11.97" />
                    <SPLIT distance="600" swimtime="00:07:52.88" />
                    <SPLIT distance="650" swimtime="00:08:32.54" />
                    <SPLIT distance="700" swimtime="00:09:12.58" />
                    <SPLIT distance="750" swimtime="00:09:52.36" />
                    <SPLIT distance="800" swimtime="00:10:32.66" />
                    <SPLIT distance="850" swimtime="00:11:12.72" />
                    <SPLIT distance="900" swimtime="00:11:52.98" />
                    <SPLIT distance="950" swimtime="00:12:32.90" />
                    <SPLIT distance="1000" swimtime="00:13:12.92" />
                    <SPLIT distance="1050" swimtime="00:13:52.93" />
                    <SPLIT distance="1100" swimtime="00:14:32.73" />
                    <SPLIT distance="1150" swimtime="00:15:12.76" />
                    <SPLIT distance="1200" swimtime="00:15:52.62" />
                    <SPLIT distance="1250" swimtime="00:16:32.19" />
                    <SPLIT distance="1300" swimtime="00:17:12.10" />
                    <SPLIT distance="1350" swimtime="00:17:51.81" />
                    <SPLIT distance="1400" swimtime="00:18:31.25" />
                    <SPLIT distance="1450" swimtime="00:19:09.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Bora" birthdate="2005-01-06" gender="F" nation="BRA" license="358252" swrid="5600153" athleteid="4304" externalid="358252">
              <RESULTS>
                <RESULT eventid="1064" points="360" swimtime="00:05:30.82" resultid="4305" heatid="5055" lane="1" entrytime="00:05:37.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:17.46" />
                    <SPLIT distance="150" swimtime="00:01:59.81" />
                    <SPLIT distance="200" swimtime="00:02:41.67" />
                    <SPLIT distance="250" swimtime="00:03:24.22" />
                    <SPLIT distance="300" swimtime="00:04:06.65" />
                    <SPLIT distance="350" swimtime="00:04:49.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="341" swimtime="00:03:00.48" resultid="4306" heatid="5191" lane="6" entrytime="00:03:01.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                    <SPLIT distance="100" swimtime="00:01:23.30" />
                    <SPLIT distance="150" swimtime="00:02:20.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="309" swimtime="00:01:24.73" resultid="4307" heatid="5248" lane="2" entrytime="00:01:24.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="315" swimtime="00:06:30.45" resultid="4308" heatid="5279" lane="2" entrytime="00:06:48.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.97" />
                    <SPLIT distance="100" swimtime="00:01:25.58" />
                    <SPLIT distance="150" swimtime="00:02:17.40" />
                    <SPLIT distance="200" swimtime="00:03:07.14" />
                    <SPLIT distance="250" swimtime="00:04:06.31" />
                    <SPLIT distance="300" swimtime="00:05:03.91" />
                    <SPLIT distance="350" swimtime="00:05:47.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="261" swimtime="00:00:38.22" resultid="4309" heatid="5324" lane="1" entrytime="00:00:37.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Stella" lastname="Magalhaes Birnbaum" birthdate="2009-05-14" gender="F" nation="BRA" license="399684" swrid="5653298" athleteid="4378" externalid="399684">
              <RESULTS>
                <RESULT eventid="1096" points="412" swimtime="00:00:31.72" resultid="4379" heatid="5102" lane="7" entrytime="00:00:32.09" entrycourse="LCM" />
                <RESULT eventid="1175" points="342" swimtime="00:01:21.94" resultid="4380" heatid="5246" lane="5" entrytime="00:01:20.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="401" swimtime="00:01:10.11" resultid="4381" heatid="5207" lane="8" entrytime="00:01:09.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1275" points="341" swimtime="00:02:56.15" resultid="4382" heatid="5341" lane="1" entrytime="00:02:54.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.14" />
                    <SPLIT distance="100" swimtime="00:01:23.20" />
                    <SPLIT distance="150" swimtime="00:02:09.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Rafaella Dos Santos" birthdate="2005-02-25" gender="F" nation="BRA" license="358849" athleteid="4238" externalid="358849">
              <RESULTS>
                <RESULT eventid="1080" points="297" swimtime="00:01:36.10" resultid="4239" heatid="5070" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="263" swimtime="00:02:56.03" resultid="4240" heatid="5145" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.39" />
                    <SPLIT distance="100" swimtime="00:01:23.90" />
                    <SPLIT distance="150" swimtime="00:02:10.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="338" swimtime="00:00:41.85" resultid="4241" heatid="5373" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lauren" lastname="Dziura" birthdate="2010-01-11" gender="F" nation="BRA" license="369416" swrid="5588668" athleteid="4315" externalid="369416">
              <RESULTS>
                <RESULT eventid="1064" points="403" swimtime="00:05:18.55" resultid="4316" heatid="5050" lane="8" entrytime="00:05:13.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.33" />
                    <SPLIT distance="100" swimtime="00:01:14.18" />
                    <SPLIT distance="150" swimtime="00:01:52.98" />
                    <SPLIT distance="200" swimtime="00:02:33.11" />
                    <SPLIT distance="250" swimtime="00:03:13.73" />
                    <SPLIT distance="300" swimtime="00:03:56.62" />
                    <SPLIT distance="350" swimtime="00:04:38.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="400" swimtime="00:00:32.04" resultid="4317" heatid="5098" lane="2" entrytime="00:00:32.76" entrycourse="LCM" />
                <RESULT eventid="1112" points="424" swimtime="00:02:30.14" resultid="4318" heatid="5140" lane="2" entrytime="00:02:28.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.58" />
                    <SPLIT distance="100" swimtime="00:01:14.18" />
                    <SPLIT distance="150" swimtime="00:01:52.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="406" swimtime="00:10:54.27" resultid="4319" heatid="5271" lane="1" entrytime="00:10:59.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                    <SPLIT distance="100" swimtime="00:01:16.32" />
                    <SPLIT distance="150" swimtime="00:01:56.30" />
                    <SPLIT distance="200" swimtime="00:02:37.34" />
                    <SPLIT distance="250" swimtime="00:03:18.92" />
                    <SPLIT distance="300" swimtime="00:03:59.58" />
                    <SPLIT distance="350" swimtime="00:04:41.97" />
                    <SPLIT distance="400" swimtime="00:05:23.89" />
                    <SPLIT distance="450" swimtime="00:06:06.71" />
                    <SPLIT distance="500" swimtime="00:06:48.51" />
                    <SPLIT distance="550" swimtime="00:07:29.89" />
                    <SPLIT distance="600" swimtime="00:08:11.90" />
                    <SPLIT distance="650" swimtime="00:08:53.69" />
                    <SPLIT distance="700" swimtime="00:09:34.40" />
                    <SPLIT distance="750" swimtime="00:10:15.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="346" swimtime="00:06:18.50" resultid="4320" heatid="5279" lane="7" entrytime="00:06:51.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.41" />
                    <SPLIT distance="100" swimtime="00:01:27.96" />
                    <SPLIT distance="150" swimtime="00:02:17.68" />
                    <SPLIT distance="200" swimtime="00:03:05.38" />
                    <SPLIT distance="250" swimtime="00:04:01.74" />
                    <SPLIT distance="300" swimtime="00:04:57.06" />
                    <SPLIT distance="350" swimtime="00:05:39.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1279" points="420" swimtime="00:20:28.45" resultid="4321" heatid="5349" lane="4" entrytime="00:20:47.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.89" />
                    <SPLIT distance="100" swimtime="00:01:15.91" />
                    <SPLIT distance="150" swimtime="00:01:56.28" />
                    <SPLIT distance="200" swimtime="00:02:36.96" />
                    <SPLIT distance="250" swimtime="00:03:18.26" />
                    <SPLIT distance="300" swimtime="00:03:59.12" />
                    <SPLIT distance="350" swimtime="00:04:39.35" />
                    <SPLIT distance="400" swimtime="00:05:19.57" />
                    <SPLIT distance="450" swimtime="00:06:00.24" />
                    <SPLIT distance="500" swimtime="00:06:40.24" />
                    <SPLIT distance="550" swimtime="00:07:20.94" />
                    <SPLIT distance="600" swimtime="00:08:02.20" />
                    <SPLIT distance="650" swimtime="00:08:43.65" />
                    <SPLIT distance="700" swimtime="00:09:24.40" />
                    <SPLIT distance="750" swimtime="00:10:06.04" />
                    <SPLIT distance="800" swimtime="00:10:47.77" />
                    <SPLIT distance="850" swimtime="00:11:29.65" />
                    <SPLIT distance="900" swimtime="00:12:11.36" />
                    <SPLIT distance="950" swimtime="00:12:52.96" />
                    <SPLIT distance="1000" swimtime="00:13:34.29" />
                    <SPLIT distance="1050" swimtime="00:14:16.12" />
                    <SPLIT distance="1100" swimtime="00:14:57.68" />
                    <SPLIT distance="1150" swimtime="00:15:38.82" />
                    <SPLIT distance="1200" swimtime="00:16:20.13" />
                    <SPLIT distance="1250" swimtime="00:17:01.91" />
                    <SPLIT distance="1300" swimtime="00:17:44.44" />
                    <SPLIT distance="1350" swimtime="00:18:26.72" />
                    <SPLIT distance="1400" swimtime="00:19:08.88" />
                    <SPLIT distance="1450" swimtime="00:19:49.54" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wilson" lastname="Soares Filho" birthdate="2007-12-20" gender="M" nation="BRA" license="414552" swrid="5755379" athleteid="4402" externalid="414552">
              <RESULTS>
                <RESULT eventid="1088" points="284" swimtime="00:01:26.44" resultid="4403" heatid="5086" lane="2" entrytime="00:01:29.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="361" swimtime="00:01:05.76" resultid="4404" heatid="5231" lane="7" entrytime="00:01:07.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="361" swimtime="00:00:36.42" resultid="4405" heatid="5367" lane="4" entrytime="00:00:38.08" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marcus" lastname="Vinicius De Almeida" birthdate="2009-06-16" gender="M" nation="BRA" license="348099" swrid="5600272" athleteid="4297" externalid="348099">
              <RESULTS>
                <RESULT eventid="1088" points="524" swimtime="00:01:10.52" resultid="4298" heatid="5085" lane="2" entrytime="00:01:09.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="457" swimtime="00:02:27.97" resultid="4299" heatid="5198" lane="1" entrytime="00:02:25.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:11.48" />
                    <SPLIT distance="150" swimtime="00:01:52.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="475" swimtime="00:01:06.10" resultid="4300" heatid="5261" lane="1" entrytime="00:01:06.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.01" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 8.3 - Movimento alternado das pernas ou pés.  (Horário: 16:50)" eventid="1198" status="DSQ" swimtime="00:05:17.49" resultid="4301" heatid="5275" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.31" />
                    <SPLIT distance="100" swimtime="00:01:15.32" />
                    <SPLIT distance="150" swimtime="00:01:57.43" />
                    <SPLIT distance="200" swimtime="00:02:39.36" />
                    <SPLIT distance="250" swimtime="00:03:22.21" />
                    <SPLIT distance="300" swimtime="00:04:05.73" />
                    <SPLIT distance="350" swimtime="00:04:42.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="458" swimtime="00:00:30.55" resultid="4302" heatid="5287" lane="7" entrytime="00:00:30.31" entrycourse="LCM" />
                <RESULT eventid="1297" points="545" swimtime="00:00:31.76" resultid="4303" heatid="5370" lane="4" entrytime="00:00:31.97" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Barros Zagonel" birthdate="2006-06-01" gender="M" nation="BRA" license="347856" swrid="5622261" athleteid="4233" externalid="347856" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1088" points="297" swimtime="00:01:25.23" resultid="4234" heatid="5086" lane="3" entrytime="00:01:23.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="314" swimtime="00:02:47.72" resultid="4235" heatid="5200" lane="1" entrytime="00:02:50.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:20.24" />
                    <SPLIT distance="150" swimtime="00:02:09.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="289" swimtime="00:03:09.77" resultid="4236" heatid="5317" lane="2" entrytime="00:03:08.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                    <SPLIT distance="100" swimtime="00:01:27.67" />
                    <SPLIT distance="150" swimtime="00:02:18.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="376" swimtime="00:00:35.95" resultid="4237" heatid="5369" lane="1" entrytime="00:00:35.42" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benito" lastname="Alves Sant&apos;Ana" birthdate="2009-06-01" gender="M" nation="BRA" license="376585" swrid="5351951" athleteid="4254" externalid="376585">
              <RESULTS>
                <RESULT eventid="1072" points="525" swimtime="00:04:32.78" resultid="4255" heatid="5062" lane="7" entrytime="00:04:28.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.86" />
                    <SPLIT distance="100" swimtime="00:01:04.75" />
                    <SPLIT distance="150" swimtime="00:01:39.42" />
                    <SPLIT distance="200" swimtime="00:02:14.27" />
                    <SPLIT distance="250" swimtime="00:02:49.19" />
                    <SPLIT distance="300" swimtime="00:03:25.02" />
                    <SPLIT distance="350" swimtime="00:04:00.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="457" swimtime="00:02:27.99" resultid="4256" heatid="5197" lane="6" entrytime="00:02:28.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:09.44" />
                    <SPLIT distance="150" swimtime="00:01:56.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="483" swimtime="00:05:09.06" resultid="4257" heatid="5277" lane="1" entrytime="00:05:10.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.01" />
                    <SPLIT distance="100" swimtime="00:01:10.12" />
                    <SPLIT distance="150" swimtime="00:01:50.45" />
                    <SPLIT distance="200" swimtime="00:02:29.52" />
                    <SPLIT distance="250" swimtime="00:03:16.33" />
                    <SPLIT distance="300" swimtime="00:04:01.51" />
                    <SPLIT distance="350" swimtime="00:04:36.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="515" swimtime="00:09:24.01" resultid="4258" heatid="5300" lane="5" entrytime="00:09:08.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.93" />
                    <SPLIT distance="100" swimtime="00:01:04.65" />
                    <SPLIT distance="150" swimtime="00:01:40.03" />
                    <SPLIT distance="200" swimtime="00:02:14.99" />
                    <SPLIT distance="250" swimtime="00:02:51.12" />
                    <SPLIT distance="300" swimtime="00:03:26.89" />
                    <SPLIT distance="350" swimtime="00:04:03.28" />
                    <SPLIT distance="400" swimtime="00:04:39.14" />
                    <SPLIT distance="450" swimtime="00:05:15.64" />
                    <SPLIT distance="500" swimtime="00:05:51.84" />
                    <SPLIT distance="550" swimtime="00:06:28.56" />
                    <SPLIT distance="600" swimtime="00:07:02.92" />
                    <SPLIT distance="650" swimtime="00:07:40.09" />
                    <SPLIT distance="700" swimtime="00:08:15.87" />
                    <SPLIT distance="750" swimtime="00:08:51.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="424" swimtime="00:02:28.97" resultid="4259" heatid="5346" lane="2" entrytime="00:02:33.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.82" />
                    <SPLIT distance="100" swimtime="00:01:12.45" />
                    <SPLIT distance="150" swimtime="00:01:51.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="551" swimtime="00:17:41.90" resultid="4260" heatid="5380" lane="4" entrytime="00:17:25.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.66" />
                    <SPLIT distance="100" swimtime="00:01:04.33" />
                    <SPLIT distance="150" swimtime="00:01:39.11" />
                    <SPLIT distance="200" swimtime="00:02:14.15" />
                    <SPLIT distance="250" swimtime="00:02:50.22" />
                    <SPLIT distance="300" swimtime="00:03:26.12" />
                    <SPLIT distance="350" swimtime="00:04:02.42" />
                    <SPLIT distance="400" swimtime="00:04:37.99" />
                    <SPLIT distance="450" swimtime="00:05:14.26" />
                    <SPLIT distance="500" swimtime="00:05:49.74" />
                    <SPLIT distance="550" swimtime="00:06:25.73" />
                    <SPLIT distance="600" swimtime="00:07:00.20" />
                    <SPLIT distance="650" swimtime="00:07:35.48" />
                    <SPLIT distance="700" swimtime="00:08:11.02" />
                    <SPLIT distance="750" swimtime="00:08:46.65" />
                    <SPLIT distance="800" swimtime="00:09:22.60" />
                    <SPLIT distance="850" swimtime="00:09:58.51" />
                    <SPLIT distance="900" swimtime="00:10:34.70" />
                    <SPLIT distance="950" swimtime="00:11:10.47" />
                    <SPLIT distance="1000" swimtime="00:11:46.32" />
                    <SPLIT distance="1050" swimtime="00:12:22.43" />
                    <SPLIT distance="1100" swimtime="00:12:58.55" />
                    <SPLIT distance="1150" swimtime="00:13:34.11" />
                    <SPLIT distance="1200" swimtime="00:14:09.95" />
                    <SPLIT distance="1250" swimtime="00:14:46.13" />
                    <SPLIT distance="1300" swimtime="00:15:22.47" />
                    <SPLIT distance="1350" swimtime="00:15:58.24" />
                    <SPLIT distance="1400" swimtime="00:16:33.77" />
                    <SPLIT distance="1450" swimtime="00:17:08.45" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Mingorance Martins" birthdate="2007-10-13" gender="M" nation="BRA" license="393920" swrid="5622295" athleteid="4364" externalid="393920">
              <RESULTS>
                <RESULT eventid="1072" points="462" swimtime="00:04:44.64" resultid="4365" heatid="5064" lane="7" entrytime="00:04:46.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                    <SPLIT distance="100" swimtime="00:01:04.07" />
                    <SPLIT distance="150" swimtime="00:01:39.27" />
                    <SPLIT distance="200" swimtime="00:02:16.06" />
                    <SPLIT distance="250" swimtime="00:02:53.33" />
                    <SPLIT distance="300" swimtime="00:03:30.77" />
                    <SPLIT distance="350" swimtime="00:04:08.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="508" swimtime="00:00:26.20" resultid="4366" heatid="5129" lane="8" entrytime="00:00:25.92" entrycourse="LCM" />
                <RESULT eventid="1120" points="502" swimtime="00:02:08.32" resultid="4367" heatid="5158" lane="1" entrytime="00:02:09.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.64" />
                    <SPLIT distance="100" swimtime="00:01:00.52" />
                    <SPLIT distance="150" swimtime="00:01:34.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="365" swimtime="00:01:12.18" resultid="4368" heatid="5262" lane="6" entrytime="00:01:12.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="558" swimtime="00:00:56.90" resultid="4369" heatid="5232" lane="7" entrytime="00:00:57.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="378" swimtime="00:02:34.70" resultid="4370" heatid="5345" lane="5" entrytime="00:02:39.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:14.42" />
                    <SPLIT distance="150" swimtime="00:01:54.87" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thiago" lastname="Kozera Chiarato" birthdate="2008-01-22" gender="M" nation="BRA" license="406728" swrid="5717276" athleteid="4395" externalid="406728">
              <RESULTS>
                <RESULT eventid="1088" points="394" swimtime="00:01:17.54" resultid="4396" heatid="5084" lane="2" entrytime="00:01:18.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="423" swimtime="00:00:27.85" resultid="4397" heatid="5123" lane="3" entrytime="00:00:27.77" entrycourse="LCM" />
                <RESULT eventid="1135" points="358" swimtime="00:01:09.64" resultid="4398" heatid="5173" lane="4" entrytime="00:01:09.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="460" swimtime="00:01:00.69" resultid="4399" heatid="5227" lane="6" entrytime="00:01:00.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="344" swimtime="00:00:31.76" resultid="4400" heatid="5332" lane="2" entrytime="00:00:32.70" entrycourse="LCM" />
                <RESULT eventid="1297" points="403" swimtime="00:00:35.13" resultid="4401" heatid="5365" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaylane" lastname="Marques Ferreira" birthdate="2010-03-06" gender="F" nation="BRA" license="391146" swrid="5600211" athleteid="4356" externalid="391146">
              <RESULTS>
                <RESULT eventid="1064" points="233" swimtime="00:06:22.07" resultid="4357" heatid="5048" lane="5" entrytime="00:06:30.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                    <SPLIT distance="100" swimtime="00:01:22.80" />
                    <SPLIT distance="150" swimtime="00:02:13.23" />
                    <SPLIT distance="200" swimtime="00:03:00.97" />
                    <SPLIT distance="250" swimtime="00:03:53.33" />
                    <SPLIT distance="300" swimtime="00:04:45.49" />
                    <SPLIT distance="350" swimtime="00:05:35.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="305" swimtime="00:00:35.04" resultid="4358" heatid="5097" lane="5" entrytime="00:00:34.55" entrycourse="LCM" />
                <RESULT eventid="1128" points="198" swimtime="00:01:35.11" resultid="4359" heatid="5160" lane="8" entrytime="00:01:27.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="300" swimtime="00:01:17.16" resultid="4360" heatid="5201" lane="4" entrytime="00:01:19.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="351" swimtime="00:00:34.60" resultid="4361" heatid="5325" lane="2" entrytime="00:00:34.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="Rodrigues Galvao" birthdate="2007-04-19" gender="M" nation="BRA" license="376586" swrid="5600247" athleteid="4248" externalid="376586">
              <RESULTS>
                <RESULT eventid="1104" points="524" swimtime="00:00:25.92" resultid="4249" heatid="5128" lane="4" entrytime="00:00:26.07" entrycourse="LCM" />
                <RESULT eventid="1135" points="480" swimtime="00:01:03.13" resultid="4250" heatid="5177" lane="1" entrytime="00:01:03.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="524" swimtime="00:00:58.11" resultid="4251" heatid="5232" lane="1" entrytime="00:00:58.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="520" swimtime="00:00:27.68" resultid="4252" heatid="5336" lane="3" entrytime="00:00:27.65" entrycourse="LCM" />
                <RESULT eventid="1293" points="371" swimtime="00:02:33.44" resultid="4253" heatid="5359" lane="7" entrytime="00:02:35.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:07.96" />
                    <SPLIT distance="150" swimtime="00:01:48.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monike" lastname="Lemos Carvalho" birthdate="2008-03-28" gender="F" nation="BRA" license="307796" swrid="5600199" athleteid="4338" externalid="307796">
              <RESULTS>
                <RESULT eventid="1064" points="384" swimtime="00:05:23.56" resultid="4339" heatid="5053" lane="2" entrytime="00:05:18.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.95" />
                    <SPLIT distance="100" swimtime="00:01:11.76" />
                    <SPLIT distance="150" swimtime="00:01:52.23" />
                    <SPLIT distance="200" swimtime="00:02:33.70" />
                    <SPLIT distance="250" swimtime="00:03:16.43" />
                    <SPLIT distance="300" swimtime="00:03:59.02" />
                    <SPLIT distance="350" swimtime="00:04:42.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="460" swimtime="00:00:30.57" resultid="4340" heatid="5101" lane="6" />
                <RESULT eventid="1112" points="479" swimtime="00:02:24.20" resultid="4341" heatid="5144" lane="8" entrytime="00:02:24.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.92" />
                    <SPLIT distance="100" swimtime="00:01:09.07" />
                    <SPLIT distance="150" swimtime="00:01:47.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Gabriel Sarmento Buski" birthdate="2010-04-05" gender="M" nation="BRA" license="399533" swrid="5717264" athleteid="4267" externalid="399533">
              <RESULTS>
                <RESULT eventid="1088" points="335" swimtime="00:01:21.86" resultid="4268" heatid="5082" lane="3" entrytime="00:01:18.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="364" swimtime="00:05:08.20" resultid="4269" heatid="5058" lane="2" entrytime="00:05:00.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.60" />
                    <SPLIT distance="100" swimtime="00:01:10.94" />
                    <SPLIT distance="150" swimtime="00:01:50.05" />
                    <SPLIT distance="200" swimtime="00:02:29.26" />
                    <SPLIT distance="250" swimtime="00:03:10.29" />
                    <SPLIT distance="300" swimtime="00:03:50.22" />
                    <SPLIT distance="350" swimtime="00:04:30.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="300" swimtime="00:02:32.34" resultid="4270" heatid="5149" lane="3" entrytime="00:02:36.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:12.60" />
                    <SPLIT distance="150" swimtime="00:01:52.82" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="346" swimtime="00:10:43.93" resultid="4271" heatid="5299" lane="8" entrytime="00:10:22.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.32" />
                    <SPLIT distance="100" swimtime="00:01:11.52" />
                    <SPLIT distance="150" swimtime="00:01:51.76" />
                    <SPLIT distance="200" swimtime="00:02:32.32" />
                    <SPLIT distance="250" swimtime="00:03:13.24" />
                    <SPLIT distance="300" swimtime="00:03:54.32" />
                    <SPLIT distance="350" swimtime="00:04:34.67" />
                    <SPLIT distance="400" swimtime="00:05:16.42" />
                    <SPLIT distance="450" swimtime="00:05:57.45" />
                    <SPLIT distance="500" swimtime="00:06:38.13" />
                    <SPLIT distance="550" swimtime="00:07:19.36" />
                    <SPLIT distance="600" swimtime="00:08:00.56" />
                    <SPLIT distance="650" swimtime="00:08:41.51" />
                    <SPLIT distance="700" swimtime="00:09:23.19" />
                    <SPLIT distance="750" swimtime="00:10:03.54" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 9:50), Na volta dos 100m." eventid="1251" status="DSQ" swimtime="00:03:00.50" resultid="4272" heatid="5316" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                    <SPLIT distance="100" swimtime="00:01:23.52" />
                    <SPLIT distance="150" swimtime="00:02:12.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="363" swimtime="00:20:20.09" resultid="4273" heatid="5379" lane="5" entrytime="00:19:48.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:01:13.48" />
                    <SPLIT distance="150" swimtime="00:01:53.46" />
                    <SPLIT distance="200" swimtime="00:02:34.62" />
                    <SPLIT distance="250" swimtime="00:03:14.81" />
                    <SPLIT distance="300" swimtime="00:03:56.04" />
                    <SPLIT distance="350" swimtime="00:04:37.61" />
                    <SPLIT distance="400" swimtime="00:05:18.69" />
                    <SPLIT distance="450" swimtime="00:06:00.63" />
                    <SPLIT distance="500" swimtime="00:06:41.74" />
                    <SPLIT distance="550" swimtime="00:07:23.47" />
                    <SPLIT distance="600" swimtime="00:08:04.56" />
                    <SPLIT distance="650" swimtime="00:08:47.52" />
                    <SPLIT distance="700" swimtime="00:09:28.88" />
                    <SPLIT distance="750" swimtime="00:10:11.22" />
                    <SPLIT distance="800" swimtime="00:10:52.58" />
                    <SPLIT distance="850" swimtime="00:11:32.96" />
                    <SPLIT distance="900" swimtime="00:12:12.80" />
                    <SPLIT distance="950" swimtime="00:12:52.52" />
                    <SPLIT distance="1000" swimtime="00:13:32.26" />
                    <SPLIT distance="1050" swimtime="00:14:13.10" />
                    <SPLIT distance="1100" swimtime="00:14:53.95" />
                    <SPLIT distance="1150" swimtime="00:15:34.02" />
                    <SPLIT distance="1200" swimtime="00:16:15.20" />
                    <SPLIT distance="1250" swimtime="00:16:57.20" />
                    <SPLIT distance="1300" swimtime="00:17:39.30" />
                    <SPLIT distance="1350" swimtime="00:18:20.83" />
                    <SPLIT distance="1400" swimtime="00:19:02.04" />
                    <SPLIT distance="1450" swimtime="00:19:41.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Kozera Chiarato" birthdate="2010-05-28" gender="M" nation="BRA" license="406722" swrid="5717275" athleteid="4388" externalid="406722">
              <RESULTS>
                <RESULT eventid="1104" points="324" swimtime="00:00:30.43" resultid="4389" heatid="5117" lane="3" entrytime="00:00:30.38" entrycourse="LCM" />
                <RESULT eventid="1135" points="303" swimtime="00:01:13.56" resultid="4390" heatid="5170" lane="5" entrytime="00:01:16.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="282" swimtime="00:02:53.81" resultid="4391" heatid="5193" lane="5" entrytime="00:02:54.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.39" />
                    <SPLIT distance="100" swimtime="00:01:25.52" />
                    <SPLIT distance="150" swimtime="00:02:18.33" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="313" swimtime="00:01:08.97" resultid="4392" heatid="5220" lane="1" entrytime="00:01:08.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="301" swimtime="00:00:33.21" resultid="4393" heatid="5332" lane="1" entrytime="00:00:33.59" entrycourse="LCM" />
                <RESULT eventid="1293" points="217" swimtime="00:03:03.59" resultid="4394" heatid="5358" lane="1" entrytime="00:03:03.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.40" />
                    <SPLIT distance="100" swimtime="00:01:26.29" />
                    <SPLIT distance="150" swimtime="00:02:16.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Geovana" lastname="Dos Santos" birthdate="2011-01-20" gender="F" nation="BRA" license="367254" swrid="5602533" athleteid="4242" externalid="367254">
              <RESULTS>
                <RESULT eventid="1096" points="321" swimtime="00:00:34.47" resultid="4243" heatid="5097" lane="3" entrytime="00:00:34.62" entrycourse="LCM" />
                <RESULT eventid="1175" points="308" swimtime="00:01:24.86" resultid="4244" heatid="5242" lane="6" entrytime="00:01:26.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="309" swimtime="00:01:16.41" resultid="4245" heatid="5202" lane="6" entrytime="00:01:15.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="320" swimtime="00:00:39.25" resultid="4246" heatid="5293" lane="1" entrytime="00:00:40.67" entrycourse="LCM" />
                <RESULT eventid="1275" points="281" swimtime="00:03:07.91" resultid="4247" heatid="5340" lane="6" entrytime="00:03:02.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                    <SPLIT distance="100" swimtime="00:01:29.85" />
                    <SPLIT distance="150" swimtime="00:02:19.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Andreis Ramos" birthdate="2007-03-26" gender="M" nation="BRA" license="406719" swrid="5717243" athleteid="4290" externalid="406719">
              <RESULTS>
                <RESULT eventid="1104" points="413" swimtime="00:00:28.07" resultid="4291" heatid="5127" lane="5" entrytime="00:00:28.31" entrycourse="LCM" />
                <RESULT eventid="1135" points="267" swimtime="00:01:16.79" resultid="4292" heatid="5176" lane="3" entrytime="00:01:18.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="359" swimtime="00:02:23.44" resultid="4293" heatid="5157" lane="5" entrytime="00:02:25.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.75" />
                    <SPLIT distance="100" swimtime="00:01:07.69" />
                    <SPLIT distance="150" swimtime="00:01:46.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="410" swimtime="00:01:03.03" resultid="4294" heatid="5231" lane="6" entrytime="00:01:03.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="275" swimtime="00:00:36.18" resultid="4295" heatid="5284" lane="4" entrytime="00:00:36.36" entrycourse="LCM" />
                <RESULT eventid="1267" points="332" swimtime="00:00:32.13" resultid="4296" heatid="5333" lane="7" entrytime="00:00:31.35" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Luiza Rimbano De Jesus" birthdate="2008-09-02" gender="F" nation="BRA" license="366819" swrid="5653297" athleteid="4371" externalid="366819">
              <RESULTS>
                <RESULT eventid="1096" points="573" swimtime="00:00:28.41" resultid="4372" heatid="5104" lane="5" entrytime="00:00:28.21" entrycourse="LCM" />
                <RESULT eventid="1112" points="468" swimtime="00:02:25.35" resultid="4373" heatid="5144" lane="7" entrytime="00:02:23.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.58" />
                    <SPLIT distance="100" swimtime="00:01:08.32" />
                    <SPLIT distance="150" swimtime="00:01:47.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="554" swimtime="00:01:02.96" resultid="4374" heatid="5208" lane="2" entrytime="00:01:02.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="437" swimtime="00:00:35.37" resultid="4375" heatid="5289" lane="4" />
                <RESULT eventid="1259" points="397" swimtime="00:00:33.22" resultid="4376" heatid="5325" lane="8" entrytime="00:00:35.69" entrycourse="LCM" />
                <RESULT eventid="1305" points="472" swimtime="00:00:37.45" resultid="4377" heatid="5376" lane="3" entrytime="00:00:38.24" entrycourse="LCM" />
                <RESULT eventid="2375" points="554" swimtime="00:00:28.73" resultid="5971" heatid="5978" lane="6" entrytime="00:00:28.41" />
                <RESULT eventid="2343" points="534" swimtime="00:01:03.70" resultid="6106" heatid="6421" lane="7" entrytime="00:01:02.96">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Andrianczik Corcini" birthdate="2008-07-19" gender="M" nation="BRA" license="406685" swrid="5736533" athleteid="4274" externalid="406685">
              <RESULTS>
                <RESULT eventid="1088" points="257" swimtime="00:01:29.44" resultid="4275" heatid="5083" lane="6" entrytime="00:01:33.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="343" swimtime="00:00:29.87" resultid="4276" heatid="5122" lane="1" entrytime="00:00:29.55" entrycourse="LCM" />
                <RESULT eventid="1167" points="333" swimtime="00:01:07.60" resultid="4277" heatid="5225" lane="8" entrytime="00:01:08.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" status="SICK" swimtime="00:00:00.00" resultid="4278" heatid="5366" lane="5" entrytime="00:00:41.28" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Lima" birthdate="2006-12-03" gender="M" nation="BRA" license="366749" swrid="5600201" athleteid="4322" externalid="366749">
              <RESULTS>
                <RESULT eventid="1104" points="550" swimtime="00:00:25.51" resultid="4323" heatid="5129" lane="2" entrytime="00:00:25.27" entrycourse="LCM" />
                <RESULT eventid="1135" points="487" swimtime="00:01:02.81" resultid="4324" heatid="5177" lane="2" entrytime="00:01:02.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="583" swimtime="00:00:56.07" resultid="4325" heatid="5232" lane="3" entrytime="00:00:55.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="537" swimtime="00:00:27.39" resultid="4326" heatid="5337" lane="7" entrytime="00:00:27.31" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Fernanda Pinto" birthdate="2004-09-17" gender="F" nation="BRA" license="391144" swrid="5600157" athleteid="4284" externalid="391144">
              <RESULTS>
                <RESULT eventid="1096" points="397" swimtime="00:00:32.10" resultid="4285" heatid="5106" lane="1" entrytime="00:00:32.41" entrycourse="LCM" />
                <RESULT eventid="1112" points="318" swimtime="00:02:45.23" resultid="4286" heatid="5146" lane="8" entrytime="00:02:46.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.07" />
                    <SPLIT distance="100" swimtime="00:01:17.11" />
                    <SPLIT distance="150" swimtime="00:02:01.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="356" swimtime="00:01:12.96" resultid="4287" heatid="5209" lane="2" entrytime="00:01:11.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="294" swimtime="00:00:40.35" resultid="4288" heatid="5293" lane="8" entrytime="00:00:40.76" entrycourse="LCM" />
                <RESULT eventid="1259" points="223" swimtime="00:00:40.23" resultid="4289" heatid="5323" lane="4" entrytime="00:00:38.69" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauan" lastname="Araujo" birthdate="2009-12-17" gender="M" nation="BRA" license="385119" swrid="5653286" athleteid="4332" externalid="385119">
              <RESULTS>
                <RESULT eventid="1104" points="352" swimtime="00:00:29.60" resultid="4333" heatid="5122" lane="2" entrytime="00:00:29.07" entrycourse="LCM" />
                <RESULT eventid="1120" points="383" swimtime="00:02:20.45" resultid="4334" heatid="5153" lane="3" entrytime="00:02:24.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.73" />
                    <SPLIT distance="100" swimtime="00:01:05.93" />
                    <SPLIT distance="150" swimtime="00:01:42.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="308" swimtime="00:02:48.74" resultid="4335" heatid="5197" lane="1" entrytime="00:02:44.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.09" />
                    <SPLIT distance="100" swimtime="00:01:18.76" />
                    <SPLIT distance="150" swimtime="00:02:12.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="392" swimtime="00:01:04.01" resultid="4336" heatid="5226" lane="8" entrytime="00:01:03.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="359" swimtime="00:10:35.66" resultid="4337" heatid="5298" lane="5" entrytime="00:10:32.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:11.34" />
                    <SPLIT distance="150" swimtime="00:01:50.82" />
                    <SPLIT distance="200" swimtime="00:02:30.49" />
                    <SPLIT distance="250" swimtime="00:03:11.06" />
                    <SPLIT distance="300" swimtime="00:03:52.01" />
                    <SPLIT distance="350" swimtime="00:04:32.18" />
                    <SPLIT distance="400" swimtime="00:05:13.51" />
                    <SPLIT distance="450" swimtime="00:05:54.19" />
                    <SPLIT distance="500" swimtime="00:06:35.68" />
                    <SPLIT distance="550" swimtime="00:07:16.76" />
                    <SPLIT distance="600" swimtime="00:07:58.02" />
                    <SPLIT distance="650" swimtime="00:08:38.74" />
                    <SPLIT distance="700" swimtime="00:09:19.36" />
                    <SPLIT distance="750" swimtime="00:09:58.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduarda" lastname="Azevedo Birsneek" birthdate="2010-03-31" gender="F" nation="BRA" license="391145" swrid="5389427" athleteid="4349" externalid="391145">
              <RESULTS>
                <RESULT eventid="1064" points="189" swimtime="00:06:49.94" resultid="4350" heatid="5048" lane="3" entrytime="00:06:51.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.77" />
                    <SPLIT distance="100" swimtime="00:01:33.85" />
                    <SPLIT distance="150" swimtime="00:02:26.34" />
                    <SPLIT distance="250" swimtime="00:04:11.46" />
                    <SPLIT distance="300" swimtime="00:05:04.57" />
                    <SPLIT distance="350" swimtime="00:05:58.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="221" swimtime="00:00:39.05" resultid="4351" heatid="5096" lane="7" entrytime="00:00:39.38" entrycourse="LCM" />
                <RESULT eventid="1128" points="135" swimtime="00:01:47.97" resultid="4352" heatid="5159" lane="7" entrytime="00:01:45.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="228" swimtime="00:00:43.93" resultid="4353" heatid="5291" lane="3" entrytime="00:00:45.37" entrycourse="LCM" />
                <RESULT eventid="1259" points="136" swimtime="00:00:47.45" resultid="4354" heatid="5322" lane="4" entrytime="00:00:49.44" entrycourse="LCM" />
                <RESULT eventid="1275" points="221" swimtime="00:03:23.39" resultid="4355" heatid="5340" lane="8" entrytime="00:03:31.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.96" />
                    <SPLIT distance="150" swimtime="00:02:33.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Henrique Opuchkevich" birthdate="2011-02-22" gender="M" nation="BRA" license="406720" swrid="5717273" athleteid="4383" externalid="406720">
              <RESULTS>
                <RESULT eventid="1088" points="311" swimtime="00:01:23.93" resultid="4384" heatid="5081" lane="5" entrytime="00:01:26.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="369" swimtime="00:05:06.59" resultid="4385" heatid="5057" lane="3" entrytime="00:05:15.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.76" />
                    <SPLIT distance="100" swimtime="00:01:09.72" />
                    <SPLIT distance="150" swimtime="00:01:49.55" />
                    <SPLIT distance="200" swimtime="00:02:28.75" />
                    <SPLIT distance="250" swimtime="00:03:09.76" />
                    <SPLIT distance="300" swimtime="00:03:49.71" />
                    <SPLIT distance="350" swimtime="00:04:29.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="316" swimtime="00:03:04.13" resultid="4386" heatid="5317" lane="6" entrytime="00:03:06.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.76" />
                    <SPLIT distance="100" swimtime="00:01:26.86" />
                    <SPLIT distance="150" swimtime="00:02:15.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="344" swimtime="00:00:37.02" resultid="4387" heatid="5367" lane="6" entrytime="00:00:40.14" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mayara" lastname="Fieber" birthdate="2008-08-20" gender="F" nation="BRA" license="391147" swrid="5600161" athleteid="4362" externalid="391147">
              <RESULTS>
                <RESULT eventid="1259" points="329" swimtime="00:00:35.36" resultid="4363" heatid="5321" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Karine" lastname="Correa" birthdate="2002-08-01" gender="F" nation="BRA" license="385191" swrid="5600141" athleteid="4279" externalid="385191">
              <RESULTS>
                <RESULT eventid="1064" points="324" swimtime="00:05:42.57" resultid="4280" heatid="5054" lane="4" entrytime="00:05:44.91" entrycourse="LCM" />
                <RESULT eventid="1096" points="393" swimtime="00:00:32.22" resultid="4281" heatid="5105" lane="3" />
                <RESULT eventid="1112" points="333" swimtime="00:02:42.67" resultid="4282" heatid="5146" lane="1" entrytime="00:02:43.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:17.20" />
                    <SPLIT distance="150" swimtime="00:02:00.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="278" swimtime="00:03:13.03" resultid="4283" heatid="5191" lane="2" entrytime="00:03:12.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.45" />
                    <SPLIT distance="100" swimtime="00:01:30.91" />
                    <SPLIT distance="150" swimtime="00:02:30.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Vitor Navarro Zanini" birthdate="2008-06-30" gender="M" nation="BRA" license="369415" swrid="5600273" athleteid="4310" externalid="369415">
              <RESULTS>
                <RESULT eventid="1088" points="377" swimtime="00:01:18.73" resultid="4311" heatid="5084" lane="1" entrytime="00:01:19.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="358" swimtime="00:10:36.28" resultid="4312" heatid="5298" lane="6" entrytime="00:10:40.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.14" />
                    <SPLIT distance="100" swimtime="00:01:14.40" />
                    <SPLIT distance="150" swimtime="00:01:54.75" />
                    <SPLIT distance="200" swimtime="00:02:35.21" />
                    <SPLIT distance="250" swimtime="00:03:15.82" />
                    <SPLIT distance="300" swimtime="00:03:56.37" />
                    <SPLIT distance="350" swimtime="00:04:36.68" />
                    <SPLIT distance="400" swimtime="00:05:17.39" />
                    <SPLIT distance="450" swimtime="00:05:58.39" />
                    <SPLIT distance="500" swimtime="00:06:39.80" />
                    <SPLIT distance="550" swimtime="00:07:20.83" />
                    <SPLIT distance="600" swimtime="00:08:02.08" />
                    <SPLIT distance="650" swimtime="00:08:42.67" />
                    <SPLIT distance="700" swimtime="00:09:23.01" />
                    <SPLIT distance="750" swimtime="00:10:00.52" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 9:58), Na volta dos 150m." eventid="1251" status="DSQ" swimtime="00:02:57.84" resultid="4313" heatid="5318" lane="1" entrytime="00:02:57.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.33" />
                    <SPLIT distance="100" swimtime="00:01:24.13" />
                    <SPLIT distance="150" swimtime="00:02:11.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="375" swimtime="00:00:35.98" resultid="4314" heatid="5368" lane="5" entrytime="00:00:35.79" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kedny" lastname="Correa" birthdate="2004-11-05" gender="M" nation="BRA" license="383858" swrid="5600142" athleteid="4327" externalid="383858">
              <RESULTS>
                <RESULT eventid="1072" points="459" swimtime="00:04:45.18" resultid="4328" heatid="5064" lane="2" entrytime="00:04:41.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="100" swimtime="00:01:06.06" />
                    <SPLIT distance="150" swimtime="00:01:41.91" />
                    <SPLIT distance="200" swimtime="00:02:18.42" />
                    <SPLIT distance="250" swimtime="00:02:55.37" />
                    <SPLIT distance="300" swimtime="00:03:33.05" />
                    <SPLIT distance="350" swimtime="00:04:10.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="439" swimtime="00:00:27.51" resultid="4329" heatid="5128" lane="1" entrytime="00:00:27.54" entrycourse="LCM" />
                <RESULT eventid="1120" points="426" swimtime="00:02:15.52" resultid="4330" heatid="5157" lane="4" entrytime="00:02:15.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                    <SPLIT distance="100" swimtime="00:01:05.47" />
                    <SPLIT distance="150" swimtime="00:01:40.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="366" swimtime="00:02:39.32" resultid="4331" heatid="5200" lane="2" entrytime="00:02:32.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.53" />
                    <SPLIT distance="100" swimtime="00:01:14.91" />
                    <SPLIT distance="150" swimtime="00:02:03.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1237" points="414" swimtime="00:04:12.56" resultid="4408" heatid="5308" lane="2" entrytime="00:04:16.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                    <SPLIT distance="100" swimtime="00:00:59.63" />
                    <SPLIT distance="150" swimtime="00:01:31.29" />
                    <SPLIT distance="200" swimtime="00:02:05.25" />
                    <SPLIT distance="250" swimtime="00:02:35.93" />
                    <SPLIT distance="300" swimtime="00:03:11.65" />
                    <SPLIT distance="350" swimtime="00:03:40.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4297" number="1" />
                    <RELAYPOSITION athleteid="4310" number="2" />
                    <RELAYPOSITION athleteid="4274" number="3" />
                    <RELAYPOSITION athleteid="4395" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1338" points="410" swimtime="00:04:38.21" resultid="4413" heatid="5388" lane="6" entrytime="00:04:55.56">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.63" />
                    <SPLIT distance="100" swimtime="00:01:08.41" />
                    <SPLIT distance="150" swimtime="00:01:45.63" />
                    <SPLIT distance="200" swimtime="00:02:26.84" />
                    <SPLIT distance="250" swimtime="00:03:00.28" />
                    <SPLIT distance="300" swimtime="00:03:37.18" />
                    <SPLIT distance="350" swimtime="00:04:06.34" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4297" number="1" />
                    <RELAYPOSITION athleteid="4310" number="2" />
                    <RELAYPOSITION athleteid="4254" number="3" />
                    <RELAYPOSITION athleteid="4395" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="19" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="M" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1239" points="525" swimtime="00:03:53.25" resultid="4409" heatid="5309" lane="4" entrytime="00:04:01.19">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                    <SPLIT distance="100" swimtime="00:00:57.55" />
                    <SPLIT distance="150" swimtime="00:01:27.19" />
                    <SPLIT distance="200" swimtime="00:02:00.08" />
                    <SPLIT distance="250" swimtime="00:02:27.39" />
                    <SPLIT distance="300" swimtime="00:02:58.05" />
                    <SPLIT distance="350" swimtime="00:03:24.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4364" number="1" />
                    <RELAYPOSITION athleteid="4290" number="2" />
                    <RELAYPOSITION athleteid="4248" number="3" />
                    <RELAYPOSITION athleteid="4322" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1340" points="423" swimtime="00:04:35.43" resultid="4411" heatid="5389" lane="4" entrytime="00:04:41.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                    <SPLIT distance="100" swimtime="00:01:11.26" />
                    <SPLIT distance="150" swimtime="00:01:49.24" />
                    <SPLIT distance="200" swimtime="00:02:37.19" />
                    <SPLIT distance="250" swimtime="00:03:06.57" />
                    <SPLIT distance="300" swimtime="00:03:40.79" />
                    <SPLIT distance="350" swimtime="00:04:06.87" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4364" number="1" />
                    <RELAYPOSITION athleteid="4402" number="2" />
                    <RELAYPOSITION athleteid="4248" number="3" />
                    <RELAYPOSITION athleteid="4322" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1233" points="351" swimtime="00:04:26.71" resultid="4410" heatid="5306" lane="7" entrytime="00:04:32.83">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.41" />
                    <SPLIT distance="100" swimtime="00:01:06.23" />
                    <SPLIT distance="150" swimtime="00:01:38.13" />
                    <SPLIT distance="200" swimtime="00:02:14.26" />
                    <SPLIT distance="250" swimtime="00:02:45.94" />
                    <SPLIT distance="300" swimtime="00:03:20.35" />
                    <SPLIT distance="350" swimtime="00:03:51.15" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4342" number="1" />
                    <RELAYPOSITION athleteid="4388" number="2" />
                    <RELAYPOSITION athleteid="4383" number="3" />
                    <RELAYPOSITION athleteid="4267" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1334" points="313" swimtime="00:05:04.43" resultid="4412" heatid="5386" lane="7" entrytime="00:05:28.10">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                    <SPLIT distance="100" swimtime="00:01:18.25" />
                    <SPLIT distance="150" swimtime="00:01:56.67" />
                    <SPLIT distance="200" swimtime="00:02:40.92" />
                    <SPLIT distance="250" swimtime="00:03:14.57" />
                    <SPLIT distance="300" swimtime="00:03:57.23" />
                    <SPLIT distance="350" swimtime="00:04:27.92" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4342" number="1" />
                    <RELAYPOSITION athleteid="4383" number="2" />
                    <RELAYPOSITION athleteid="4388" number="3" />
                    <RELAYPOSITION athleteid="4267" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1221" points="300" swimtime="00:05:10.61" resultid="4406" heatid="5302" lane="7" entrytime="00:05:15.43">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                    <SPLIT distance="100" swimtime="00:01:11.65" />
                    <SPLIT distance="150" swimtime="00:01:54.37" />
                    <SPLIT distance="200" swimtime="00:02:42.83" />
                    <SPLIT distance="250" swimtime="00:03:17.85" />
                    <SPLIT distance="300" swimtime="00:04:01.19" />
                    <SPLIT distance="350" swimtime="00:04:33.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4315" number="1" />
                    <RELAYPOSITION athleteid="4349" number="2" />
                    <RELAYPOSITION athleteid="4356" number="3" />
                    <RELAYPOSITION athleteid="4261" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1322" points="334" swimtime="00:05:31.99" resultid="4407" heatid="5382" lane="2" entrytime="00:05:55.27">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.95" />
                    <SPLIT distance="100" swimtime="00:01:37.66" />
                    <SPLIT distance="150" swimtime="00:02:14.92" />
                    <SPLIT distance="200" swimtime="00:02:58.19" />
                    <SPLIT distance="250" swimtime="00:03:32.83" />
                    <SPLIT distance="300" swimtime="00:04:22.44" />
                    <SPLIT distance="350" swimtime="00:04:55.65" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4349" number="1" />
                    <RELAYPOSITION athleteid="4261" number="2" />
                    <RELAYPOSITION athleteid="4356" number="3" />
                    <RELAYPOSITION athleteid="4315" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1287" points="370" swimtime="00:05:02.85" resultid="4414" heatid="5354" lane="6" entrytime="00:05:03.15">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.74" />
                    <SPLIT distance="100" swimtime="00:01:19.51" />
                    <SPLIT distance="150" swimtime="00:01:56.71" />
                    <SPLIT distance="200" swimtime="00:02:39.59" />
                    <SPLIT distance="250" swimtime="00:03:12.53" />
                    <SPLIT distance="300" swimtime="00:03:50.60" />
                    <SPLIT distance="350" swimtime="00:04:24.69" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4371" number="1" />
                    <RELAYPOSITION athleteid="4310" number="2" />
                    <RELAYPOSITION athleteid="4395" number="3" />
                    <RELAYPOSITION athleteid="4362" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="19" agemin="17" agetotalmax="-1" agetotalmin="-1" gender="X" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1289" points="399" swimtime="00:04:55.45" resultid="4415" heatid="5355" lane="4" entrytime="00:04:58.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.18" />
                    <SPLIT distance="100" swimtime="00:01:24.26" />
                    <SPLIT distance="150" swimtime="00:02:06.94" />
                    <SPLIT distance="200" swimtime="00:02:57.07" />
                    <SPLIT distance="250" swimtime="00:03:27.06" />
                    <SPLIT distance="300" swimtime="00:04:00.64" />
                    <SPLIT distance="350" swimtime="00:04:27.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4304" number="1" />
                    <RELAYPOSITION athleteid="4238" number="2" />
                    <RELAYPOSITION athleteid="4248" number="3" />
                    <RELAYPOSITION athleteid="4322" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="MORGENAU &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1283" points="317" swimtime="00:05:18.77" resultid="4416" heatid="5352" lane="1" entrytime="00:05:06.39">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.65" />
                    <SPLIT distance="100" swimtime="00:01:30.42" />
                    <SPLIT distance="150" swimtime="00:02:08.12" />
                    <SPLIT distance="200" swimtime="00:02:51.75" />
                    <SPLIT distance="250" swimtime="00:03:26.36" />
                    <SPLIT distance="300" swimtime="00:04:07.59" />
                    <SPLIT distance="350" swimtime="00:04:41.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="4267" number="1" />
                    <RELAYPOSITION athleteid="4261" number="2" />
                    <RELAYPOSITION athleteid="4388" number="3" />
                    <RELAYPOSITION athleteid="4315" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="13038" nation="BRA" region="PR" clubid="2693" swrid="93759" name="Associação De Pais E Atletas De Natação Ws/Crb" shortname="Apan/Ws">
          <ATHLETES>
            <ATHLETE firstname="Heloisa" lastname="Daniele Silva" birthdate="2010-07-06" gender="F" nation="BRA" license="359593" swrid="5588628" athleteid="2724" externalid="359593" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1096" points="517" swimtime="00:00:29.40" resultid="2725" heatid="5100" lane="5" entrytime="00:00:29.13" entrycourse="LCM" />
                <RESULT eventid="1175" points="394" swimtime="00:01:18.20" resultid="2726" heatid="5243" lane="4" entrytime="00:01:17.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="480" swimtime="00:01:06.02" resultid="2727" heatid="5205" lane="8" entrytime="00:01:06.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="469" swimtime="00:00:34.55" resultid="2728" heatid="5295" lane="8" entrytime="00:00:35.05" entrycourse="LCM" />
                <RESULT eventid="1259" points="338" swimtime="00:00:35.06" resultid="2729" heatid="5321" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="De Reginalda" birthdate="2011-07-22" gender="M" nation="BRA" license="400323" swrid="5717257" athleteid="2743" externalid="400323">
              <RESULTS>
                <RESULT eventid="1104" points="457" swimtime="00:00:27.14" resultid="2744" heatid="5119" lane="5" entrytime="00:00:27.61" entrycourse="LCM" />
                <RESULT eventid="1182" points="347" swimtime="00:01:13.36" resultid="2745" heatid="5257" lane="6" entrytime="00:01:12.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="428" swimtime="00:01:02.15" resultid="2746" heatid="5222" lane="1" entrytime="00:01:02.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="371" swimtime="00:00:32.77" resultid="2747" heatid="5285" lane="4" entrytime="00:00:32.96" entrycourse="LCM" />
                <RESULT eventid="1277" points="348" swimtime="00:02:39.07" resultid="2748" heatid="5345" lane="3" entrytime="00:02:40.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.65" />
                    <SPLIT distance="100" swimtime="00:01:16.57" />
                    <SPLIT distance="150" swimtime="00:01:58.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Marjori" lastname="Leticia Oliveira" birthdate="2011-05-23" gender="F" nation="BRA" license="406869" swrid="5717279" athleteid="2760" externalid="406869">
              <RESULTS>
                <RESULT eventid="1096" points="293" swimtime="00:00:35.54" resultid="2761" heatid="5097" lane="7" entrytime="00:00:35.29" entrycourse="LCM" />
                <RESULT eventid="1112" points="253" swimtime="00:02:58.20" resultid="2762" heatid="5138" lane="7" entrytime="00:02:57.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.71" />
                    <SPLIT distance="100" swimtime="00:01:25.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="251" swimtime="00:01:30.86" resultid="2763" heatid="5241" lane="5" entrytime="00:01:33.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="278" swimtime="00:01:19.21" resultid="2764" heatid="5201" lane="5" entrytime="00:01:20.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="256" swimtime="00:00:42.26" resultid="2765" heatid="5292" lane="1" entrytime="00:00:43.72" entrycourse="LCM" />
                <RESULT eventid="1259" points="157" swimtime="00:00:45.21" resultid="2766" heatid="5322" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luana" lastname="Zeclhynski Silva" birthdate="2006-09-14" gender="F" nation="BRA" license="330727" swrid="5600283" athleteid="2694" externalid="330727" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1096" points="630" swimtime="00:00:27.54" resultid="2695" heatid="5106" lane="4" entrytime="00:00:27.78" entrycourse="LCM" />
                <RESULT eventid="1143" points="475" swimtime="00:02:41.58" resultid="2696" heatid="5191" lane="5" entrytime="00:02:42.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                    <SPLIT distance="100" swimtime="00:01:10.08" />
                    <SPLIT distance="150" swimtime="00:02:04.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="560" swimtime="00:01:09.55" resultid="2697" heatid="5248" lane="4" entrytime="00:01:06.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="638" swimtime="00:01:00.04" resultid="2698" heatid="5209" lane="3" entrytime="00:01:00.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="602" swimtime="00:00:31.81" resultid="2699" heatid="5295" lane="4" entrytime="00:00:30.32" entrycourse="LCM" />
                <RESULT eventid="2375" points="625" swimtime="00:00:27.60" resultid="5969" heatid="5978" lane="5" entrytime="00:00:27.54" />
                <RESULT eventid="2343" points="632" swimtime="00:01:00.24" resultid="6101" heatid="6421" lane="4" entrytime="00:01:00.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2391" points="603" swimtime="00:01:07.85" resultid="6129" heatid="6424" lane="3" entrytime="00:01:09.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Da Costa Riekes" birthdate="2008-06-19" gender="F" nation="BRA" license="331686" swrid="5600143" athleteid="2706" externalid="331686" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1096" points="549" swimtime="00:00:28.82" resultid="2707" heatid="5104" lane="7" entrytime="00:00:29.28" entrycourse="LCM" />
                <RESULT eventid="1128" points="394" swimtime="00:01:15.66" resultid="2708" heatid="5161" lane="3" entrytime="00:01:13.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="499" swimtime="00:02:22.27" resultid="2709" heatid="5144" lane="6" entrytime="00:02:20.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.73" />
                    <SPLIT distance="100" swimtime="00:01:08.27" />
                    <SPLIT distance="150" swimtime="00:01:45.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="435" swimtime="00:01:15.62" resultid="2710" heatid="5247" lane="7" entrytime="00:01:13.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="541" swimtime="00:01:03.46" resultid="2711" heatid="5208" lane="7" entrytime="00:01:03.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2375" points="560" swimtime="00:00:28.63" resultid="5974" heatid="5978" lane="7" entrytime="00:00:28.82" />
                <RESULT eventid="2328" swimtime="00:00:00.00" resultid="6006" entrytime="00:01:15.66" />
                <RESULT eventid="2343" swimtime="00:00:00.00" resultid="6109" entrytime="00:01:03.46" />
                <RESULT eventid="2391" points="421" swimtime="00:01:16.48" resultid="6136" entrytime="00:01:15.62">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Fernandes Ferreira" birthdate="2008-07-28" gender="M" nation="BRA" license="414578" swrid="5755373" athleteid="2767" externalid="414578">
              <RESULTS>
                <RESULT eventid="1104" points="405" swimtime="00:00:28.26" resultid="2768" heatid="5122" lane="4" entrytime="00:00:28.45" entrycourse="LCM" />
                <RESULT eventid="1167" points="407" swimtime="00:01:03.20" resultid="2769" heatid="5225" lane="5" entrytime="00:01:04.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="384" swimtime="00:00:32.39" resultid="2770" heatid="5283" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Sieck" birthdate="2011-01-20" gender="F" nation="BRA" license="382234" swrid="5602584" athleteid="2737" externalid="382234">
              <RESULTS>
                <RESULT eventid="1096" points="302" swimtime="00:00:35.18" resultid="2738" heatid="5096" lane="3" entrytime="00:00:37.15" entrycourse="LCM" />
                <RESULT eventid="1128" points="185" swimtime="00:01:37.33" resultid="2739" heatid="5159" lane="2" entrytime="00:01:45.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="205" swimtime="00:00:45.50" resultid="2740" heatid="5289" lane="5" />
                <RESULT eventid="1259" points="206" swimtime="00:00:41.33" resultid="2741" heatid="5323" lane="2" entrytime="00:00:42.22" entrycourse="LCM" />
                <RESULT eventid="1295" points="162" swimtime="00:03:43.32" resultid="2742" heatid="5361" lane="5" entrytime="00:04:14.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.73" />
                    <SPLIT distance="100" swimtime="00:01:40.96" />
                    <SPLIT distance="150" swimtime="00:02:44.37" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Rosa Silva" birthdate="2011-03-25" gender="F" nation="BRA" license="392120" swrid="5602579" athleteid="2718" externalid="392120">
              <RESULTS>
                <RESULT eventid="1080" points="228" swimtime="00:01:44.97" resultid="2719" heatid="5065" lane="3" entrytime="00:01:47.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="265" swimtime="00:00:36.75" resultid="2720" heatid="5096" lane="4" entrytime="00:00:36.86" entrycourse="LCM" />
                <RESULT eventid="1143" points="225" swimtime="00:03:27.23" resultid="2721" heatid="5186" lane="6" entrytime="00:03:36.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.94" />
                    <SPLIT distance="100" swimtime="00:01:38.97" />
                    <SPLIT distance="150" swimtime="00:02:42.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="240" swimtime="00:01:23.14" resultid="2722" heatid="5201" lane="6" entrytime="00:01:21.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="229" swimtime="00:00:47.62" resultid="2723" heatid="5373" lane="4" entrytime="00:00:51.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Zanchetta Silva" birthdate="2010-08-05" gender="F" nation="BRA" license="406865" swrid="5717308" athleteid="2749" externalid="406865">
              <RESULTS>
                <RESULT eventid="1096" points="252" swimtime="00:00:37.34" resultid="2750" heatid="5096" lane="5" entrytime="00:00:37.13" entrycourse="LCM" />
                <RESULT eventid="1175" points="154" swimtime="00:01:46.88" resultid="2751" heatid="5241" lane="6" entrytime="00:01:41.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="240" swimtime="00:01:23.20" resultid="2752" heatid="5201" lane="3" entrytime="00:01:21.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="197" swimtime="00:00:46.10" resultid="2753" heatid="5291" lane="6" entrytime="00:00:46.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniel" lastname="Cravcenco Marcondes" birthdate="2011-05-06" gender="M" nation="BRA" license="406867" swrid="5723023" athleteid="2754" externalid="406867">
              <RESULTS>
                <RESULT eventid="1104" points="286" swimtime="00:00:31.73" resultid="2755" heatid="5116" lane="5" entrytime="00:00:31.31" entrycourse="LCM" />
                <RESULT eventid="1167" points="290" swimtime="00:01:10.73" resultid="2756" heatid="5219" lane="6" entrytime="00:01:12.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="230" swimtime="00:00:38.42" resultid="2757" heatid="5284" lane="7" entrytime="00:00:42.45" entrycourse="LCM" />
                <RESULT eventid="1267" points="237" swimtime="00:00:35.94" resultid="2758" heatid="5331" lane="1" entrytime="00:00:36.93" entrycourse="LCM" />
                <RESULT eventid="1297" points="181" swimtime="00:00:45.81" resultid="2759" heatid="5366" lane="1" entrytime="00:00:49.09" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Reis" birthdate="2008-04-07" gender="F" nation="BRA" license="378820" swrid="5600243" athleteid="2730" externalid="378820" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1096" points="308" swimtime="00:00:34.93" resultid="2731" heatid="5102" lane="8" entrytime="00:00:35.56" entrycourse="LCM" />
                <RESULT eventid="1128" points="187" swimtime="00:01:36.96" resultid="2732" heatid="5161" lane="7" entrytime="00:01:44.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="250" swimtime="00:01:30.99" resultid="2733" heatid="5245" lane="5" entrytime="00:01:30.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="268" swimtime="00:01:20.14" resultid="2734" heatid="5206" lane="3" entrytime="00:01:21.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="260" swimtime="00:00:42.05" resultid="2735" heatid="5292" lane="8" entrytime="00:00:43.74" entrycourse="LCM" />
                <RESULT eventid="1259" points="190" swimtime="00:00:42.43" resultid="2736" heatid="5323" lane="7" entrytime="00:00:42.86" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonia" lastname="Adam  Fracaro" birthdate="2010-04-27" gender="F" nation="BRA" license="382212" swrid="5588512" athleteid="2700" externalid="382212">
              <RESULTS>
                <RESULT eventid="1080" points="149" swimtime="00:02:00.76" resultid="2701" heatid="5065" lane="2" entrytime="00:01:58.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" points="311" swimtime="00:05:47.36" resultid="2702" heatid="5049" lane="8" entrytime="00:05:59.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="100" swimtime="00:01:19.44" />
                    <SPLIT distance="150" swimtime="00:02:03.03" />
                    <SPLIT distance="200" swimtime="00:02:48.10" />
                    <SPLIT distance="250" swimtime="00:03:32.54" />
                    <SPLIT distance="300" swimtime="00:04:18.75" />
                    <SPLIT distance="350" swimtime="00:05:04.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="300" swimtime="00:02:48.39" resultid="2703" heatid="5138" lane="3" entrytime="00:02:43.66" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                    <SPLIT distance="100" swimtime="00:01:21.51" />
                    <SPLIT distance="150" swimtime="00:02:06.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="313" swimtime="00:01:16.13" resultid="2704" heatid="5202" lane="5" entrytime="00:01:13.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="180" swimtime="00:00:51.62" resultid="2705" heatid="5373" lane="5" entrytime="00:00:52.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabelly" lastname="Mendonca Bello" birthdate="2008-04-15" gender="F" nation="BRA" license="376996" swrid="5600217" athleteid="2712" externalid="376996" level="SMELJ CURI">
              <RESULTS>
                <RESULT eventid="1080" points="400" swimtime="00:01:26.98" resultid="2713" heatid="5068" lane="5" entrytime="00:01:24.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="463" swimtime="00:00:30.50" resultid="2714" heatid="5103" lane="6" entrytime="00:00:30.10" entrycourse="LCM" />
                <RESULT eventid="1143" points="377" swimtime="00:02:54.44" resultid="2715" heatid="5189" lane="3" entrytime="00:02:51.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.85" />
                    <SPLIT distance="100" swimtime="00:01:25.65" />
                    <SPLIT distance="150" swimtime="00:02:17.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="379" swimtime="00:03:09.91" resultid="2716" heatid="5312" lane="7" entrytime="00:03:11.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.35" />
                    <SPLIT distance="100" swimtime="00:01:31.23" />
                    <SPLIT distance="150" swimtime="00:02:21.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="387" swimtime="00:00:40.00" resultid="2717" heatid="5376" lane="6" entrytime="00:00:38.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2864" nation="BRA" region="PR" clubid="2441" swrid="93756" name="Associacao De Pais E Amigos Da Natacao De Ponta Gr" shortname="Apan Ponta Grossa">
          <ATHLETES>
            <ATHLETE firstname="Felipe" lastname="Chi Kravchychyn" birthdate="2009-09-27" gender="M" nation="BRA" license="344268" swrid="5600134" athleteid="2448" externalid="344268">
              <RESULTS>
                <RESULT eventid="1088" points="524" swimtime="00:01:10.51" resultid="2449" heatid="5085" lane="5" entrytime="00:01:09.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="524" swimtime="00:01:01.32" resultid="2450" heatid="5175" lane="1" entrytime="00:01:01.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="532" swimtime="00:02:20.66" resultid="2451" heatid="5198" lane="6" entrytime="00:02:17.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.06" />
                    <SPLIT distance="100" swimtime="00:01:06.71" />
                    <SPLIT distance="150" swimtime="00:01:47.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="493" swimtime="00:05:06.81" resultid="2452" heatid="5277" lane="3" entrytime="00:04:51.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.14" />
                    <SPLIT distance="100" swimtime="00:01:07.08" />
                    <SPLIT distance="150" swimtime="00:01:47.93" />
                    <SPLIT distance="200" swimtime="00:02:28.23" />
                    <SPLIT distance="250" swimtime="00:03:12.76" />
                    <SPLIT distance="300" swimtime="00:03:55.03" />
                    <SPLIT distance="350" swimtime="00:04:31.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="521" swimtime="00:02:35.94" resultid="2453" heatid="5320" lane="2" entrytime="00:02:30.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.78" />
                    <SPLIT distance="100" swimtime="00:01:14.56" />
                    <SPLIT distance="150" swimtime="00:01:55.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1293" status="DNS" swimtime="00:00:00.00" resultid="2454" heatid="5360" lane="2" entrytime="00:02:16.82" entrycourse="LCM" />
                <RESULT eventid="2320" swimtime="00:00:00.00" resultid="5962" entrytime="00:01:10.51" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yohan" lastname="Rigoni Moraes" birthdate="2002-04-03" gender="M" nation="BRA" license="272187" swrid="5600245" athleteid="2455" externalid="272187" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1088" points="606" swimtime="00:01:07.21" resultid="2456" heatid="5087" lane="3" entrytime="00:01:06.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="713" swimtime="00:00:29.04" resultid="2457" heatid="5371" lane="4" entrytime="00:00:28.71" entrycourse="LCM" />
                <RESULT eventid="2320" points="619" swimtime="00:01:06.74" resultid="5954" heatid="6414" lane="5" entrytime="00:01:07.21">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Lievore" birthdate="2010-06-07" gender="F" nation="BRA" license="414856" athleteid="2516" externalid="414856">
              <RESULTS>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 11:50)" eventid="1096" status="DSQ" swimtime="00:00:32.76" resultid="2517" heatid="5095" lane="5" />
                <RESULT eventid="1159" points="327" swimtime="00:01:15.00" resultid="2518" heatid="5201" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Carraro Borges" birthdate="2009-05-11" gender="M" nation="BRA" license="345590" swrid="5622267" athleteid="2487" externalid="345590" level="SAGRADA FA">
              <RESULTS>
                <RESULT eventid="1072" points="385" swimtime="00:05:02.36" resultid="2488" heatid="5061" lane="6" entrytime="00:04:47.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                    <SPLIT distance="100" swimtime="00:01:08.51" />
                    <SPLIT distance="150" swimtime="00:01:46.05" />
                    <SPLIT distance="200" swimtime="00:02:25.50" />
                    <SPLIT distance="250" swimtime="00:03:06.37" />
                    <SPLIT distance="300" swimtime="00:03:45.11" />
                    <SPLIT distance="350" swimtime="00:04:24.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="413" swimtime="00:02:16.94" resultid="2489" heatid="5155" lane="8" entrytime="00:02:15.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                    <SPLIT distance="100" swimtime="00:01:04.80" />
                    <SPLIT distance="150" swimtime="00:01:40.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="438" swimtime="00:01:01.68" resultid="2490" heatid="5227" lane="8" entrytime="00:01:01.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="354" swimtime="00:10:39.11" resultid="2491" heatid="5299" lane="6" entrytime="00:10:01.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                    <SPLIT distance="100" swimtime="00:01:09.79" />
                    <SPLIT distance="150" swimtime="00:01:47.50" />
                    <SPLIT distance="200" swimtime="00:02:26.64" />
                    <SPLIT distance="250" swimtime="00:03:06.44" />
                    <SPLIT distance="300" swimtime="00:03:45.92" />
                    <SPLIT distance="400" swimtime="00:05:08.08" />
                    <SPLIT distance="450" swimtime="00:05:49.67" />
                    <SPLIT distance="500" swimtime="00:06:31.45" />
                    <SPLIT distance="600" swimtime="00:07:55.28" />
                    <SPLIT distance="650" swimtime="00:08:37.08" />
                    <SPLIT distance="700" swimtime="00:09:18.46" />
                    <SPLIT distance="750" swimtime="00:09:59.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" status="DNS" swimtime="00:00:00.00" resultid="2492" heatid="5380" lane="1" entrytime="00:19:19.25" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Carolina Babiuki" birthdate="2007-02-06" gender="F" nation="BRA" license="316227" swrid="5600131" athleteid="2472" externalid="316227" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1096" points="553" swimtime="00:00:28.75" resultid="2473" heatid="5106" lane="5" entrytime="00:00:28.74" entrycourse="LCM" />
                <RESULT eventid="1175" points="502" swimtime="00:01:12.11" resultid="2474" heatid="5248" lane="3" entrytime="00:01:12.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="570" swimtime="00:00:32.39" resultid="2475" heatid="5295" lane="6" entrytime="00:00:32.70" entrycourse="LCM" />
                <RESULT eventid="2375" points="539" swimtime="00:00:29.01" resultid="5973" heatid="5978" lane="2" entrytime="00:00:28.75" />
                <RESULT eventid="2391" points="498" swimtime="00:01:12.31" resultid="6132" heatid="6424" lane="2" entrytime="00:01:12.11">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Allana" lastname="Lacerda" birthdate="2005-03-15" gender="F" nation="BRA" license="295186" swrid="5600197" athleteid="2458" externalid="295186" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1080" points="432" swimtime="00:01:24.80" resultid="2459" heatid="5070" lane="3" entrytime="00:01:22.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="418" swimtime="00:02:30.91" resultid="2460" heatid="5146" lane="7" entrytime="00:02:30.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.56" />
                    <SPLIT distance="100" swimtime="00:01:13.64" />
                    <SPLIT distance="150" swimtime="00:01:53.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="424" swimtime="00:03:03.04" resultid="2461" heatid="5313" lane="6" entrytime="00:02:58.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                    <SPLIT distance="100" swimtime="00:01:28.93" />
                    <SPLIT distance="150" swimtime="00:02:16.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="423" swimtime="00:00:38.84" resultid="2462" heatid="5376" lane="2" entrytime="00:00:38.77" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Brenda" lastname="Gabriele Carvalho" birthdate="2010-04-11" gender="F" nation="BRA" license="399557" swrid="5658060" athleteid="2496" externalid="399557">
              <RESULTS>
                <RESULT eventid="1175" points="272" swimtime="00:01:28.44" resultid="2497" heatid="5242" lane="8" entrytime="00:01:29.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="311" swimtime="00:01:16.26" resultid="2498" heatid="5202" lane="7" entrytime="00:01:18.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="291" swimtime="00:00:40.51" resultid="2499" heatid="5292" lane="4" entrytime="00:00:40.96" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Fegert" birthdate="2009-04-13" gender="M" nation="BRA" license="353813" swrid="5622279" athleteid="2482" externalid="353813">
              <RESULTS>
                <RESULT eventid="1104" points="489" swimtime="00:00:26.53" resultid="2483" heatid="5124" lane="4" entrytime="00:00:26.58" entrycourse="LCM" />
                <RESULT eventid="1135" points="430" swimtime="00:01:05.47" resultid="2484" heatid="5174" lane="1" entrytime="00:01:05.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="488" swimtime="00:00:59.50" resultid="2485" heatid="5228" lane="1" entrytime="00:00:59.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="495" swimtime="00:00:28.15" resultid="2486" heatid="5334" lane="2" entrytime="00:00:29.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Augusto" lastname="Tramontin" birthdate="2011-11-29" gender="M" nation="BRA" license="399691" swrid="5652901" athleteid="2500" externalid="399691">
              <RESULTS>
                <RESULT eventid="1088" points="302" swimtime="00:01:24.76" resultid="2501" heatid="5082" lane="8" entrytime="00:01:23.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="383" swimtime="00:00:28.78" resultid="2502" heatid="5118" lane="4" entrytime="00:00:28.73" entrycourse="LCM" />
                <RESULT eventid="1167" points="389" swimtime="00:01:04.15" resultid="2503" heatid="5221" lane="5" entrytime="00:01:04.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="374" swimtime="00:00:35.99" resultid="2504" heatid="5367" lane="5" entrytime="00:00:38.38" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Delinski" birthdate="2009-11-28" gender="F" nation="BRA" license="385190" swrid="5600150" athleteid="2476" externalid="385190">
              <RESULTS>
                <RESULT eventid="1080" points="388" swimtime="00:01:27.92" resultid="2477" heatid="5068" lane="3" entrytime="00:01:28.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="327" swimtime="00:01:23.13" resultid="2478" heatid="5246" lane="6" entrytime="00:01:21.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="367" swimtime="00:00:37.51" resultid="2479" heatid="5293" lane="5" entrytime="00:00:37.58" entrycourse="LCM" />
                <RESULT eventid="1243" points="288" swimtime="00:03:28.15" resultid="2480" heatid="5311" lane="6" entrytime="00:03:21.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.70" />
                    <SPLIT distance="100" swimtime="00:01:41.41" />
                    <SPLIT distance="150" swimtime="00:02:38.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="384" swimtime="00:00:40.10" resultid="2481" heatid="5375" lane="2" entrytime="00:00:42.30" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Franca Berger" birthdate="2010-05-07" gender="F" nation="BRA" license="399692" swrid="5653290" athleteid="2505" externalid="399692">
              <RESULTS>
                <RESULT eventid="1096" points="323" swimtime="00:00:34.39" resultid="2506" heatid="5097" lane="2" entrytime="00:00:35.17" entrycourse="LCM" />
                <RESULT eventid="1159" points="296" swimtime="00:01:17.55" resultid="2507" heatid="5202" lane="8" entrytime="00:01:19.05" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="136" swimtime="00:00:47.50" resultid="2508" heatid="5323" lane="1" entrytime="00:00:44.81" entrycourse="LCM" />
                <RESULT eventid="1305" points="273" swimtime="00:00:44.90" resultid="2509" heatid="5374" lane="7" entrytime="00:00:47.88" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carolina" lastname="Reda" birthdate="2007-05-21" gender="F" nation="BRA" license="316228" swrid="5600241" athleteid="2468" externalid="316228">
              <RESULTS>
                <RESULT eventid="1096" points="384" swimtime="00:00:32.46" resultid="2469" heatid="5106" lane="7" entrytime="00:00:32.08" entrycourse="LCM" />
                <RESULT eventid="1159" points="381" swimtime="00:01:11.29" resultid="2470" heatid="5209" lane="7" entrytime="00:01:11.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="369" swimtime="00:00:37.43" resultid="2471" heatid="5294" lane="1" entrytime="00:00:36.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Gueiber Montes" birthdate="2009-03-09" gender="M" nation="BRA" license="342154" swrid="5600179" athleteid="2442" externalid="342154">
              <RESULTS>
                <RESULT eventid="1104" points="583" swimtime="00:00:25.03" resultid="2443" heatid="5126" lane="5" entrytime="00:00:24.54" entrycourse="LCM" />
                <RESULT eventid="1120" points="593" swimtime="00:02:01.40" resultid="2444" heatid="5156" lane="4" entrytime="00:02:00.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.66" />
                    <SPLIT distance="100" swimtime="00:00:57.95" />
                    <SPLIT distance="150" swimtime="00:01:30.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="646" swimtime="00:00:54.20" resultid="2445" heatid="5230" lane="3" entrytime="00:00:54.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="550" swimtime="00:00:28.73" resultid="2446" heatid="5288" lane="8" entrytime="00:00:28.83" entrycourse="LCM" />
                <RESULT eventid="1267" points="553" swimtime="00:00:27.13" resultid="2447" heatid="5329" lane="1" />
                <RESULT eventid="2351" swimtime="00:00:00.00" resultid="6125" entrytime="00:00:54.20" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Sabedotti" birthdate="2011-04-20" gender="F" nation="BRA" license="390877" swrid="5602580" athleteid="2512" externalid="390877">
              <RESULTS>
                <RESULT eventid="1175" points="402" swimtime="00:01:17.65" resultid="2513" heatid="5243" lane="6" entrytime="00:01:18.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="434" swimtime="00:00:35.46" resultid="2514" heatid="5295" lane="1" entrytime="00:00:34.92" entrycourse="LCM" />
                <RESULT eventid="1259" points="399" swimtime="00:00:33.16" resultid="2515" heatid="5321" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Pontes Mattioli" birthdate="2011-09-10" gender="F" nation="BRA" license="366914" swrid="5602572" athleteid="2510" externalid="366914">
              <RESULTS>
                <RESULT eventid="1259" points="341" swimtime="00:00:34.96" resultid="2511" heatid="5324" lane="3" entrytime="00:00:35.82" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yoseph" lastname="Rigoni Moraes" birthdate="2006-04-17" gender="M" nation="BRA" license="295182" swrid="5622302" athleteid="2493" externalid="295182" level="POSITIVO M">
              <RESULTS>
                <RESULT eventid="1267" points="522" swimtime="00:00:27.65" resultid="2494" heatid="5336" lane="4" entrytime="00:00:27.50" entrycourse="LCM" />
                <RESULT eventid="1297" points="471" swimtime="00:00:33.33" resultid="2495" heatid="5370" lane="3" entrytime="00:00:32.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Barbara" lastname="Campagnoli" birthdate="2009-04-13" gender="F" nation="BRA" license="366915" swrid="5600128" athleteid="2463" externalid="366915">
              <RESULTS>
                <RESULT eventid="1096" points="536" swimtime="00:00:29.05" resultid="2464" heatid="5104" lane="2" entrytime="00:00:29.10" entrycourse="LCM" />
                <RESULT eventid="1112" points="500" swimtime="00:02:22.09" resultid="2465" heatid="5144" lane="3" entrytime="00:02:19.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.93" />
                    <SPLIT distance="100" swimtime="00:01:08.11" />
                    <SPLIT distance="150" swimtime="00:01:45.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="521" swimtime="00:01:11.22" resultid="2466" heatid="5247" lane="6" entrytime="00:01:11.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="515" swimtime="00:00:33.49" resultid="2467" heatid="5295" lane="7" entrytime="00:00:33.45" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/PONTA GROSSA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1235" points="516" swimtime="00:03:54.66" resultid="2520" heatid="5307" lane="5" entrytime="00:03:54.97">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.13" />
                    <SPLIT distance="100" swimtime="00:01:00.14" />
                    <SPLIT distance="150" swimtime="00:01:26.78" />
                    <SPLIT distance="200" swimtime="00:01:57.85" />
                    <SPLIT distance="250" swimtime="00:02:26.88" />
                    <SPLIT distance="300" swimtime="00:02:59.47" />
                    <SPLIT distance="350" swimtime="00:03:25.67" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2482" number="1" />
                    <RELAYPOSITION athleteid="2448" number="2" />
                    <RELAYPOSITION athleteid="2487" number="3" />
                    <RELAYPOSITION athleteid="2442" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1336" status="WDR" swimtime="00:00:00.00" resultid="2521" heatid="5387" lane="5" entrytime="00:04:23.71" />
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="APAN/PONTA GROSSA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1221" points="352" swimtime="00:04:54.28" resultid="2519" heatid="5302" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.52" />
                    <SPLIT distance="100" swimtime="00:01:06.59" />
                    <SPLIT distance="150" swimtime="00:01:41.46" />
                    <SPLIT distance="200" swimtime="00:02:22.74" />
                    <SPLIT distance="250" swimtime="00:02:55.62" />
                    <SPLIT distance="300" swimtime="00:03:34.94" />
                    <SPLIT distance="350" swimtime="00:04:11.79" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2512" number="1" />
                    <RELAYPOSITION athleteid="2505" number="2" />
                    <RELAYPOSITION athleteid="2516" number="3" />
                    <RELAYPOSITION athleteid="2496" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="20" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/PONTA GROSSA &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1291" points="430" swimtime="00:04:48.18" resultid="2522" heatid="5356" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.24" />
                    <SPLIT distance="100" swimtime="00:01:15.89" />
                    <SPLIT distance="150" swimtime="00:01:49.79" />
                    <SPLIT distance="200" swimtime="00:02:25.88" />
                    <SPLIT distance="250" swimtime="00:02:57.24" />
                    <SPLIT distance="300" swimtime="00:03:36.46" />
                    <SPLIT distance="350" swimtime="00:04:10.29" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2472" number="1" />
                    <RELAYPOSITION athleteid="2455" number="2" />
                    <RELAYPOSITION athleteid="2493" number="3" />
                    <RELAYPOSITION athleteid="2458" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="2416" nation="BRA" region="PR" clubid="2523" swrid="93758" name="Apan/Maringá">
          <ATHLETES>
            <ATHLETE firstname="Gabriel" lastname="Casavechia Carraro" birthdate="2009-07-28" gender="M" nation="BRA" license="368150" swrid="5384752" athleteid="2524" externalid="368150">
              <RESULTS>
                <RESULT eventid="1104" points="585" swimtime="00:00:25.00" resultid="2525" heatid="5126" lane="2" entrytime="00:00:24.82" entrycourse="LCM" />
                <RESULT eventid="1135" points="584" swimtime="00:00:59.14" resultid="2526" heatid="5175" lane="5" entrytime="00:00:58.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="682" swimtime="00:00:53.23" resultid="2527" heatid="5230" lane="4" entrytime="00:00:53.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="569" swimtime="00:00:26.87" resultid="2528" heatid="5337" lane="3" entrytime="00:00:27.02" entrycourse="LCM" />
                <RESULT eventid="1293" points="390" swimtime="00:02:30.95" resultid="2529" heatid="5357" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.60" />
                    <SPLIT distance="100" swimtime="00:01:08.23" />
                    <SPLIT distance="150" swimtime="00:01:49.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2335" swimtime="00:00:00.00" resultid="6016" entrytime="00:00:59.14" />
                <RESULT eventid="2351" points="667" swimtime="00:00:53.61" resultid="6119" heatid="6422" lane="6" entrytime="00:00:53.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Sol Reolon Gomes" birthdate="2011-02-28" gender="F" nation="BRA" license="392100" swrid="5603914" athleteid="2656" externalid="392100">
              <RESULTS>
                <RESULT eventid="1096" points="503" swimtime="00:00:29.67" resultid="2657" heatid="5100" lane="2" entrytime="00:00:29.73" entrycourse="LCM" />
                <RESULT eventid="1112" points="411" swimtime="00:02:31.74" resultid="2658" heatid="5139" lane="6" entrytime="00:02:33.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:12.26" />
                    <SPLIT distance="150" swimtime="00:01:53.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="409" swimtime="00:01:17.18" resultid="2659" heatid="5244" lane="6" entrytime="00:01:15.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="488" swimtime="00:00:34.11" resultid="2660" heatid="5294" lane="8" entrytime="00:00:36.89" entrycourse="LCM" />
                <RESULT eventid="1259" points="407" swimtime="00:00:32.96" resultid="2661" heatid="5324" lane="4" entrytime="00:00:35.74" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Passafaro" birthdate="2009-02-01" gender="F" nation="BRA" license="370673" swrid="5603885" athleteid="2595" externalid="370673">
              <RESULTS>
                <RESULT eventid="1096" points="391" swimtime="00:00:32.28" resultid="2596" heatid="5103" lane="7" entrytime="00:00:30.34" entrycourse="LCM" />
                <RESULT eventid="1128" points="232" swimtime="00:01:30.20" resultid="2597" heatid="5161" lane="2" entrytime="00:01:29.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" status="DNS" swimtime="00:00:00.00" resultid="2598" heatid="5206" lane="5" entrytime="00:01:10.85" entrycourse="LCM" />
                <RESULT eventid="1259" points="358" swimtime="00:00:34.38" resultid="2599" heatid="5325" lane="5" entrytime="00:00:34.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Garcia Cavalcante" birthdate="2011-11-21" gender="M" nation="BRA" license="378200" swrid="5603840" athleteid="2555" externalid="378200">
              <RESULTS>
                <RESULT eventid="1088" points="281" swimtime="00:01:26.75" resultid="2556" heatid="5081" lane="6" entrytime="00:01:27.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="289" swimtime="00:02:34.25" resultid="2557" heatid="5147" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.75" />
                    <SPLIT distance="100" swimtime="00:01:13.50" />
                    <SPLIT distance="150" swimtime="00:01:54.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="323" swimtime="00:01:08.23" resultid="2558" heatid="5218" lane="4" entrytime="00:01:17.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="287" swimtime="00:03:10.10" resultid="2559" heatid="5317" lane="8" entrytime="00:03:13.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.74" />
                    <SPLIT distance="100" swimtime="00:01:35.54" />
                    <SPLIT distance="150" swimtime="00:02:24.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="286" swimtime="00:00:39.38" resultid="2560" heatid="5367" lane="2" entrytime="00:00:40.56" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Corsine Ferreira" birthdate="2010-03-10" gender="F" nation="BRA" license="353591" swrid="5588608" athleteid="2636" externalid="353591">
              <RESULTS>
                <RESULT eventid="1080" points="357" swimtime="00:01:30.38" resultid="2637" heatid="5065" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="353" swimtime="00:02:39.53" resultid="2638" heatid="5139" lane="8" entrytime="00:02:39.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.30" />
                    <SPLIT distance="100" swimtime="00:01:15.46" />
                    <SPLIT distance="150" swimtime="00:01:57.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="387" swimtime="00:01:18.61" resultid="2639" heatid="5244" lane="8" entrytime="00:01:16.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="436" swimtime="00:00:35.40" resultid="2640" heatid="5294" lane="4" entrytime="00:00:35.38" entrycourse="LCM" />
                <RESULT eventid="1275" points="374" swimtime="00:02:50.80" resultid="2641" heatid="5342" lane="6" entrytime="00:02:46.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:23.76" />
                    <SPLIT distance="150" swimtime="00:02:07.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="368" swimtime="00:00:40.69" resultid="2642" heatid="5375" lane="5" entrytime="00:00:40.21" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Antônio Boeing" birthdate="2004-06-04" gender="M" nation="BRA" license="317474" swrid="5184340" athleteid="2561" externalid="317474">
              <RESULTS>
                <RESULT eventid="1088" points="581" swimtime="00:01:08.13" resultid="2562" heatid="5086" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="667" swimtime="00:00:23.93" resultid="2563" heatid="5130" lane="2" entrytime="00:00:23.96" entrycourse="LCM" />
                <RESULT eventid="1135" points="691" swimtime="00:00:55.92" resultid="2564" heatid="5178" lane="4" entrytime="00:00:54.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="678" swimtime="00:00:26.80" resultid="2565" heatid="5288" lane="5" entrytime="00:00:26.92" entrycourse="LCM" />
                <RESULT eventid="1267" points="727" swimtime="00:00:24.76" resultid="2566" heatid="5338" lane="4" entrytime="00:00:24.81" entrycourse="LCM" />
                <RESULT eventid="1297" points="650" swimtime="00:00:29.95" resultid="2567" heatid="5364" lane="3" />
                <RESULT eventid="2320" points="597" swimtime="00:01:07.54" resultid="5957" heatid="6414" lane="2" entrytime="00:01:08.13">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2383" points="693" swimtime="00:00:23.62" resultid="5981" heatid="6425" lane="3" entrytime="00:00:23.93" />
                <RESULT eventid="2335" points="691" swimtime="00:00:55.92" resultid="6009" heatid="6417" lane="5" entrytime="00:00:55.92">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Furuchi Martins" birthdate="2011-10-05" gender="F" nation="BRA" license="367001" swrid="5602616" athleteid="2668" externalid="367001">
              <RESULTS>
                <RESULT eventid="1080" points="317" swimtime="00:01:34.02" resultid="2669" heatid="5066" lane="1" entrytime="00:01:32.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="277" swimtime="00:03:13.28" resultid="2670" heatid="5186" lane="4" entrytime="00:03:17.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:39.23" />
                    <SPLIT distance="150" swimtime="00:02:31.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="265" swimtime="00:00:41.80" resultid="2671" heatid="5291" lane="7" entrytime="00:00:48.15" entrycourse="LCM" />
                <RESULT eventid="1243" points="293" swimtime="00:03:26.87" resultid="2672" heatid="5311" lane="7" entrytime="00:03:26.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.49" />
                    <SPLIT distance="100" swimtime="00:01:40.79" />
                    <SPLIT distance="150" swimtime="00:02:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="335" swimtime="00:00:41.97" resultid="2673" heatid="5374" lane="5" entrytime="00:00:43.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanni" lastname="Lazzari Mariotti" birthdate="2006-08-14" gender="M" nation="BRA" license="341929" swrid="5615873" athleteid="2572" externalid="341929">
              <RESULTS>
                <RESULT eventid="1088" points="556" swimtime="00:01:09.17" resultid="2573" heatid="5087" lane="6" entrytime="00:01:07.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" status="DNS" swimtime="00:00:00.00" resultid="2574" heatid="5200" lane="6" entrytime="00:02:27.38" entrycourse="LCM" />
                <RESULT eventid="1251" points="483" swimtime="00:02:39.87" resultid="2575" heatid="5320" lane="7" entrytime="00:02:33.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.03" />
                    <SPLIT distance="100" swimtime="00:01:15.59" />
                    <SPLIT distance="150" swimtime="00:01:57.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="562" swimtime="00:00:31.44" resultid="2576" heatid="5371" lane="8" entrytime="00:00:31.55" entrycourse="LCM" />
                <RESULT eventid="2320" points="559" swimtime="00:01:09.01" resultid="5959" heatid="6414" lane="1" entrytime="00:01:09.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.91" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Chaim" birthdate="2011-05-29" gender="F" nation="BRA" license="370662" swrid="5409721" athleteid="2629" externalid="370662">
              <RESULTS>
                <RESULT eventid="1096" points="362" swimtime="00:00:33.11" resultid="2630" heatid="5098" lane="8" entrytime="00:00:33.29" entrycourse="LCM" />
                <RESULT eventid="1112" points="301" swimtime="00:02:48.29" resultid="2631" heatid="5138" lane="6" entrytime="00:02:49.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="100" swimtime="00:01:20.62" />
                    <SPLIT distance="150" swimtime="00:02:06.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="246" swimtime="00:01:31.49" resultid="2632" heatid="5241" lane="4" entrytime="00:01:31.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="331" swimtime="00:01:14.73" resultid="2633" heatid="5202" lane="2" entrytime="00:01:16.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="295" swimtime="00:00:40.34" resultid="2634" heatid="5292" lane="6" entrytime="00:00:42.99" entrycourse="LCM" />
                <RESULT eventid="1259" points="209" swimtime="00:00:41.16" resultid="2635" heatid="5323" lane="5" entrytime="00:00:39.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carina" lastname="Costa Profeta" birthdate="2008-03-20" gender="F" nation="BRA" license="366964" swrid="5591584" athleteid="2584" externalid="366964">
              <RESULTS>
                <RESULT eventid="1080" points="491" swimtime="00:01:21.25" resultid="2585" heatid="5069" lane="2" entrytime="00:01:19.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="468" swimtime="00:00:30.39" resultid="2586" heatid="5103" lane="5" entrytime="00:00:29.73" entrycourse="LCM" />
                <RESULT eventid="1215" points="370" swimtime="00:00:37.40" resultid="2587" heatid="5290" lane="4" />
                <RESULT eventid="1259" points="462" swimtime="00:00:31.60" resultid="2588" heatid="5326" lane="2" entrytime="00:00:32.88" entrycourse="LCM" />
                <RESULT eventid="1305" points="514" swimtime="00:00:36.38" resultid="2589" heatid="5377" lane="5" entrytime="00:00:35.61" entrycourse="LCM" />
                <RESULT eventid="2312" swimtime="00:00:00.00" resultid="5947" entrytime="00:01:21.25" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Biason Santana" birthdate="2009-01-21" gender="M" nation="BRA" license="366969" swrid="5317765" athleteid="2606" externalid="366969">
              <RESULTS>
                <RESULT eventid="1104" points="462" swimtime="00:00:27.04" resultid="2607" heatid="5123" lane="5" entrytime="00:00:27.68" entrycourse="LCM" />
                <RESULT eventid="1135" points="476" swimtime="00:01:03.31" resultid="2608" heatid="5174" lane="3" entrytime="00:01:02.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="470" swimtime="00:01:00.24" resultid="2609" heatid="5227" lane="1" entrytime="00:01:01.25" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="516" swimtime="00:00:27.76" resultid="2610" heatid="5335" lane="7" entrytime="00:00:28.72" entrycourse="LCM" />
                <RESULT eventid="1293" points="372" swimtime="00:02:33.39" resultid="2611" heatid="5359" lane="8" entrytime="00:02:38.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.70" />
                    <SPLIT distance="100" swimtime="00:01:11.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Campelo" birthdate="2011-09-12" gender="M" nation="BRA" license="366963" swrid="5588742" athleteid="2617" externalid="366963">
              <RESULTS>
                <RESULT eventid="1104" points="514" swimtime="00:00:26.10" resultid="2618" heatid="5120" lane="5" entrytime="00:00:26.49" entrycourse="LCM" />
                <RESULT eventid="1120" points="420" swimtime="00:02:16.15" resultid="2619" heatid="5147" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                    <SPLIT distance="100" swimtime="00:01:06.79" />
                    <SPLIT distance="150" swimtime="00:01:42.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="506" swimtime="00:00:58.80" resultid="2620" heatid="5223" lane="3" entrytime="00:00:57.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="404" swimtime="00:00:31.84" resultid="2621" heatid="5286" lane="7" entrytime="00:00:31.97" entrycourse="LCM" />
                <RESULT eventid="1267" points="399" swimtime="00:00:30.24" resultid="2622" heatid="5333" lane="4" entrytime="00:00:30.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietro" lastname="Nabas De Assis" birthdate="2011-07-09" gender="M" nation="BRA" license="366968" swrid="5603878" athleteid="2623" externalid="366968">
              <RESULTS>
                <RESULT eventid="1088" points="339" swimtime="00:01:21.51" resultid="2624" heatid="5082" lane="5" entrytime="00:01:18.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="302" swimtime="00:02:31.88" resultid="2625" heatid="5147" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                    <SPLIT distance="100" swimtime="00:01:12.87" />
                    <SPLIT distance="150" swimtime="00:01:52.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="269" swimtime="00:06:15.26" resultid="2626" heatid="5275" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.60" />
                    <SPLIT distance="100" swimtime="00:01:25.85" />
                    <SPLIT distance="150" swimtime="00:02:17.36" />
                    <SPLIT distance="200" swimtime="00:03:06.75" />
                    <SPLIT distance="300" swimtime="00:04:50.46" />
                    <SPLIT distance="350" swimtime="00:05:33.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="274" swimtime="00:03:13.05" resultid="2627" heatid="5318" lane="7" entrytime="00:02:56.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.35" />
                    <SPLIT distance="100" swimtime="00:01:31.45" />
                    <SPLIT distance="150" swimtime="00:02:23.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="382" swimtime="00:00:35.74" resultid="2628" heatid="5368" lane="6" entrytime="00:00:36.22" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mochiutti Carneiro" birthdate="2010-04-22" gender="F" nation="BRA" license="370670" swrid="5588817" athleteid="2643" externalid="370670">
              <RESULTS>
                <RESULT eventid="1096" points="478" swimtime="00:00:30.18" resultid="2644" heatid="5100" lane="7" entrytime="00:00:29.92" entrycourse="LCM" />
                <RESULT eventid="1128" points="337" swimtime="00:01:19.69" resultid="2645" heatid="5160" lane="3" entrytime="00:01:13.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="478" swimtime="00:02:24.27" resultid="2646" heatid="5141" lane="1" entrytime="00:02:24.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                    <SPLIT distance="100" swimtime="00:01:10.91" />
                    <SPLIT distance="150" swimtime="00:01:48.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="488" swimtime="00:01:05.66" resultid="2647" heatid="5205" lane="5" entrytime="00:01:04.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="332" swimtime="00:06:23.89" resultid="2648" heatid="5279" lane="6" entrytime="00:06:32.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                    <SPLIT distance="100" swimtime="00:01:21.91" />
                    <SPLIT distance="150" swimtime="00:02:17.04" />
                    <SPLIT distance="200" swimtime="00:03:08.72" />
                    <SPLIT distance="250" swimtime="00:04:05.68" />
                    <SPLIT distance="300" swimtime="00:05:00.72" />
                    <SPLIT distance="350" swimtime="00:05:43.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="390" swimtime="00:00:33.42" resultid="2649" heatid="5326" lane="1" entrytime="00:00:33.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felype" lastname="Gongora Zago" birthdate="2011-09-14" gender="M" nation="BRA" license="392099" swrid="5603848" athleteid="2650" externalid="392099">
              <RESULTS>
                <RESULT eventid="1104" points="241" swimtime="00:00:33.56" resultid="2651" heatid="5116" lane="8" entrytime="00:00:34.34" entrycourse="LCM" />
                <RESULT eventid="1151" points="176" swimtime="00:03:23.23" resultid="2652" heatid="5192" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.25" />
                    <SPLIT distance="100" swimtime="00:01:34.20" />
                    <SPLIT distance="150" swimtime="00:02:40.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="251" swimtime="00:01:14.26" resultid="2653" heatid="5219" lane="2" entrytime="00:01:14.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="196" swimtime="00:00:40.52" resultid="2654" heatid="5283" lane="5" entrytime="00:00:44.70" entrycourse="LCM" />
                <RESULT eventid="1267" points="216" swimtime="00:00:37.06" resultid="2655" heatid="5330" lane="4" entrytime="00:00:51.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Quental De Meireles" birthdate="2008-11-20" gender="M" nation="BRA" license="392103" swrid="5603898" athleteid="2662" externalid="392103">
              <RESULTS>
                <RESULT eventid="1088" points="333" swimtime="00:01:22.06" resultid="2663" heatid="5083" lane="5" entrytime="00:01:22.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="387" swimtime="00:00:28.67" resultid="2664" heatid="5121" lane="4" entrytime="00:00:30.32" entrycourse="LCM" />
                <RESULT eventid="1135" points="371" swimtime="00:01:08.80" resultid="2665" heatid="5172" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="393" swimtime="00:00:30.39" resultid="2666" heatid="5334" lane="8" entrytime="00:00:29.96" entrycourse="LCM" />
                <RESULT eventid="1297" points="375" swimtime="00:00:35.96" resultid="2667" heatid="5368" lane="2" entrytime="00:00:36.80" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Marques Picolo Vinha" birthdate="2010-07-01" gender="M" nation="BRA" license="366990" swrid="5603869" athleteid="2674" externalid="366990">
              <RESULTS>
                <RESULT eventid="1104" points="358" swimtime="00:00:29.43" resultid="2675" heatid="5117" lane="4" entrytime="00:00:30.22" entrycourse="LCM" />
                <RESULT eventid="1120" points="301" swimtime="00:02:32.16" resultid="2676" heatid="5150" lane="7" entrytime="00:02:27.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                    <SPLIT distance="100" swimtime="00:01:11.69" />
                    <SPLIT distance="150" swimtime="00:01:51.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="355" swimtime="00:01:06.12" resultid="2677" heatid="5221" lane="6" entrytime="00:01:05.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="292" swimtime="00:11:20.76" resultid="2678" heatid="5297" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.35" />
                    <SPLIT distance="100" swimtime="00:01:15.85" />
                    <SPLIT distance="150" swimtime="00:01:59.21" />
                    <SPLIT distance="200" swimtime="00:02:43.09" />
                    <SPLIT distance="250" swimtime="00:03:24.76" />
                    <SPLIT distance="300" swimtime="00:04:07.18" />
                    <SPLIT distance="350" swimtime="00:04:50.88" />
                    <SPLIT distance="400" swimtime="00:05:35.04" />
                    <SPLIT distance="450" swimtime="00:06:19.28" />
                    <SPLIT distance="500" swimtime="00:07:04.96" />
                    <SPLIT distance="550" swimtime="00:07:48.70" />
                    <SPLIT distance="600" swimtime="00:08:32.37" />
                    <SPLIT distance="650" swimtime="00:09:17.50" />
                    <SPLIT distance="700" swimtime="00:09:59.62" />
                    <SPLIT distance="750" swimtime="00:10:39.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="307" swimtime="00:00:33.01" resultid="2679" heatid="5332" lane="8" entrytime="00:00:35.00" entrycourse="LCM" />
                <RESULT eventid="1297" points="258" swimtime="00:00:40.72" resultid="2680" heatid="5364" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Pacheco" birthdate="2006-12-20" gender="M" nation="BRA" license="336850" swrid="5603854" athleteid="2577" externalid="336850">
              <RESULTS>
                <RESULT eventid="1104" points="476" swimtime="00:00:26.78" resultid="2578" heatid="5128" lane="3" entrytime="00:00:27.07" entrycourse="LCM" />
                <RESULT eventid="1135" points="458" swimtime="00:01:04.11" resultid="2579" heatid="5177" lane="8" entrytime="00:01:03.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="508" swimtime="00:00:58.70" resultid="2580" heatid="5231" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="335" swimtime="00:05:48.91" resultid="2581" heatid="5276" lane="5" entrytime="00:05:27.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                    <SPLIT distance="100" swimtime="00:01:11.67" />
                    <SPLIT distance="150" swimtime="00:01:56.45" />
                    <SPLIT distance="200" swimtime="00:02:41.55" />
                    <SPLIT distance="250" swimtime="00:03:35.03" />
                    <SPLIT distance="300" swimtime="00:04:27.46" />
                    <SPLIT distance="350" swimtime="00:05:07.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="474" swimtime="00:00:28.55" resultid="2582" heatid="5335" lane="6" entrytime="00:00:28.20" entrycourse="LCM" />
                <RESULT eventid="1297" points="387" swimtime="00:00:35.59" resultid="2583" heatid="5368" lane="7" entrytime="00:00:36.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Camila Cuenca" birthdate="2005-10-06" gender="F" nation="BRA" license="308081" swrid="5357445" athleteid="2568" externalid="308081">
              <RESULTS>
                <RESULT eventid="1096" points="474" swimtime="00:00:30.26" resultid="2569" heatid="5106" lane="2" entrytime="00:00:29.59" entrycourse="LCM" />
                <RESULT eventid="1275" points="377" swimtime="00:02:50.44" resultid="2570" heatid="5342" lane="3" entrytime="00:02:46.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.77" />
                    <SPLIT distance="100" swimtime="00:01:24.37" />
                    <SPLIT distance="150" swimtime="00:02:08.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="326" swimtime="00:00:42.33" resultid="2571" heatid="5375" lane="6" entrytime="00:00:40.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Donato De Morais" birthdate="2009-03-28" gender="F" nation="BRA" license="345588" swrid="5485198" athleteid="2590" externalid="345588">
              <RESULTS>
                <RESULT eventid="1096" points="384" swimtime="00:00:32.46" resultid="2591" heatid="5102" lane="1" entrytime="00:00:32.51" entrycourse="LCM" />
                <RESULT eventid="1175" points="375" swimtime="00:01:19.49" resultid="2592" heatid="5246" lane="4" entrytime="00:01:18.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="398" swimtime="00:00:36.51" resultid="2593" heatid="5294" lane="7" entrytime="00:00:36.43" entrycourse="LCM" />
                <RESULT eventid="1275" points="312" swimtime="00:03:01.39" resultid="2594" heatid="5341" lane="3" entrytime="00:02:50.64" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Antonio Mendes" birthdate="2008-12-04" gender="M" nation="BRA" license="366962" swrid="5196287" athleteid="2600" externalid="366962">
              <RESULTS>
                <RESULT eventid="1088" points="567" swimtime="00:01:08.69" resultid="2601" heatid="5085" lane="3" entrytime="00:01:09.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="461" swimtime="00:02:27.54" resultid="2602" heatid="5197" lane="3" entrytime="00:02:28.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                    <SPLIT distance="100" swimtime="00:01:08.99" />
                    <SPLIT distance="150" swimtime="00:01:49.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="443" swimtime="00:00:30.89" resultid="2603" heatid="5286" lane="2" entrytime="00:00:31.88" entrycourse="LCM" />
                <RESULT eventid="1251" points="539" swimtime="00:02:34.11" resultid="2604" heatid="5320" lane="1" entrytime="00:02:34.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:13.81" />
                    <SPLIT distance="150" swimtime="00:01:53.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="591" swimtime="00:00:30.92" resultid="2605" heatid="5371" lane="6" entrytime="00:00:30.98" entrycourse="LCM" />
                <RESULT eventid="2320" points="552" swimtime="00:01:09.30" resultid="5958" heatid="6414" lane="7" entrytime="00:01:08.69">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wellington" lastname="De Lima" birthdate="2008-03-01" gender="M" nation="BRA" license="370024" swrid="5470912" athleteid="2537" externalid="370024">
              <RESULTS>
                <RESULT eventid="1104" points="514" swimtime="00:00:26.09" resultid="2538" heatid="5125" lane="7" entrytime="00:00:26.30" entrycourse="LCM" />
                <RESULT eventid="1135" points="371" swimtime="00:01:08.77" resultid="2539" heatid="5174" lane="8" entrytime="00:01:07.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="364" swimtime="00:01:12.26" resultid="2540" heatid="5260" lane="7" entrytime="00:01:11.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="544" swimtime="00:00:57.38" resultid="2541" heatid="5229" lane="7" entrytime="00:00:57.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="428" swimtime="00:00:31.23" resultid="2542" heatid="5286" lane="1" entrytime="00:00:32.24" entrycourse="LCM" />
                <RESULT eventid="1267" points="438" swimtime="00:00:29.31" resultid="2543" heatid="5334" lane="4" entrytime="00:00:28.83" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Ficher Delmont Pais" birthdate="2010-07-15" gender="M" nation="BRA" license="338533" swrid="5588701" athleteid="2530" externalid="338533">
              <RESULTS>
                <RESULT eventid="1104" points="557" swimtime="00:00:25.41" resultid="2531" heatid="5120" lane="4" entrytime="00:00:25.14" entrycourse="LCM" />
                <RESULT eventid="1135" points="538" swimtime="00:01:00.80" resultid="2532" heatid="5171" lane="4" entrytime="00:00:59.28" entrycourse="LCM" />
                <RESULT eventid="1120" points="551" swimtime="00:02:04.41" resultid="2533" heatid="5152" lane="3" entrytime="00:02:08.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.06" />
                    <SPLIT distance="100" swimtime="00:01:00.63" />
                    <SPLIT distance="150" swimtime="00:01:32.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="610" swimtime="00:00:55.23" resultid="2534" heatid="5223" lane="4" entrytime="00:00:54.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="559" swimtime="00:00:27.02" resultid="2535" heatid="5337" lane="2" entrytime="00:00:27.28" entrycourse="LCM" />
                <RESULT eventid="1293" points="364" swimtime="00:02:34.48" resultid="2536" heatid="5359" lane="2" entrytime="00:02:33.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.85" />
                    <SPLIT distance="100" swimtime="00:01:14.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Inoue" birthdate="2008-10-31" gender="F" nation="BRA" license="378348" swrid="5603856" athleteid="2612" externalid="378348">
              <RESULTS>
                <RESULT eventid="1096" points="430" swimtime="00:00:31.26" resultid="2613" heatid="5102" lane="3" entrytime="00:00:31.67" entrycourse="LCM" />
                <RESULT eventid="1175" points="301" swimtime="00:01:25.53" resultid="2614" heatid="5246" lane="7" entrytime="00:01:24.40" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="354" swimtime="00:00:37.95" resultid="2615" heatid="5293" lane="6" entrytime="00:00:37.96" entrycourse="LCM" />
                <RESULT eventid="1259" points="299" swimtime="00:00:36.51" resultid="2616" heatid="5324" lane="5" entrytime="00:00:35.76" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Garcia Cavalcante" birthdate="2008-08-11" gender="M" nation="BRA" license="369676" swrid="5603841" athleteid="2549" externalid="369676">
              <RESULTS>
                <RESULT eventid="1088" points="344" swimtime="00:01:21.14" resultid="2550" heatid="5084" lane="6" entrytime="00:01:16.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="375" swimtime="00:02:21.33" resultid="2551" heatid="5154" lane="2" entrytime="00:02:19.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:07.71" />
                    <SPLIT distance="150" swimtime="00:01:44.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" status="DNS" swimtime="00:00:00.00" resultid="2552" heatid="5224" lane="6" />
                <RESULT eventid="1251" status="DNS" swimtime="00:00:00.00" resultid="2553" heatid="5319" lane="7" entrytime="00:02:43.93" entrycourse="LCM" />
                <RESULT eventid="1297" points="388" swimtime="00:00:35.56" resultid="2554" heatid="5369" lane="2" entrytime="00:00:35.06" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Batista Sanchez" birthdate="2009-05-22" gender="M" nation="BRA" license="370668" swrid="5255779" athleteid="2544" externalid="370668">
              <RESULTS>
                <RESULT eventid="1088" points="437" swimtime="00:01:14.92" resultid="2545" heatid="5084" lane="5" entrytime="00:01:15.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="345" swimtime="00:01:10.50" resultid="2546" heatid="5173" lane="2" entrytime="00:01:14.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="411" swimtime="00:02:48.66" resultid="2547" heatid="5318" lane="5" entrytime="00:02:45.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.13" />
                    <SPLIT distance="100" swimtime="00:01:20.78" />
                    <SPLIT distance="150" swimtime="00:02:05.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="452" swimtime="00:00:33.80" resultid="2548" heatid="5368" lane="4" entrytime="00:00:35.65" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1237" points="471" swimtime="00:04:01.90" resultid="2685" heatid="5308" lane="6" entrytime="00:04:05.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.93" />
                    <SPLIT distance="100" swimtime="00:00:58.14" />
                    <SPLIT distance="150" swimtime="00:01:25.30" />
                    <SPLIT distance="200" swimtime="00:01:56.75" />
                    <SPLIT distance="250" swimtime="00:02:26.05" />
                    <SPLIT distance="300" swimtime="00:02:59.10" />
                    <SPLIT distance="350" swimtime="00:03:28.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2537" number="1" />
                    <RELAYPOSITION athleteid="2600" number="2" />
                    <RELAYPOSITION athleteid="2549" number="3" />
                    <RELAYPOSITION athleteid="2662" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1338" points="462" swimtime="00:04:27.43" resultid="2688" heatid="5388" lane="3" entrytime="00:04:34.34">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.57" />
                    <SPLIT distance="100" swimtime="00:01:10.70" />
                    <SPLIT distance="150" swimtime="00:01:42.15" />
                    <SPLIT distance="200" swimtime="00:02:18.67" />
                    <SPLIT distance="250" swimtime="00:02:49.34" />
                    <SPLIT distance="300" swimtime="00:03:24.84" />
                    <SPLIT distance="350" swimtime="00:03:53.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2537" number="1" />
                    <RELAYPOSITION athleteid="2600" number="2" />
                    <RELAYPOSITION athleteid="2662" number="3" />
                    <RELAYPOSITION athleteid="2549" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1231" points="357" swimtime="00:04:25.21" resultid="2686" heatid="5305" lane="2" entrytime="00:04:38.72">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.00" />
                    <SPLIT distance="100" swimtime="00:00:58.54" />
                    <SPLIT distance="150" swimtime="00:01:28.97" />
                    <SPLIT distance="200" swimtime="00:02:04.24" />
                    <SPLIT distance="250" swimtime="00:02:39.05" />
                    <SPLIT distance="300" swimtime="00:03:18.08" />
                    <SPLIT distance="350" swimtime="00:03:49.59" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2617" number="1" />
                    <RELAYPOSITION athleteid="2623" number="2" />
                    <RELAYPOSITION athleteid="2650" number="3" />
                    <RELAYPOSITION athleteid="2555" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 18:59), Na volta dos 250m (Revezamento Medley, Borboleta)." eventid="1332" status="DSQ" swimtime="00:05:15.79" resultid="2687" heatid="5385" lane="2" entrytime="00:05:23.55">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.08" />
                    <SPLIT distance="100" swimtime="00:01:09.02" />
                    <SPLIT distance="150" swimtime="00:01:48.82" />
                    <SPLIT distance="200" swimtime="00:02:34.87" />
                    <SPLIT distance="250" swimtime="00:03:12.45" />
                    <SPLIT distance="350" swimtime="00:04:36.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2617" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="2623" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="2555" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="2650" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1221" points="410" swimtime="00:04:39.73" resultid="2681" heatid="5302" lane="6" entrytime="00:04:41.23">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.57" />
                    <SPLIT distance="100" swimtime="00:01:07.67" />
                    <SPLIT distance="150" swimtime="00:01:39.74" />
                    <SPLIT distance="200" swimtime="00:02:14.20" />
                    <SPLIT distance="250" swimtime="00:02:48.83" />
                    <SPLIT distance="300" swimtime="00:03:28.19" />
                    <SPLIT distance="350" swimtime="00:04:01.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2656" number="1" />
                    <RELAYPOSITION athleteid="2643" number="2" />
                    <RELAYPOSITION athleteid="2629" number="3" />
                    <RELAYPOSITION athleteid="2636" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1322" points="392" swimtime="00:05:14.63" resultid="2684" heatid="5382" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                    <SPLIT distance="150" swimtime="00:02:03.61" />
                    <SPLIT distance="200" swimtime="00:02:52.17" />
                    <SPLIT distance="250" swimtime="00:03:27.87" />
                    <SPLIT distance="300" swimtime="00:04:08.69" />
                    <SPLIT distance="350" swimtime="00:04:39.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2636" number="1" />
                    <RELAYPOSITION athleteid="2668" number="2" />
                    <RELAYPOSITION athleteid="2643" number="3" />
                    <RELAYPOSITION athleteid="2656" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="F" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1225" points="377" swimtime="00:04:47.73" resultid="2682" heatid="5304" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:14.90" />
                    <SPLIT distance="150" swimtime="00:01:46.78" />
                    <SPLIT distance="200" swimtime="00:02:24.07" />
                    <SPLIT distance="250" swimtime="00:02:57.66" />
                    <SPLIT distance="300" swimtime="00:03:35.44" />
                    <SPLIT distance="350" swimtime="00:04:09.12" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2595" number="1" />
                    <RELAYPOSITION athleteid="2584" number="2" />
                    <RELAYPOSITION athleteid="2590" number="3" />
                    <RELAYPOSITION athleteid="2612" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1326" points="359" swimtime="00:05:23.92" resultid="2683" heatid="5384" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.96" />
                    <SPLIT distance="100" swimtime="00:01:19.50" />
                    <SPLIT distance="150" swimtime="00:01:58.76" />
                    <SPLIT distance="200" swimtime="00:02:44.17" />
                    <SPLIT distance="250" swimtime="00:03:22.38" />
                    <SPLIT distance="300" swimtime="00:04:12.84" />
                    <SPLIT distance="350" swimtime="00:04:46.18" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2590" number="1" />
                    <RELAYPOSITION athleteid="2584" number="2" />
                    <RELAYPOSITION athleteid="2595" number="3" />
                    <RELAYPOSITION athleteid="2612" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1287" points="437" swimtime="00:04:46.55" resultid="2689" heatid="5354" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                    <SPLIT distance="100" swimtime="00:01:06.96" />
                    <SPLIT distance="150" swimtime="00:01:45.05" />
                    <SPLIT distance="200" swimtime="00:02:29.66" />
                    <SPLIT distance="250" swimtime="00:03:00.42" />
                    <SPLIT distance="300" swimtime="00:03:37.42" />
                    <SPLIT distance="350" swimtime="00:04:09.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2600" number="1" />
                    <RELAYPOSITION athleteid="2584" number="2" />
                    <RELAYPOSITION athleteid="2662" number="3" />
                    <RELAYPOSITION athleteid="2612" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1285" points="399" swimtime="00:04:55.46" resultid="2690" heatid="5353" lane="2" entrytime="00:04:38.17">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.79" />
                    <SPLIT distance="150" swimtime="00:01:56.57" />
                    <SPLIT distance="200" swimtime="00:02:36.43" />
                    <SPLIT distance="250" swimtime="00:03:05.98" />
                    <SPLIT distance="300" swimtime="00:03:40.49" />
                    <SPLIT distance="350" swimtime="00:04:14.94" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2590" number="1" />
                    <RELAYPOSITION athleteid="2544" number="2" />
                    <RELAYPOSITION athleteid="2606" number="3" />
                    <RELAYPOSITION athleteid="2595" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1283" points="381" swimtime="00:05:00.01" resultid="2691" heatid="5352" lane="3" entrytime="00:04:52.99">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.84" />
                    <SPLIT distance="100" swimtime="00:01:18.13" />
                    <SPLIT distance="150" swimtime="00:01:54.80" />
                    <SPLIT distance="200" swimtime="00:02:35.82" />
                    <SPLIT distance="250" swimtime="00:03:12.88" />
                    <SPLIT distance="300" swimtime="00:03:54.95" />
                    <SPLIT distance="350" swimtime="00:04:25.53" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2636" number="1" />
                    <RELAYPOSITION athleteid="2530" number="2" />
                    <RELAYPOSITION athleteid="2643" number="3" />
                    <RELAYPOSITION athleteid="2674" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="APAN/MARINGÁ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1281" points="373" swimtime="00:05:02.09" resultid="2692" heatid="5351" lane="5" entrytime="00:04:58.04">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:16.61" />
                    <SPLIT distance="150" swimtime="00:01:57.21" />
                    <SPLIT distance="200" swimtime="00:02:39.46" />
                    <SPLIT distance="250" swimtime="00:03:11.84" />
                    <SPLIT distance="300" swimtime="00:03:49.27" />
                    <SPLIT distance="350" swimtime="00:04:22.66" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2656" number="1" />
                    <RELAYPOSITION athleteid="2623" number="2" />
                    <RELAYPOSITION athleteid="2617" number="3" />
                    <RELAYPOSITION athleteid="2629" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="36" nation="BRA" region="PR" clubid="3236" swrid="93753" name="Associação Atlética Comercial" shortname="Comercial Cascavel">
          <ATHLETES>
            <ATHLETE firstname="Raul" lastname="Bonamigo" birthdate="2010-12-01" gender="M" nation="BRA" license="344397" swrid="5588559" athleteid="3386" externalid="344397">
              <RESULTS>
                <RESULT eventid="1072" points="465" swimtime="00:04:43.96" resultid="3387" heatid="5059" lane="2" entrytime="00:04:44.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:06.64" />
                    <SPLIT distance="150" swimtime="00:01:42.58" />
                    <SPLIT distance="200" swimtime="00:02:19.04" />
                    <SPLIT distance="250" swimtime="00:02:55.23" />
                    <SPLIT distance="300" swimtime="00:03:32.09" />
                    <SPLIT distance="350" swimtime="00:04:08.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="443" swimtime="00:02:29.54" resultid="3388" heatid="5195" lane="2" entrytime="00:02:32.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.44" />
                    <SPLIT distance="100" swimtime="00:01:10.39" />
                    <SPLIT distance="150" swimtime="00:01:55.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="451" swimtime="00:01:07.27" resultid="3389" heatid="5257" lane="2" entrytime="00:01:12.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="441" swimtime="00:05:18.46" resultid="3390" heatid="5276" lane="4" entrytime="00:05:23.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.16" />
                    <SPLIT distance="100" swimtime="00:01:12.73" />
                    <SPLIT distance="150" swimtime="00:01:53.67" />
                    <SPLIT distance="200" swimtime="00:02:32.88" />
                    <SPLIT distance="250" swimtime="00:03:20.10" />
                    <SPLIT distance="300" swimtime="00:04:08.51" />
                    <SPLIT distance="350" swimtime="00:04:45.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="373" swimtime="00:00:32.71" resultid="3391" heatid="5283" lane="1" />
                <RESULT eventid="1277" points="435" swimtime="00:02:27.61" resultid="3392" heatid="5347" lane="6" entrytime="00:02:25.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:11.94" />
                    <SPLIT distance="150" swimtime="00:01:50.60" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Assakura" birthdate="2010-06-29" gender="F" nation="BRA" license="376473" swrid="5596868" athleteid="3379" externalid="376473">
              <RESULTS>
                <RESULT eventid="1080" points="416" swimtime="00:01:25.88" resultid="3380" heatid="5067" lane="7" entrytime="00:01:23.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" points="440" swimtime="00:05:09.31" resultid="3381" heatid="5049" lane="5" entrytime="00:05:19.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.27" />
                    <SPLIT distance="100" swimtime="00:01:09.29" />
                    <SPLIT distance="150" swimtime="00:01:49.58" />
                    <SPLIT distance="200" swimtime="00:02:30.02" />
                    <SPLIT distance="250" swimtime="00:03:10.96" />
                    <SPLIT distance="300" swimtime="00:03:50.32" />
                    <SPLIT distance="350" swimtime="00:04:29.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="465" swimtime="00:02:25.62" resultid="3382" heatid="5140" lane="8" entrytime="00:02:29.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                    <SPLIT distance="100" swimtime="00:01:09.60" />
                    <SPLIT distance="150" swimtime="00:01:47.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="445" swimtime="00:02:45.14" resultid="3383" heatid="5188" lane="6" entrytime="00:02:44.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.16" />
                    <SPLIT distance="100" swimtime="00:01:19.99" />
                    <SPLIT distance="150" swimtime="00:02:08.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="423" swimtime="00:01:16.36" resultid="3384" heatid="5244" lane="7" entrytime="00:01:16.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="464" swimtime="00:02:57.64" resultid="3385" heatid="5314" lane="2" entrytime="00:02:55.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.50" />
                    <SPLIT distance="100" swimtime="00:01:24.07" />
                    <SPLIT distance="150" swimtime="00:02:10.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Gamero Prado" birthdate="2007-05-16" gender="F" nation="BRA" license="305973" swrid="5596903" athleteid="3248" externalid="305973">
              <RESULTS>
                <RESULT eventid="1128" points="398" swimtime="00:01:15.37" resultid="3249" heatid="5162" lane="5" entrytime="00:01:15.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="435" swimtime="00:10:39.76" resultid="3250" heatid="5273" lane="6" entrytime="00:10:25.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.61" />
                    <SPLIT distance="100" swimtime="00:01:13.31" />
                    <SPLIT distance="150" swimtime="00:01:52.51" />
                    <SPLIT distance="200" swimtime="00:02:32.85" />
                    <SPLIT distance="250" swimtime="00:03:13.27" />
                    <SPLIT distance="300" swimtime="00:03:54.03" />
                    <SPLIT distance="350" swimtime="00:04:35.31" />
                    <SPLIT distance="400" swimtime="00:05:16.81" />
                    <SPLIT distance="450" swimtime="00:05:58.62" />
                    <SPLIT distance="500" swimtime="00:06:39.91" />
                    <SPLIT distance="550" swimtime="00:07:20.47" />
                    <SPLIT distance="600" swimtime="00:08:01.72" />
                    <SPLIT distance="650" swimtime="00:08:42.35" />
                    <SPLIT distance="700" swimtime="00:09:23.48" />
                    <SPLIT distance="750" swimtime="00:10:04.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="359" swimtime="00:06:13.89" resultid="3251" heatid="5279" lane="4" entrytime="00:06:04.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.00" />
                    <SPLIT distance="100" swimtime="00:01:19.77" />
                    <SPLIT distance="150" swimtime="00:02:07.41" />
                    <SPLIT distance="200" swimtime="00:02:54.81" />
                    <SPLIT distance="250" swimtime="00:03:53.99" />
                    <SPLIT distance="300" swimtime="00:04:52.48" />
                    <SPLIT distance="350" swimtime="00:05:33.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="390" swimtime="00:00:33.42" resultid="3252" heatid="5325" lane="1" entrytime="00:00:35.14" entrycourse="LCM" />
                <RESULT eventid="1279" points="400" swimtime="00:20:48.90" resultid="3253" heatid="5350" lane="8" entrytime="00:20:42.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.79" />
                    <SPLIT distance="100" swimtime="00:01:15.64" />
                    <SPLIT distance="150" swimtime="00:01:56.91" />
                    <SPLIT distance="200" swimtime="00:02:39.00" />
                    <SPLIT distance="250" swimtime="00:03:20.59" />
                    <SPLIT distance="300" swimtime="00:04:03.20" />
                    <SPLIT distance="350" swimtime="00:04:45.61" />
                    <SPLIT distance="400" swimtime="00:05:28.90" />
                    <SPLIT distance="450" swimtime="00:06:12.15" />
                    <SPLIT distance="500" swimtime="00:06:55.80" />
                    <SPLIT distance="550" swimtime="00:07:39.20" />
                    <SPLIT distance="600" swimtime="00:08:22.50" />
                    <SPLIT distance="650" swimtime="00:09:06.08" />
                    <SPLIT distance="700" swimtime="00:09:49.79" />
                    <SPLIT distance="750" swimtime="00:10:33.72" />
                    <SPLIT distance="800" swimtime="00:11:15.12" />
                    <SPLIT distance="850" swimtime="00:11:56.45" />
                    <SPLIT distance="900" swimtime="00:12:38.58" />
                    <SPLIT distance="950" swimtime="00:13:20.34" />
                    <SPLIT distance="1000" swimtime="00:14:02.12" />
                    <SPLIT distance="1050" swimtime="00:14:44.04" />
                    <SPLIT distance="1100" swimtime="00:15:24.43" />
                    <SPLIT distance="1150" swimtime="00:16:05.84" />
                    <SPLIT distance="1200" swimtime="00:16:47.63" />
                    <SPLIT distance="1250" swimtime="00:17:28.90" />
                    <SPLIT distance="1300" swimtime="00:18:10.20" />
                    <SPLIT distance="1350" swimtime="00:18:50.47" />
                    <SPLIT distance="1400" swimtime="00:19:30.42" />
                    <SPLIT distance="1450" swimtime="00:20:10.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1295" points="326" swimtime="00:02:56.90" resultid="3254" heatid="5362" lane="6" entrytime="00:02:49.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.66" />
                    <SPLIT distance="100" swimtime="00:01:23.91" />
                    <SPLIT distance="150" swimtime="00:02:13.56" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2328" swimtime="00:00:00.00" resultid="6005" entrytime="00:01:15.37" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hendrik" lastname="Alteiro Groenwold" birthdate="2011-03-23" gender="M" nation="BRA" license="365756" swrid="5588520" athleteid="3309" externalid="365756">
              <RESULTS>
                <RESULT eventid="1072" points="494" swimtime="00:04:38.26" resultid="3310" heatid="5058" lane="5" entrytime="00:04:56.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.46" />
                    <SPLIT distance="100" swimtime="00:01:05.08" />
                    <SPLIT distance="150" swimtime="00:01:40.48" />
                    <SPLIT distance="200" swimtime="00:02:16.70" />
                    <SPLIT distance="250" swimtime="00:02:52.22" />
                    <SPLIT distance="300" swimtime="00:03:28.97" />
                    <SPLIT distance="350" swimtime="00:04:03.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="491" swimtime="00:02:09.29" resultid="3311" heatid="5151" lane="3" entrytime="00:02:18.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.57" />
                    <SPLIT distance="100" swimtime="00:01:02.35" />
                    <SPLIT distance="150" swimtime="00:01:36.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="477" swimtime="00:01:06.04" resultid="3312" heatid="5258" lane="3" entrytime="00:01:06.70" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="443" swimtime="00:05:17.88" resultid="3313" heatid="5276" lane="3" entrytime="00:05:37.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.58" />
                    <SPLIT distance="100" swimtime="00:01:10.14" />
                    <SPLIT distance="150" swimtime="00:01:50.32" />
                    <SPLIT distance="200" swimtime="00:02:29.66" />
                    <SPLIT distance="250" swimtime="00:03:17.46" />
                    <SPLIT distance="300" swimtime="00:04:07.19" />
                    <SPLIT distance="350" swimtime="00:04:43.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="442" swimtime="00:02:26.85" resultid="3314" heatid="5346" lane="7" entrytime="00:02:33.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                    <SPLIT distance="100" swimtime="00:01:13.19" />
                    <SPLIT distance="150" swimtime="00:01:50.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1293" points="418" swimtime="00:02:27.54" resultid="3315" heatid="5359" lane="5" entrytime="00:02:26.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.62" />
                    <SPLIT distance="100" swimtime="00:01:10.65" />
                    <SPLIT distance="150" swimtime="00:01:50.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Bortoli Da Silva" birthdate="2010-09-30" gender="M" nation="BRA" license="365500" swrid="4675666" athleteid="3435" externalid="365500">
              <RESULTS>
                <RESULT eventid="1104" points="337" swimtime="00:00:30.03" resultid="3436" heatid="5114" lane="3" />
                <RESULT eventid="1135" points="310" swimtime="00:01:13.01" resultid="3437" heatid="5169" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="348" swimtime="00:01:06.61" resultid="3438" heatid="5218" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="356" swimtime="00:05:41.97" resultid="3439" heatid="5275" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.84" />
                    <SPLIT distance="100" swimtime="00:01:15.58" />
                    <SPLIT distance="150" swimtime="00:02:01.86" />
                    <SPLIT distance="200" swimtime="00:02:47.60" />
                    <SPLIT distance="250" swimtime="00:03:35.11" />
                    <SPLIT distance="300" swimtime="00:04:25.04" />
                    <SPLIT distance="350" swimtime="00:05:04.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="297" swimtime="00:00:33.37" resultid="3440" heatid="5329" lane="7" />
                <RESULT eventid="1297" points="306" swimtime="00:00:38.48" resultid="3441" heatid="5364" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Cordeiro Silva" birthdate="2011-09-04" gender="M" nation="BRA" license="380664" swrid="5596877" athleteid="3365" externalid="380664">
              <RESULTS>
                <RESULT eventid="1088" points="281" swimtime="00:01:26.74" resultid="3366" heatid="5080" lane="1" entrytime="00:01:32.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="266" swimtime="00:02:57.11" resultid="3367" heatid="5193" lane="3" entrytime="00:03:06.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.19" />
                    <SPLIT distance="100" swimtime="00:01:28.08" />
                    <SPLIT distance="150" swimtime="00:02:15.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="249" swimtime="00:01:14.42" resultid="3368" heatid="5219" lane="8" entrytime="00:01:17.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="277" swimtime="00:06:11.63" resultid="3369" heatid="5275" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.28" />
                    <SPLIT distance="100" swimtime="00:01:28.22" />
                    <SPLIT distance="150" swimtime="00:02:20.85" />
                    <SPLIT distance="200" swimtime="00:03:07.75" />
                    <SPLIT distance="250" swimtime="00:03:57.00" />
                    <SPLIT distance="300" swimtime="00:04:47.05" />
                    <SPLIT distance="350" swimtime="00:05:30.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="291" swimtime="00:03:09.14" resultid="3370" heatid="5316" lane="3" entrytime="00:03:18.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.72" />
                    <SPLIT distance="100" swimtime="00:01:32.64" />
                    <SPLIT distance="150" swimtime="00:02:21.42" />
                  </SPLITS>
                </RESULT>
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 16:52), Nos 50m." eventid="1297" status="DSQ" swimtime="00:00:39.36" resultid="3371" heatid="5367" lane="1" entrytime="00:00:40.75" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Tolentino Smarczewski" birthdate="2008-09-01" gender="M" nation="BRA" license="378818" swrid="5596941" athleteid="3358" externalid="378818">
              <RESULTS>
                <RESULT eventid="1088" points="390" swimtime="00:01:17.80" resultid="3359" heatid="5084" lane="7" entrytime="00:01:18.53" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="493" swimtime="00:02:09.08" resultid="3360" heatid="5155" lane="6" entrytime="00:02:11.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.63" />
                    <SPLIT distance="100" swimtime="00:01:03.41" />
                    <SPLIT distance="150" swimtime="00:01:36.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="482" swimtime="00:00:59.73" resultid="3361" heatid="5226" lane="4" entrytime="00:01:01.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="459" swimtime="00:09:45.72" resultid="3362" heatid="5299" lane="5" entrytime="00:09:41.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.10" />
                    <SPLIT distance="100" swimtime="00:01:07.75" />
                    <SPLIT distance="150" swimtime="00:01:44.25" />
                    <SPLIT distance="200" swimtime="00:02:21.48" />
                    <SPLIT distance="250" swimtime="00:02:59.06" />
                    <SPLIT distance="300" swimtime="00:03:36.59" />
                    <SPLIT distance="350" swimtime="00:04:14.13" />
                    <SPLIT distance="400" swimtime="00:04:51.84" />
                    <SPLIT distance="450" swimtime="00:05:29.09" />
                    <SPLIT distance="500" swimtime="00:06:06.23" />
                    <SPLIT distance="550" swimtime="00:06:44.15" />
                    <SPLIT distance="600" swimtime="00:07:20.59" />
                    <SPLIT distance="650" swimtime="00:07:57.66" />
                    <SPLIT distance="700" swimtime="00:08:34.55" />
                    <SPLIT distance="750" swimtime="00:09:11.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="393" swimtime="00:02:51.20" resultid="3363" heatid="5318" lane="3" entrytime="00:02:46.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.55" />
                    <SPLIT distance="100" swimtime="00:01:23.59" />
                    <SPLIT distance="150" swimtime="00:02:09.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="354" swimtime="00:00:36.68" resultid="3364" heatid="5364" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Do Prado Martins" birthdate="2008-10-17" gender="F" nation="BRA" license="369419" swrid="5596893" athleteid="3316" externalid="369419">
              <RESULTS>
                <RESULT eventid="1080" points="501" swimtime="00:01:20.70" resultid="3317" heatid="5069" lane="8" entrytime="00:01:21.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="533" swimtime="00:02:35.47" resultid="3318" heatid="5190" lane="5" entrytime="00:02:35.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                    <SPLIT distance="100" swimtime="00:01:12.00" />
                    <SPLIT distance="150" swimtime="00:01:57.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="500" swimtime="00:01:05.15" resultid="3319" heatid="5207" lane="3" entrytime="00:01:06.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="451" swimtime="00:05:46.60" resultid="3320" heatid="5280" lane="6" entrytime="00:05:35.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                    <SPLIT distance="100" swimtime="00:01:19.18" />
                    <SPLIT distance="150" swimtime="00:02:05.41" />
                    <SPLIT distance="200" swimtime="00:02:50.36" />
                    <SPLIT distance="250" swimtime="00:03:39.64" />
                    <SPLIT distance="300" swimtime="00:04:28.08" />
                    <SPLIT distance="350" swimtime="00:05:08.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="463" swimtime="00:00:31.56" resultid="3321" heatid="5321" lane="8" />
                <RESULT eventid="1305" points="502" swimtime="00:00:36.69" resultid="3322" heatid="5373" lane="7" />
                <RESULT eventid="2312" points="498" swimtime="00:01:20.89" resultid="5946" heatid="6416" lane="8" entrytime="00:01:20.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.57" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Sehn Uren" birthdate="2009-10-15" gender="F" nation="BRA" license="357159" swrid="5596937" athleteid="3281" externalid="357159">
              <RESULTS>
                <RESULT eventid="1080" points="353" swimtime="00:01:30.73" resultid="3282" heatid="5068" lane="6" entrytime="00:01:28.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="452" swimtime="00:02:44.32" resultid="3283" heatid="5189" lane="4" entrytime="00:02:47.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.01" />
                    <SPLIT distance="100" swimtime="00:01:18.45" />
                    <SPLIT distance="150" swimtime="00:02:05.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="408" swimtime="00:01:17.25" resultid="3284" heatid="5246" lane="3" entrytime="00:01:21.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" status="DNS" swimtime="00:00:00.00" resultid="3285" heatid="5280" lane="8" entrytime="00:06:00.38" entrycourse="LCM" />
                <RESULT eventid="1243" points="355" swimtime="00:03:14.20" resultid="3286" heatid="5312" lane="1" entrytime="00:03:15.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.38" />
                    <SPLIT distance="100" swimtime="00:01:31.69" />
                    <SPLIT distance="150" swimtime="00:02:21.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1275" points="386" swimtime="00:02:49.03" resultid="3287" heatid="5342" lane="1" entrytime="00:02:47.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.64" />
                    <SPLIT distance="100" swimtime="00:01:23.40" />
                    <SPLIT distance="150" swimtime="00:02:06.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Zital" birthdate="1991-05-03" gender="M" nation="BRA" license="093924" swrid="5727652" athleteid="3237" externalid="093924">
              <RESULTS>
                <RESULT eventid="1182" points="492" swimtime="00:01:05.32" resultid="3238" heatid="5262" lane="5" entrytime="00:01:07.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="477" swimtime="00:00:30.12" resultid="3239" heatid="5287" lane="6" entrytime="00:00:29.66" entrycourse="LCM" />
                <RESULT eventid="1277" points="443" swimtime="00:02:26.80" resultid="3240" heatid="5347" lane="2" entrytime="00:02:25.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.97" />
                    <SPLIT distance="100" swimtime="00:01:08.97" />
                    <SPLIT distance="150" swimtime="00:01:48.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Rinaldini" birthdate="2009-04-09" gender="M" nation="BRA" license="348289" swrid="5596932" athleteid="3267" externalid="348289">
              <RESULTS>
                <RESULT eventid="1072" points="577" swimtime="00:04:24.25" resultid="3268" heatid="5062" lane="6" entrytime="00:04:23.82" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.15" />
                    <SPLIT distance="100" swimtime="00:01:02.49" />
                    <SPLIT distance="150" swimtime="00:01:35.81" />
                    <SPLIT distance="200" swimtime="00:02:09.14" />
                    <SPLIT distance="250" swimtime="00:02:42.29" />
                    <SPLIT distance="300" swimtime="00:03:16.08" />
                    <SPLIT distance="350" swimtime="00:03:50.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="497" swimtime="00:01:02.40" resultid="3269" heatid="5174" lane="2" entrytime="00:01:03.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="534" swimtime="00:04:58.89" resultid="3270" heatid="5277" lane="6" entrytime="00:05:04.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.53" />
                    <SPLIT distance="100" swimtime="00:01:05.43" />
                    <SPLIT distance="150" swimtime="00:01:46.44" />
                    <SPLIT distance="200" swimtime="00:02:26.05" />
                    <SPLIT distance="250" swimtime="00:03:09.42" />
                    <SPLIT distance="300" swimtime="00:03:52.88" />
                    <SPLIT distance="350" swimtime="00:04:25.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="575" swimtime="00:09:03.53" resultid="3271" heatid="5300" lane="3" entrytime="00:09:08.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.90" />
                    <SPLIT distance="100" swimtime="00:01:04.24" />
                    <SPLIT distance="150" swimtime="00:01:38.16" />
                    <SPLIT distance="200" swimtime="00:02:12.35" />
                    <SPLIT distance="250" swimtime="00:02:47.13" />
                    <SPLIT distance="300" swimtime="00:03:21.89" />
                    <SPLIT distance="350" swimtime="00:03:56.93" />
                    <SPLIT distance="400" swimtime="00:04:31.48" />
                    <SPLIT distance="450" swimtime="00:05:05.87" />
                    <SPLIT distance="500" swimtime="00:05:40.17" />
                    <SPLIT distance="550" swimtime="00:06:14.97" />
                    <SPLIT distance="600" swimtime="00:06:49.11" />
                    <SPLIT distance="650" swimtime="00:07:23.25" />
                    <SPLIT distance="700" swimtime="00:07:57.72" />
                    <SPLIT distance="750" swimtime="00:08:31.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="439" swimtime="00:00:29.28" resultid="3272" heatid="5334" lane="7" entrytime="00:00:29.57" entrycourse="LCM" />
                <RESULT eventid="1293" points="520" swimtime="00:02:17.20" resultid="3273" heatid="5360" lane="6" entrytime="00:02:16.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.70" />
                    <SPLIT distance="100" swimtime="00:01:05.24" />
                    <SPLIT distance="150" swimtime="00:01:41.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Borille Busetti" birthdate="2010-02-17" gender="F" nation="BRA" license="392830" swrid="5622263" athleteid="3428" externalid="392830">
              <RESULTS>
                <RESULT eventid="1096" points="422" swimtime="00:00:31.47" resultid="3429" heatid="5095" lane="4" />
                <RESULT eventid="1112" points="403" swimtime="00:02:32.70" resultid="3430" heatid="5139" lane="2" entrytime="00:02:33.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.16" />
                    <SPLIT distance="100" swimtime="00:01:14.74" />
                    <SPLIT distance="150" swimtime="00:01:54.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="294" swimtime="00:01:26.14" resultid="3431" heatid="5242" lane="4" entrytime="00:01:23.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="424" swimtime="00:01:08.78" resultid="3432" heatid="5203" lane="4" entrytime="00:01:09.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="347" swimtime="00:00:38.22" resultid="3433" heatid="5292" lane="5" entrytime="00:00:41.38" entrycourse="LCM" />
                <RESULT eventid="1275" points="293" swimtime="00:03:05.20" resultid="3434" heatid="5340" lane="2" entrytime="00:03:03.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.26" />
                    <SPLIT distance="100" swimtime="00:01:29.64" />
                    <SPLIT distance="150" swimtime="00:02:17.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Luisa Lottermann" birthdate="2011-08-26" gender="F" nation="BRA" license="382238" swrid="5596909" athleteid="3372" externalid="382238">
              <RESULTS>
                <RESULT eventid="1080" points="370" swimtime="00:01:29.28" resultid="3373" heatid="5066" lane="5" entrytime="00:01:28.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" points="237" swimtime="00:01:29.61" resultid="3374" heatid="5159" lane="6" entrytime="00:01:38.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="294" swimtime="00:03:09.66" resultid="3375" heatid="5187" lane="7" entrytime="00:03:02.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.77" />
                    <SPLIT distance="100" swimtime="00:01:38.34" />
                    <SPLIT distance="150" swimtime="00:02:26.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="355" swimtime="00:06:15.45" resultid="3376" heatid="5279" lane="3" entrytime="00:06:10.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.97" />
                    <SPLIT distance="100" swimtime="00:01:32.26" />
                    <SPLIT distance="150" swimtime="00:02:24.12" />
                    <SPLIT distance="200" swimtime="00:03:16.75" />
                    <SPLIT distance="250" swimtime="00:04:04.18" />
                    <SPLIT distance="300" swimtime="00:04:52.25" />
                    <SPLIT distance="350" swimtime="00:05:34.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="402" swimtime="00:03:06.31" resultid="3377" heatid="5313" lane="8" entrytime="00:03:04.15" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.63" />
                    <SPLIT distance="100" swimtime="00:01:30.50" />
                    <SPLIT distance="150" swimtime="00:02:18.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1295" points="247" swimtime="00:03:14.08" resultid="3378" heatid="5361" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.71" />
                    <SPLIT distance="100" swimtime="00:01:33.31" />
                    <SPLIT distance="150" swimtime="00:02:24.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Colaco Da Conceicao" birthdate="2011-05-25" gender="F" nation="BRA" license="369535" swrid="5588601" athleteid="3337" externalid="369535">
              <RESULTS>
                <RESULT eventid="1064" points="454" swimtime="00:05:06.17" resultid="3338" heatid="5050" lane="4" entrytime="00:05:07.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.94" />
                    <SPLIT distance="100" swimtime="00:01:11.87" />
                    <SPLIT distance="150" swimtime="00:01:51.56" />
                    <SPLIT distance="200" swimtime="00:02:30.82" />
                    <SPLIT distance="250" swimtime="00:03:10.47" />
                    <SPLIT distance="300" swimtime="00:03:49.93" />
                    <SPLIT distance="350" swimtime="00:04:29.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="425" swimtime="00:02:30.05" resultid="3339" heatid="5139" lane="5" entrytime="00:02:31.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.88" />
                    <SPLIT distance="100" swimtime="00:01:12.06" />
                    <SPLIT distance="150" swimtime="00:01:51.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="427" swimtime="00:10:43.71" resultid="3340" heatid="5271" lane="5" entrytime="00:10:24.10" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:13.41" />
                    <SPLIT distance="150" swimtime="00:01:53.29" />
                    <SPLIT distance="200" swimtime="00:02:33.54" />
                    <SPLIT distance="250" swimtime="00:03:14.39" />
                    <SPLIT distance="300" swimtime="00:03:54.72" />
                    <SPLIT distance="350" swimtime="00:04:36.16" />
                    <SPLIT distance="400" swimtime="00:05:17.41" />
                    <SPLIT distance="450" swimtime="00:05:58.40" />
                    <SPLIT distance="500" swimtime="00:06:39.75" />
                    <SPLIT distance="550" swimtime="00:07:21.41" />
                    <SPLIT distance="600" swimtime="00:08:02.47" />
                    <SPLIT distance="650" swimtime="00:08:43.41" />
                    <SPLIT distance="700" swimtime="00:09:25.18" />
                    <SPLIT distance="750" swimtime="00:10:05.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="320" swimtime="00:00:39.23" resultid="3341" heatid="5292" lane="7" entrytime="00:00:43.45" entrycourse="LCM" />
                <RESULT eventid="1279" points="423" swimtime="00:20:25.82" resultid="3342" heatid="5350" lane="6" entrytime="00:20:00.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:13.33" />
                    <SPLIT distance="150" swimtime="00:01:54.15" />
                    <SPLIT distance="200" swimtime="00:02:34.33" />
                    <SPLIT distance="250" swimtime="00:03:15.26" />
                    <SPLIT distance="300" swimtime="00:03:56.25" />
                    <SPLIT distance="350" swimtime="00:04:37.92" />
                    <SPLIT distance="400" swimtime="00:05:19.76" />
                    <SPLIT distance="450" swimtime="00:06:00.89" />
                    <SPLIT distance="500" swimtime="00:06:42.31" />
                    <SPLIT distance="550" swimtime="00:07:24.01" />
                    <SPLIT distance="600" swimtime="00:08:05.16" />
                    <SPLIT distance="650" swimtime="00:08:46.71" />
                    <SPLIT distance="700" swimtime="00:09:27.63" />
                    <SPLIT distance="750" swimtime="00:10:09.33" />
                    <SPLIT distance="800" swimtime="00:10:50.59" />
                    <SPLIT distance="850" swimtime="00:11:32.06" />
                    <SPLIT distance="900" swimtime="00:12:13.67" />
                    <SPLIT distance="950" swimtime="00:12:55.00" />
                    <SPLIT distance="1000" swimtime="00:13:36.47" />
                    <SPLIT distance="1050" swimtime="00:14:18.60" />
                    <SPLIT distance="1100" swimtime="00:15:00.11" />
                    <SPLIT distance="1150" swimtime="00:15:42.22" />
                    <SPLIT distance="1200" swimtime="00:16:23.87" />
                    <SPLIT distance="1250" swimtime="00:17:05.36" />
                    <SPLIT distance="1300" swimtime="00:17:46.16" />
                    <SPLIT distance="1350" swimtime="00:18:27.01" />
                    <SPLIT distance="1400" swimtime="00:19:07.69" />
                    <SPLIT distance="1450" swimtime="00:19:47.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1295" points="286" swimtime="00:03:04.72" resultid="3343" heatid="5361" lane="4" entrytime="00:03:06.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.00" />
                    <SPLIT distance="100" swimtime="00:01:26.86" />
                    <SPLIT distance="150" swimtime="00:02:17.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Bertelli Weirich" birthdate="2011-03-18" gender="F" nation="BRA" license="369534" swrid="5588552" athleteid="3330" externalid="369534">
              <RESULTS>
                <RESULT eventid="1064" points="455" swimtime="00:05:05.99" resultid="3331" heatid="5050" lane="3" entrytime="00:05:08.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.79" />
                    <SPLIT distance="150" swimtime="00:01:51.49" />
                    <SPLIT distance="250" swimtime="00:03:10.48" />
                    <SPLIT distance="350" swimtime="00:04:29.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" points="409" swimtime="00:01:14.73" resultid="3332" heatid="5160" lane="7" entrytime="00:01:20.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="448" swimtime="00:02:44.79" resultid="3333" heatid="5188" lane="3" entrytime="00:02:44.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.13" />
                    <SPLIT distance="100" swimtime="00:01:18.92" />
                    <SPLIT distance="150" swimtime="00:02:08.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="402" swimtime="00:01:17.62" resultid="3334" heatid="5242" lane="5" entrytime="00:01:23.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="430" swimtime="00:05:52.02" resultid="3335" heatid="5280" lane="1" entrytime="00:05:52.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.71" />
                    <SPLIT distance="100" swimtime="00:01:21.15" />
                    <SPLIT distance="150" swimtime="00:02:05.90" />
                    <SPLIT distance="200" swimtime="00:02:51.00" />
                    <SPLIT distance="250" swimtime="00:03:42.36" />
                    <SPLIT distance="300" swimtime="00:04:34.72" />
                    <SPLIT distance="350" swimtime="00:05:13.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1295" points="395" swimtime="00:02:45.89" resultid="3336" heatid="5362" lane="1" entrytime="00:03:01.13" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.53" />
                    <SPLIT distance="100" swimtime="00:01:19.52" />
                    <SPLIT distance="150" swimtime="00:02:02.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2328" points="385" swimtime="00:01:16.24" resultid="6004" heatid="6418" lane="8" entrytime="00:01:14.73">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Zimmermann" birthdate="2010-01-19" gender="M" nation="BRA" license="357160" swrid="5588977" athleteid="3288" externalid="357160">
              <RESULTS>
                <RESULT eventid="1072" points="525" swimtime="00:04:32.73" resultid="3289" heatid="5059" lane="6" entrytime="00:04:38.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.95" />
                    <SPLIT distance="100" swimtime="00:01:03.39" />
                    <SPLIT distance="150" swimtime="00:01:38.40" />
                    <SPLIT distance="200" swimtime="00:02:13.20" />
                    <SPLIT distance="250" swimtime="00:02:48.40" />
                    <SPLIT distance="300" swimtime="00:03:23.88" />
                    <SPLIT distance="350" swimtime="00:03:58.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="519" swimtime="00:02:06.85" resultid="3290" heatid="5152" lane="8" entrytime="00:02:12.96" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.95" />
                    <SPLIT distance="100" swimtime="00:01:01.05" />
                    <SPLIT distance="150" swimtime="00:01:34.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="523" swimtime="00:02:21.49" resultid="3291" heatid="5195" lane="5" entrytime="00:02:24.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.39" />
                    <SPLIT distance="100" swimtime="00:01:07.67" />
                    <SPLIT distance="150" swimtime="00:01:50.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="461" swimtime="00:01:06.76" resultid="3292" heatid="5258" lane="6" entrytime="00:01:06.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="497" swimtime="00:09:30.40" resultid="3293" heatid="5299" lane="3" entrytime="00:09:41.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:06.27" />
                    <SPLIT distance="150" swimtime="00:01:41.93" />
                    <SPLIT distance="200" swimtime="00:02:17.59" />
                    <SPLIT distance="250" swimtime="00:02:52.41" />
                    <SPLIT distance="300" swimtime="00:03:28.13" />
                    <SPLIT distance="350" swimtime="00:04:04.80" />
                    <SPLIT distance="400" swimtime="00:04:41.67" />
                    <SPLIT distance="450" swimtime="00:05:17.79" />
                    <SPLIT distance="500" swimtime="00:05:54.44" />
                    <SPLIT distance="550" swimtime="00:06:29.65" />
                    <SPLIT distance="600" swimtime="00:07:06.15" />
                    <SPLIT distance="650" swimtime="00:07:43.40" />
                    <SPLIT distance="700" swimtime="00:08:20.44" />
                    <SPLIT distance="750" swimtime="00:08:54.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="474" swimtime="00:02:23.50" resultid="3294" heatid="5348" lane="8" entrytime="00:02:22.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.51" />
                    <SPLIT distance="100" swimtime="00:01:09.47" />
                    <SPLIT distance="150" swimtime="00:01:47.32" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luann" lastname="Miguel Mazur" birthdate="2007-01-10" gender="M" nation="BRA" license="365682" swrid="5596915" athleteid="3302" externalid="365682">
              <RESULTS>
                <RESULT eventid="1088" points="448" swimtime="00:01:14.29" resultid="3303" heatid="5087" lane="8" entrytime="00:01:15.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="471" swimtime="00:02:26.49" resultid="3304" heatid="5200" lane="3" entrytime="00:02:25.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.57" />
                    <SPLIT distance="100" swimtime="00:01:10.04" />
                    <SPLIT distance="150" swimtime="00:01:53.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="376" swimtime="00:01:11.43" resultid="3305" heatid="5262" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="451" swimtime="00:05:16.15" resultid="3306" heatid="5277" lane="2" entrytime="00:05:07.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.34" />
                    <SPLIT distance="100" swimtime="00:01:09.79" />
                    <SPLIT distance="150" swimtime="00:01:51.25" />
                    <SPLIT distance="200" swimtime="00:02:32.06" />
                    <SPLIT distance="250" swimtime="00:03:17.12" />
                    <SPLIT distance="300" swimtime="00:04:01.96" />
                    <SPLIT distance="350" swimtime="00:04:38.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="432" swimtime="00:02:45.98" resultid="3307" heatid="5319" lane="5" entrytime="00:02:39.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.22" />
                    <SPLIT distance="100" swimtime="00:01:20.52" />
                    <SPLIT distance="150" swimtime="00:02:03.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="399" swimtime="00:00:35.24" resultid="3308" heatid="5369" lane="4" entrytime="00:00:34.21" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Claudio" lastname="Rohnelt" birthdate="2010-03-08" gender="M" nation="BRA" license="357954" swrid="5596935" athleteid="3295" externalid="357954">
              <RESULTS>
                <RESULT eventid="1072" points="355" swimtime="00:05:10.80" resultid="3296" heatid="5057" lane="5" entrytime="00:05:12.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                    <SPLIT distance="100" swimtime="00:01:11.21" />
                    <SPLIT distance="150" swimtime="00:01:50.17" />
                    <SPLIT distance="200" swimtime="00:02:29.74" />
                    <SPLIT distance="250" swimtime="00:03:10.04" />
                    <SPLIT distance="300" swimtime="00:03:50.60" />
                    <SPLIT distance="350" swimtime="00:04:30.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="323" swimtime="00:01:12.06" resultid="3297" heatid="5171" lane="8" entrytime="00:01:13.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="404" swimtime="00:02:17.94" resultid="3298" heatid="5150" lane="5" entrytime="00:02:26.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                    <SPLIT distance="100" swimtime="00:01:05.92" />
                    <SPLIT distance="150" swimtime="00:01:41.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="391" swimtime="00:01:04.08" resultid="3299" heatid="5221" lane="1" entrytime="00:01:06.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="340" swimtime="00:00:31.90" resultid="3300" heatid="5328" lane="7" />
                <RESULT eventid="1293" points="316" swimtime="00:02:41.89" resultid="3301" heatid="5358" lane="2" entrytime="00:02:50.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.88" />
                    <SPLIT distance="100" swimtime="00:01:16.44" />
                    <SPLIT distance="150" swimtime="00:01:59.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Vitoria Gugel" birthdate="2011-12-08" gender="F" nation="BRA" license="365490" swrid="5588960" athleteid="3421" externalid="365490">
              <RESULTS>
                <RESULT eventid="1080" points="339" swimtime="00:01:31.95" resultid="3422" heatid="5065" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" points="284" swimtime="00:01:24.33" resultid="3423" heatid="5160" lane="1" entrytime="00:01:24.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="384" swimtime="00:06:05.77" resultid="3424" heatid="5279" lane="5" entrytime="00:06:06.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.29" />
                    <SPLIT distance="100" swimtime="00:01:23.18" />
                    <SPLIT distance="150" swimtime="00:02:11.68" />
                    <SPLIT distance="200" swimtime="00:02:58.08" />
                    <SPLIT distance="250" swimtime="00:03:48.30" />
                    <SPLIT distance="300" swimtime="00:04:38.94" />
                    <SPLIT distance="350" swimtime="00:05:23.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="288" swimtime="00:00:36.96" resultid="3425" heatid="5324" lane="7" entrytime="00:00:37.21" entrycourse="LCM" />
                <RESULT eventid="1243" points="347" swimtime="00:03:15.68" resultid="3426" heatid="5311" lane="4" entrytime="00:03:16.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.42" />
                    <SPLIT distance="100" swimtime="00:01:34.07" />
                    <SPLIT distance="150" swimtime="00:02:25.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1295" points="284" swimtime="00:03:05.11" resultid="3427" heatid="5362" lane="8" entrytime="00:03:04.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.36" />
                    <SPLIT distance="100" swimtime="00:01:26.71" />
                    <SPLIT distance="150" swimtime="00:02:18.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Emanuel" lastname="Ranieri" birthdate="2011-01-24" gender="M" nation="BRA" license="390838" swrid="5596930" athleteid="3400" externalid="390838">
              <RESULTS>
                <RESULT eventid="1088" points="269" swimtime="00:01:28.05" resultid="3401" heatid="5080" lane="4" entrytime="00:01:29.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="351" swimtime="00:02:41.61" resultid="3402" heatid="5194" lane="2" entrytime="00:02:46.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.00" />
                    <SPLIT distance="100" swimtime="00:01:16.01" />
                    <SPLIT distance="150" swimtime="00:02:05.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="307" swimtime="00:01:16.47" resultid="3403" heatid="5256" lane="6" entrytime="00:01:20.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="356" swimtime="00:05:42.09" resultid="3404" heatid="5276" lane="7" entrytime="00:05:41.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.58" />
                    <SPLIT distance="150" swimtime="00:02:02.93" />
                    <SPLIT distance="250" swimtime="00:03:37.60" />
                    <SPLIT distance="350" swimtime="00:05:05.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="279" swimtime="00:03:11.83" resultid="3405" heatid="5317" lane="1" entrytime="00:03:11.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.85" />
                    <SPLIT distance="100" swimtime="00:01:32.67" />
                    <SPLIT distance="150" swimtime="00:02:22.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="298" swimtime="00:02:47.55" resultid="3406" heatid="5345" lane="7" entrytime="00:02:48.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.13" />
                    <SPLIT distance="100" swimtime="00:01:22.91" />
                    <SPLIT distance="150" swimtime="00:02:06.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Ramirez Vasconcelos" birthdate="2011-04-06" gender="M" nation="BRA" license="392013" swrid="4863662" athleteid="3414" externalid="392013">
              <RESULTS>
                <RESULT eventid="1088" points="322" swimtime="00:01:22.91" resultid="3415" heatid="5082" lane="1" entrytime="00:01:21.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="337" swimtime="00:02:43.81" resultid="3416" heatid="5194" lane="3" entrytime="00:02:44.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                    <SPLIT distance="100" swimtime="00:01:16.93" />
                    <SPLIT distance="150" swimtime="00:02:04.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="325" swimtime="00:05:52.49" resultid="3417" heatid="5276" lane="8" entrytime="00:05:53.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.63" />
                    <SPLIT distance="100" swimtime="00:01:18.56" />
                    <SPLIT distance="150" swimtime="00:02:06.33" />
                    <SPLIT distance="200" swimtime="00:02:53.51" />
                    <SPLIT distance="250" swimtime="00:03:42.66" />
                    <SPLIT distance="300" swimtime="00:04:32.87" />
                    <SPLIT distance="350" swimtime="00:05:13.25" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="312" swimtime="00:00:32.83" resultid="3418" heatid="5327" lane="3" />
                <RESULT eventid="1251" points="346" swimtime="00:02:58.60" resultid="3419" heatid="5317" lane="4" entrytime="00:02:58.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.10" />
                    <SPLIT distance="100" swimtime="00:01:24.49" />
                    <SPLIT distance="150" swimtime="00:02:11.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="316" swimtime="00:00:38.07" resultid="3420" heatid="5365" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Paiz Ribeiro" birthdate="2006-02-17" gender="M" nation="BRA" license="297583" swrid="5596921" athleteid="3241" externalid="297583">
              <RESULTS>
                <RESULT eventid="1088" points="385" swimtime="00:01:18.14" resultid="3242" heatid="5086" lane="5" entrytime="00:01:19.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1072" points="499" swimtime="00:04:37.30" resultid="3243" heatid="5063" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                    <SPLIT distance="100" swimtime="00:01:05.75" />
                    <SPLIT distance="150" swimtime="00:01:41.06" />
                    <SPLIT distance="200" swimtime="00:02:16.18" />
                    <SPLIT distance="250" swimtime="00:02:51.69" />
                    <SPLIT distance="300" swimtime="00:03:27.02" />
                    <SPLIT distance="350" swimtime="00:04:02.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="498" swimtime="00:01:02.38" resultid="3244" heatid="5177" lane="6" entrytime="00:01:02.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="483" swimtime="00:09:36.08" resultid="3245" heatid="5300" lane="1" entrytime="00:09:36.03" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                    <SPLIT distance="100" swimtime="00:01:06.71" />
                    <SPLIT distance="150" swimtime="00:01:42.50" />
                    <SPLIT distance="200" swimtime="00:02:18.75" />
                    <SPLIT distance="250" swimtime="00:02:55.12" />
                    <SPLIT distance="300" swimtime="00:03:31.73" />
                    <SPLIT distance="350" swimtime="00:04:07.82" />
                    <SPLIT distance="400" swimtime="00:04:44.29" />
                    <SPLIT distance="450" swimtime="00:05:20.84" />
                    <SPLIT distance="500" swimtime="00:05:57.76" />
                    <SPLIT distance="550" swimtime="00:06:34.07" />
                    <SPLIT distance="600" swimtime="00:07:11.13" />
                    <SPLIT distance="650" swimtime="00:07:47.54" />
                    <SPLIT distance="700" swimtime="00:08:24.31" />
                    <SPLIT distance="750" swimtime="00:09:00.71" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="483" swimtime="00:00:28.37" resultid="3246" heatid="5328" lane="6" />
                <RESULT eventid="1251" points="427" swimtime="00:02:46.60" resultid="3247" heatid="5319" lane="8" entrytime="00:02:44.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.07" />
                    <SPLIT distance="100" swimtime="00:01:18.89" />
                    <SPLIT distance="150" swimtime="00:02:02.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Danilo" lastname="Rodrigues" birthdate="2011-05-23" gender="M" nation="BRA" license="370763" swrid="5596934" athleteid="3344" externalid="370763">
              <RESULTS>
                <RESULT eventid="1088" points="303" swimtime="00:01:24.64" resultid="3345" heatid="5081" lane="1" entrytime="00:01:28.55" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="304" swimtime="00:01:13.48" resultid="3346" heatid="5171" lane="2" entrytime="00:01:10.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="316" swimtime="00:02:47.25" resultid="3347" heatid="5192" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.72" />
                    <SPLIT distance="150" swimtime="00:02:10.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="356" swimtime="00:05:42.01" resultid="3348" heatid="5276" lane="6" entrytime="00:05:39.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.05" />
                    <SPLIT distance="100" swimtime="00:01:16.31" />
                    <SPLIT distance="150" swimtime="00:02:03.92" />
                    <SPLIT distance="250" swimtime="00:03:38.49" />
                    <SPLIT distance="300" swimtime="00:04:27.60" />
                    <SPLIT distance="350" swimtime="00:05:04.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="333" swimtime="00:03:00.97" resultid="3349" heatid="5317" lane="5" entrytime="00:03:00.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.73" />
                    <SPLIT distance="100" swimtime="00:01:28.11" />
                    <SPLIT distance="150" swimtime="00:02:15.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1293" points="319" swimtime="00:02:41.39" resultid="3350" heatid="5359" lane="1" entrytime="00:02:37.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.75" />
                    <SPLIT distance="100" swimtime="00:01:17.53" />
                    <SPLIT distance="150" swimtime="00:01:59.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Balduíno" birthdate="2009-06-24" gender="M" nation="BRA" license="370764" swrid="5596870" athleteid="3351" externalid="370764">
              <RESULTS>
                <RESULT eventid="1135" points="531" swimtime="00:01:01.06" resultid="3352" heatid="5175" lane="8" entrytime="00:01:02.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="487" swimtime="00:02:24.81" resultid="3353" heatid="5197" lane="5" entrytime="00:02:27.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.12" />
                    <SPLIT distance="100" swimtime="00:01:08.30" />
                    <SPLIT distance="150" swimtime="00:01:51.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="439" swimtime="00:01:07.88" resultid="3354" heatid="5260" lane="5" entrytime="00:01:07.19" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="471" swimtime="00:05:11.61" resultid="3355" heatid="5277" lane="7" entrytime="00:05:07.87" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.45" />
                    <SPLIT distance="150" swimtime="00:01:47.64" />
                    <SPLIT distance="250" swimtime="00:03:13.83" />
                    <SPLIT distance="350" swimtime="00:04:38.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="458" swimtime="00:02:25.16" resultid="3356" heatid="5345" lane="4" entrytime="00:02:37.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.71" />
                    <SPLIT distance="100" swimtime="00:01:11.50" />
                    <SPLIT distance="150" swimtime="00:01:49.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1293" points="469" swimtime="00:02:21.92" resultid="3357" heatid="5360" lane="7" entrytime="00:02:21.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.17" />
                    <SPLIT distance="100" swimtime="00:01:07.42" />
                    <SPLIT distance="150" swimtime="00:01:45.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Stein Duarte" birthdate="2010-10-03" gender="F" nation="BRA" license="351635" swrid="5588923" athleteid="3274" externalid="351635">
              <RESULTS>
                <RESULT eventid="1064" points="385" swimtime="00:05:23.48" resultid="3275" heatid="5049" lane="6" entrytime="00:05:29.64" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.91" />
                    <SPLIT distance="100" swimtime="00:01:13.39" />
                    <SPLIT distance="150" swimtime="00:01:54.88" />
                    <SPLIT distance="200" swimtime="00:02:36.78" />
                    <SPLIT distance="250" swimtime="00:03:18.29" />
                    <SPLIT distance="300" swimtime="00:03:59.98" />
                    <SPLIT distance="350" swimtime="00:04:42.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="458" swimtime="00:02:43.54" resultid="3276" heatid="5188" lane="5" entrytime="00:02:39.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.24" />
                    <SPLIT distance="100" swimtime="00:01:17.97" />
                    <SPLIT distance="150" swimtime="00:02:07.07" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="489" swimtime="00:01:12.76" resultid="3277" heatid="5244" lane="4" entrytime="00:01:13.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1205" points="445" swimtime="00:05:48.07" resultid="3278" heatid="5280" lane="2" entrytime="00:05:41.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.14" />
                    <SPLIT distance="100" swimtime="00:01:20.12" />
                    <SPLIT distance="150" swimtime="00:02:03.00" />
                    <SPLIT distance="200" swimtime="00:02:44.97" />
                    <SPLIT distance="250" swimtime="00:03:36.37" />
                    <SPLIT distance="300" swimtime="00:04:26.52" />
                    <SPLIT distance="350" swimtime="00:05:07.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="461" swimtime="00:00:34.76" resultid="3279" heatid="5289" lane="3" />
                <RESULT eventid="1275" points="475" swimtime="00:02:37.81" resultid="3280" heatid="5343" lane="6" entrytime="00:02:35.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.80" />
                    <SPLIT distance="100" swimtime="00:01:16.97" />
                    <SPLIT distance="150" swimtime="00:01:58.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2391" points="446" swimtime="00:01:14.99" resultid="6134" heatid="6424" lane="1" entrytime="00:01:12.76">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Alves Serafini" birthdate="2008-04-15" gender="M" nation="BRA" license="351644" swrid="5596867" athleteid="3393" externalid="351644">
              <RESULTS>
                <RESULT eventid="1072" points="526" swimtime="00:04:32.47" resultid="3394" heatid="5061" lane="4" entrytime="00:04:36.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:02.20" />
                    <SPLIT distance="150" swimtime="00:01:35.07" />
                    <SPLIT distance="200" swimtime="00:02:08.71" />
                    <SPLIT distance="250" swimtime="00:02:43.11" />
                    <SPLIT distance="300" swimtime="00:03:17.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="530" swimtime="00:01:01.07" resultid="3395" heatid="5175" lane="6" entrytime="00:01:00.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="502" swimtime="00:00:58.93" resultid="3396" heatid="5228" lane="5" entrytime="00:00:58.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="448" swimtime="00:05:16.91" resultid="3397" heatid="5275" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.11" />
                    <SPLIT distance="150" swimtime="00:01:45.57" />
                    <SPLIT distance="250" swimtime="00:03:15.60" />
                    <SPLIT distance="350" swimtime="00:04:42.16" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="485" swimtime="00:00:28.33" resultid="3398" heatid="5335" lane="2" entrytime="00:00:28.26" entrycourse="LCM" />
                <RESULT eventid="1293" points="532" swimtime="00:02:16.13" resultid="3399" heatid="5360" lane="3" entrytime="00:02:15.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.61" />
                    <SPLIT distance="100" swimtime="00:01:03.11" />
                    <SPLIT distance="150" swimtime="00:01:39.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Souza Garute Da Silva" birthdate="2009-01-07" gender="F" nation="BRA" license="329307" swrid="5596940" athleteid="3262" externalid="329307">
              <RESULTS>
                <RESULT eventid="1175" points="400" swimtime="00:01:17.79" resultid="3263" heatid="5247" lane="2" entrytime="00:01:13.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="415" swimtime="00:00:36.01" resultid="3264" heatid="5290" lane="8" />
                <RESULT eventid="1275" points="404" swimtime="00:02:46.45" resultid="3265" heatid="5343" lane="7" entrytime="00:02:39.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.58" />
                    <SPLIT distance="100" swimtime="00:01:20.34" />
                    <SPLIT distance="150" swimtime="00:02:04.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="355" swimtime="00:00:41.17" resultid="3266" heatid="5373" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Mariotti De Castro" birthdate="2008-06-27" gender="M" nation="BRA" license="329200" swrid="5596912" athleteid="3255" externalid="329200">
              <RESULTS>
                <RESULT eventid="1072" points="625" swimtime="00:04:17.28" resultid="3256" heatid="5062" lane="4" entrytime="00:04:12.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.70" />
                    <SPLIT distance="100" swimtime="00:01:00.01" />
                    <SPLIT distance="200" swimtime="00:02:06.33" />
                    <SPLIT distance="250" swimtime="00:02:39.43" />
                    <SPLIT distance="300" swimtime="00:03:12.11" />
                    <SPLIT distance="350" swimtime="00:03:44.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="616" swimtime="00:01:59.87" resultid="3257" heatid="5156" lane="6" entrytime="00:02:02.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.92" />
                    <SPLIT distance="100" swimtime="00:00:58.13" />
                    <SPLIT distance="150" swimtime="00:01:28.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="508" swimtime="00:02:22.80" resultid="3258" heatid="5198" lane="5" entrytime="00:02:15.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.46" />
                    <SPLIT distance="100" swimtime="00:01:04.82" />
                    <SPLIT distance="150" swimtime="00:01:50.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="578" swimtime="00:00:56.23" resultid="3259" heatid="5228" lane="4" entrytime="00:00:57.78" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="433" swimtime="00:00:31.11" resultid="3260" heatid="5281" lane="3" />
                <RESULT eventid="1277" points="520" swimtime="00:02:19.12" resultid="3261" heatid="5344" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:09.15" />
                    <SPLIT distance="150" swimtime="00:01:44.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Flavia" lastname="De Metz" birthdate="2011-01-07" gender="F" nation="BRA" license="390846" swrid="5596887" athleteid="3407" externalid="390846">
              <RESULTS>
                <RESULT eventid="1064" points="393" swimtime="00:05:21.27" resultid="3408" heatid="5050" lane="7" entrytime="00:05:11.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.74" />
                    <SPLIT distance="100" swimtime="00:01:13.77" />
                    <SPLIT distance="150" swimtime="00:01:54.50" />
                    <SPLIT distance="200" swimtime="00:02:35.35" />
                    <SPLIT distance="250" swimtime="00:03:16.56" />
                    <SPLIT distance="300" swimtime="00:03:59.07" />
                    <SPLIT distance="350" swimtime="00:04:40.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="434" swimtime="00:02:29.05" resultid="3409" heatid="5141" lane="8" entrytime="00:02:24.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                    <SPLIT distance="100" swimtime="00:01:10.25" />
                    <SPLIT distance="150" swimtime="00:01:48.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="441" swimtime="00:01:07.90" resultid="3410" heatid="5204" lane="5" entrytime="00:01:06.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="385" swimtime="00:11:05.84" resultid="3411" heatid="5271" lane="7" entrytime="00:10:45.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.93" />
                    <SPLIT distance="100" swimtime="00:01:15.48" />
                    <SPLIT distance="150" swimtime="00:01:57.16" />
                    <SPLIT distance="200" swimtime="00:02:39.93" />
                    <SPLIT distance="250" swimtime="00:03:23.47" />
                    <SPLIT distance="300" swimtime="00:04:07.27" />
                    <SPLIT distance="350" swimtime="00:04:49.77" />
                    <SPLIT distance="400" swimtime="00:05:32.36" />
                    <SPLIT distance="450" swimtime="00:06:15.57" />
                    <SPLIT distance="500" swimtime="00:06:58.40" />
                    <SPLIT distance="550" swimtime="00:07:41.06" />
                    <SPLIT distance="600" swimtime="00:08:22.97" />
                    <SPLIT distance="650" swimtime="00:09:04.60" />
                    <SPLIT distance="700" swimtime="00:09:46.75" />
                    <SPLIT distance="750" swimtime="00:10:27.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="353" swimtime="00:00:37.97" resultid="3412" heatid="5289" lane="2" />
                <RESULT eventid="1275" points="361" swimtime="00:02:52.82" resultid="3413" heatid="5341" lane="2" entrytime="00:02:52.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.75" />
                    <SPLIT distance="100" swimtime="00:01:24.58" />
                    <SPLIT distance="150" swimtime="00:02:09.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Breno" lastname="Zanella Janke" birthdate="2011-04-26" gender="M" nation="BRA" license="365697" swrid="5588970" athleteid="3323" externalid="365697">
              <RESULTS>
                <RESULT eventid="1072" points="440" swimtime="00:04:49.33" resultid="3324" heatid="5059" lane="1" entrytime="00:04:48.92" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.29" />
                    <SPLIT distance="100" swimtime="00:01:07.64" />
                    <SPLIT distance="150" swimtime="00:01:44.10" />
                    <SPLIT distance="200" swimtime="00:02:20.78" />
                    <SPLIT distance="250" swimtime="00:02:56.80" />
                    <SPLIT distance="300" swimtime="00:03:33.93" />
                    <SPLIT distance="350" swimtime="00:04:11.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="414" swimtime="00:02:32.91" resultid="3325" heatid="5195" lane="3" entrytime="00:02:30.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="100" swimtime="00:01:13.62" />
                    <SPLIT distance="150" swimtime="00:01:58.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="386" swimtime="00:01:04.34" resultid="3326" heatid="5222" lane="2" entrytime="00:01:01.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="420" swimtime="00:10:03.36" resultid="3327" heatid="5297" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.54" />
                    <SPLIT distance="100" swimtime="00:01:12.03" />
                    <SPLIT distance="150" swimtime="00:01:49.78" />
                    <SPLIT distance="200" swimtime="00:02:27.16" />
                    <SPLIT distance="250" swimtime="00:03:05.08" />
                    <SPLIT distance="300" swimtime="00:03:43.11" />
                    <SPLIT distance="350" swimtime="00:04:21.59" />
                    <SPLIT distance="400" swimtime="00:04:59.87" />
                    <SPLIT distance="450" swimtime="00:05:38.36" />
                    <SPLIT distance="500" swimtime="00:06:16.51" />
                    <SPLIT distance="550" swimtime="00:06:55.13" />
                    <SPLIT distance="600" swimtime="00:07:33.69" />
                    <SPLIT distance="650" swimtime="00:08:12.04" />
                    <SPLIT distance="700" swimtime="00:08:50.34" />
                    <SPLIT distance="750" swimtime="00:09:28.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="366" swimtime="00:02:36.41" resultid="3328" heatid="5344" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                    <SPLIT distance="100" swimtime="00:01:16.45" />
                    <SPLIT distance="150" swimtime="00:01:56.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="372" swimtime="00:00:36.08" resultid="3329" heatid="5365" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1237" points="512" swimtime="00:03:55.20" resultid="3447" heatid="5308" lane="5" entrytime="00:03:57.40">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.09" />
                    <SPLIT distance="100" swimtime="00:00:58.43" />
                    <SPLIT distance="150" swimtime="00:01:26.71" />
                    <SPLIT distance="200" swimtime="00:01:57.50" />
                    <SPLIT distance="250" swimtime="00:02:26.58" />
                    <SPLIT distance="300" swimtime="00:02:57.72" />
                    <SPLIT distance="350" swimtime="00:03:25.41" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3393" number="1" />
                    <RELAYPOSITION athleteid="3351" number="2" />
                    <RELAYPOSITION athleteid="3358" number="3" />
                    <RELAYPOSITION athleteid="3255" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1338" points="493" swimtime="00:04:21.73" resultid="3452" heatid="5388" lane="5" entrytime="00:04:23.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.72" />
                    <SPLIT distance="150" swimtime="00:01:43.83" />
                    <SPLIT distance="200" swimtime="00:02:24.77" />
                    <SPLIT distance="250" swimtime="00:02:53.97" />
                    <SPLIT distance="300" swimtime="00:03:25.70" />
                    <SPLIT distance="350" swimtime="00:03:52.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3351" number="1" />
                    <RELAYPOSITION athleteid="3358" number="2" />
                    <RELAYPOSITION athleteid="3393" number="3" />
                    <RELAYPOSITION athleteid="3255" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1233" points="416" swimtime="00:04:12.10" resultid="3448" heatid="5306" lane="2" entrytime="00:04:24.41">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.44" />
                    <SPLIT distance="100" swimtime="00:01:01.37" />
                    <SPLIT distance="150" swimtime="00:01:29.85" />
                    <SPLIT distance="200" swimtime="00:02:01.28" />
                    <SPLIT distance="250" swimtime="00:02:31.56" />
                    <SPLIT distance="300" swimtime="00:03:05.69" />
                    <SPLIT distance="350" swimtime="00:03:36.77" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3386" number="1" />
                    <RELAYPOSITION athleteid="3288" number="2" />
                    <RELAYPOSITION athleteid="3295" number="3" />
                    <RELAYPOSITION athleteid="3435" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="SW 8.4 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 19:07), Na volta dos 250m (Revezamento Medley, Borboleta)." eventid="1334" status="DSQ" swimtime="00:04:44.89" resultid="3451" heatid="5386" lane="3" entrytime="00:04:39.35">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.64" />
                    <SPLIT distance="100" swimtime="00:01:10.46" />
                    <SPLIT distance="150" swimtime="00:01:47.17" />
                    <SPLIT distance="200" swimtime="00:02:28.46" />
                    <SPLIT distance="250" swimtime="00:03:00.16" />
                    <SPLIT distance="300" swimtime="00:03:38.74" />
                    <SPLIT distance="350" swimtime="00:04:10.47" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3386" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="3288" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="3295" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="3435" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1231" points="406" swimtime="00:04:14.13" resultid="3449" heatid="5305" lane="3" entrytime="00:04:17.63">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.49" />
                    <SPLIT distance="100" swimtime="00:01:02.65" />
                    <SPLIT distance="150" swimtime="00:01:31.45" />
                    <SPLIT distance="200" swimtime="00:02:03.33" />
                    <SPLIT distance="250" swimtime="00:02:33.78" />
                    <SPLIT distance="300" swimtime="00:03:07.00" />
                    <SPLIT distance="350" swimtime="00:03:38.46" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3323" number="1" />
                    <RELAYPOSITION athleteid="3309" number="2" />
                    <RELAYPOSITION athleteid="3400" number="3" />
                    <RELAYPOSITION athleteid="3344" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT comment="SW 10.12 - Os pés perderam contato com a plataforma de partida antes que o colega de equipe anterior tocasse a borda.  (Horário: 18:59)" eventid="1332" status="DSQ" swimtime="00:04:44.96" resultid="3450" heatid="5385" lane="4" entrytime="00:04:48.04">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.44" />
                    <SPLIT distance="100" swimtime="00:01:09.39" />
                    <SPLIT distance="150" swimtime="00:01:45.94" />
                    <SPLIT distance="200" swimtime="00:02:29.32" />
                    <SPLIT distance="250" swimtime="00:03:01.60" />
                    <SPLIT distance="300" swimtime="00:03:39.49" />
                    <SPLIT distance="350" swimtime="00:04:10.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3309" number="1" status="DSQ" />
                    <RELAYPOSITION athleteid="3414" number="2" status="DSQ" />
                    <RELAYPOSITION athleteid="3344" number="3" status="DSQ" />
                    <RELAYPOSITION athleteid="3400" number="4" status="DSQ" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="F" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1221" points="455" swimtime="00:04:30.28" resultid="3443" heatid="5302" lane="2" entrytime="00:04:42.25">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                    <SPLIT distance="100" swimtime="00:01:08.52" />
                    <SPLIT distance="150" swimtime="00:01:39.77" />
                    <SPLIT distance="200" swimtime="00:02:14.77" />
                    <SPLIT distance="250" swimtime="00:02:46.81" />
                    <SPLIT distance="300" swimtime="00:03:22.79" />
                    <SPLIT distance="350" swimtime="00:03:55.38" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3428" number="1" />
                    <RELAYPOSITION athleteid="3379" number="2" />
                    <RELAYPOSITION athleteid="3274" number="3" />
                    <RELAYPOSITION athleteid="3407" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1322" points="438" swimtime="00:05:03.35" resultid="3445" heatid="5382" lane="6" entrytime="00:05:18.24">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.04" />
                    <SPLIT distance="100" swimtime="00:01:16.58" />
                    <SPLIT distance="150" swimtime="00:01:54.93" />
                    <SPLIT distance="200" swimtime="00:02:40.33" />
                    <SPLIT distance="250" swimtime="00:03:14.70" />
                    <SPLIT distance="300" swimtime="00:03:55.87" />
                    <SPLIT distance="350" swimtime="00:04:28.05" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3274" number="1" />
                    <RELAYPOSITION athleteid="3379" number="2" />
                    <RELAYPOSITION athleteid="3330" number="3" />
                    <RELAYPOSITION athleteid="3428" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="F" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1219" points="359" swimtime="00:04:52.44" resultid="3444" heatid="5301" lane="3" entrytime="00:04:55.64">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.06" />
                    <SPLIT distance="100" swimtime="00:01:15.84" />
                    <SPLIT distance="150" swimtime="00:01:47.51" />
                    <SPLIT distance="200" swimtime="00:02:22.96" />
                    <SPLIT distance="250" swimtime="00:02:55.99" />
                    <SPLIT distance="300" swimtime="00:03:32.67" />
                    <SPLIT distance="350" swimtime="00:04:10.32" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3421" number="1" />
                    <RELAYPOSITION athleteid="3330" number="2" />
                    <RELAYPOSITION athleteid="3337" number="3" />
                    <RELAYPOSITION athleteid="3372" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1320" points="346" swimtime="00:05:28.02" resultid="3446" heatid="5381" lane="3" entrytime="00:05:28.88">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.74" />
                    <SPLIT distance="100" swimtime="00:01:22.89" />
                    <SPLIT distance="150" swimtime="00:02:05.75" />
                    <SPLIT distance="200" swimtime="00:02:53.97" />
                    <SPLIT distance="250" swimtime="00:03:32.13" />
                    <SPLIT distance="300" swimtime="00:04:16.53" />
                    <SPLIT distance="350" swimtime="00:04:50.52" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3407" number="1" />
                    <RELAYPOSITION athleteid="3372" number="2" />
                    <RELAYPOSITION athleteid="3421" number="3" />
                    <RELAYPOSITION athleteid="3337" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="15" agemin="15" agetotalmax="-1" agetotalmin="-1" gender="X" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1285" points="437" swimtime="00:04:46.62" resultid="3453" heatid="5353" lane="5" entrytime="00:04:32.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.54" />
                    <SPLIT distance="100" swimtime="00:01:16.65" />
                    <SPLIT distance="150" swimtime="00:01:57.85" />
                    <SPLIT distance="200" swimtime="00:02:45.21" />
                    <SPLIT distance="250" swimtime="00:03:15.22" />
                    <SPLIT distance="300" swimtime="00:03:48.93" />
                    <SPLIT distance="350" swimtime="00:04:16.56" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3262" number="1" />
                    <RELAYPOSITION athleteid="3281" number="2" />
                    <RELAYPOSITION athleteid="3267" number="3" />
                    <RELAYPOSITION athleteid="3351" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1283" points="416" swimtime="00:04:51.44" resultid="3454" heatid="5352" lane="2" entrytime="00:04:53.53">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.06" />
                    <SPLIT distance="100" swimtime="00:01:17.50" />
                    <SPLIT distance="150" swimtime="00:01:54.74" />
                    <SPLIT distance="200" swimtime="00:02:40.76" />
                    <SPLIT distance="250" swimtime="00:03:13.19" />
                    <SPLIT distance="300" swimtime="00:03:50.70" />
                    <SPLIT distance="350" swimtime="00:04:19.33" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3274" number="1" />
                    <RELAYPOSITION athleteid="3379" number="2" />
                    <RELAYPOSITION athleteid="3288" number="3" />
                    <RELAYPOSITION athleteid="3386" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="COMERCIAL CASCAVEL &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1281" points="392" swimtime="00:04:57.09" resultid="3455" heatid="5351" lane="3" entrytime="00:05:04.16">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.44" />
                    <SPLIT distance="100" swimtime="00:01:21.25" />
                    <SPLIT distance="150" swimtime="00:02:00.10" />
                    <SPLIT distance="200" swimtime="00:02:42.96" />
                    <SPLIT distance="250" swimtime="00:03:13.22" />
                    <SPLIT distance="300" swimtime="00:03:50.69" />
                    <SPLIT distance="350" swimtime="00:04:21.96" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3407" number="1" />
                    <RELAYPOSITION athleteid="3323" number="2" />
                    <RELAYPOSITION athleteid="3309" number="3" />
                    <RELAYPOSITION athleteid="3330" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="X" name="COMERCIAL CASCAVEL &quot;B&quot;" number="2">
              <RESULTS>
                <RESULT eventid="1281" points="317" swimtime="00:05:18.96" resultid="3442" heatid="5351" lane="2" entrytime="00:05:14.58">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.32" />
                    <SPLIT distance="100" swimtime="00:01:29.05" />
                    <SPLIT distance="150" swimtime="00:02:06.50" />
                    <SPLIT distance="200" swimtime="00:02:52.53" />
                    <SPLIT distance="250" swimtime="00:03:25.43" />
                    <SPLIT distance="300" swimtime="00:04:04.03" />
                    <SPLIT distance="350" swimtime="00:04:38.86" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3337" number="1" />
                    <RELAYPOSITION athleteid="3414" number="2" />
                    <RELAYPOSITION athleteid="3344" number="3" />
                    <RELAYPOSITION athleteid="3421" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="12782" nation="BRA" region="PR" clubid="4026" swrid="93773" name="Clube Duque De Caxias" shortname="Duque De Caxias">
          <ATHLETES>
            <ATHLETE firstname="Joao" lastname="Vitor Girelli" birthdate="2009-08-01" gender="M" nation="BRA" license="387965" swrid="5622312" athleteid="4031" externalid="387965">
              <RESULTS>
                <RESULT eventid="1072" points="393" swimtime="00:05:00.41" resultid="4032" heatid="5061" lane="7" entrytime="00:04:58.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.59" />
                    <SPLIT distance="100" swimtime="00:01:07.38" />
                    <SPLIT distance="150" swimtime="00:01:44.88" />
                    <SPLIT distance="200" swimtime="00:02:23.70" />
                    <SPLIT distance="250" swimtime="00:03:03.51" />
                    <SPLIT distance="300" swimtime="00:03:42.73" />
                    <SPLIT distance="350" swimtime="00:04:21.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="415" swimtime="00:00:28.03" resultid="4033" heatid="5122" lane="5" entrytime="00:00:28.53" entrycourse="LCM" />
                <RESULT eventid="1120" points="393" swimtime="00:02:19.23" resultid="4034" heatid="5154" lane="8" entrytime="00:02:20.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.38" />
                    <SPLIT distance="100" swimtime="00:01:05.58" />
                    <SPLIT distance="150" swimtime="00:01:42.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="441" swimtime="00:01:01.53" resultid="4035" heatid="5227" lane="7" entrytime="00:01:01.20" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="356" swimtime="00:00:33.22" resultid="4036" heatid="5285" lane="7" entrytime="00:00:35.39" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ian" lastname="Berger" birthdate="2011-07-27" gender="M" nation="BRA" license="387966" swrid="5652879" athleteid="4037" externalid="387966">
              <RESULTS>
                <RESULT eventid="1104" points="307" swimtime="00:00:30.98" resultid="4038" heatid="5116" lane="3" entrytime="00:00:31.47" entrycourse="LCM" />
                <RESULT eventid="1120" points="320" swimtime="00:02:29.09" resultid="4039" heatid="5150" lane="1" entrytime="00:02:29.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.30" />
                    <SPLIT distance="100" swimtime="00:01:09.60" />
                    <SPLIT distance="150" swimtime="00:01:48.90" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="345" swimtime="00:01:06.78" resultid="4040" heatid="5220" lane="4" entrytime="00:01:07.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.67" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Bulgarelli Castro" birthdate="2009-04-20" gender="M" nation="BRA" license="401867" swrid="5658058" athleteid="4041" externalid="401867">
              <RESULTS>
                <RESULT eventid="1104" points="340" swimtime="00:00:29.93" resultid="4042" heatid="5122" lane="8" entrytime="00:00:29.74" entrycourse="LCM" />
                <RESULT eventid="1120" points="281" swimtime="00:02:35.60" resultid="4043" heatid="5153" lane="6" entrytime="00:02:32.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.08" />
                    <SPLIT distance="100" swimtime="00:01:13.73" />
                    <SPLIT distance="150" swimtime="00:01:56.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="332" swimtime="00:01:07.61" resultid="4044" heatid="5225" lane="2" entrytime="00:01:06.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" status="DNS" swimtime="00:00:00.00" resultid="4045" heatid="5282" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Ana" lastname="Flavia Braz" birthdate="2004-10-25" gender="F" nation="BRA" license="280573" swrid="5622281" athleteid="4027" externalid="280573">
              <RESULTS>
                <RESULT eventid="1080" points="466" swimtime="00:01:22.69" resultid="4028" heatid="5070" lane="6" entrytime="00:01:23.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="447" swimtime="00:02:59.80" resultid="4029" heatid="5312" lane="5" entrytime="00:03:04.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.33" />
                    <SPLIT distance="100" swimtime="00:01:23.97" />
                    <SPLIT distance="150" swimtime="00:02:12.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="537" swimtime="00:00:35.86" resultid="4030" heatid="5377" lane="3" entrytime="00:00:36.50" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tayla" lastname="Kalluf Oliveira" birthdate="2011-12-05" gender="F" nation="BRA" license="414583" swrid="5755374" athleteid="4046" externalid="414583">
              <RESULTS>
                <RESULT eventid="1096" points="450" swimtime="00:00:30.81" resultid="4047" heatid="5099" lane="7" entrytime="00:00:31.61" entrycourse="LCM" />
                <RESULT eventid="1159" points="430" swimtime="00:01:08.50" resultid="4048" heatid="5204" lane="1" entrytime="00:01:08.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="385" swimtime="00:00:33.57" resultid="4049" heatid="5321" lane="5" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="15981" nation="BRA" region="PR" clubid="2398" swrid="93783" name="Quinto Nado" shortname="5º Nado">
          <ATHLETES>
            <ATHLETE firstname="Guilherme" lastname="Kikuchi Fujii" birthdate="2007-01-04" gender="M" nation="BRA" license="297805" swrid="5603863" athleteid="2399" externalid="297805" level="G-OLIMPICA">
              <RESULTS>
                <RESULT eventid="1088" points="638" swimtime="00:01:06.07" resultid="2400" heatid="5087" lane="5" entrytime="00:01:05.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="603" swimtime="00:00:58.52" resultid="2401" heatid="5178" lane="1" entrytime="00:00:58.41" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="526" swimtime="00:01:03.91" resultid="2402" heatid="5263" lane="8" entrytime="00:01:05.52" entrycourse="LCM" />
                <RESULT eventid="1267" points="596" swimtime="00:00:26.45" resultid="2403" heatid="5336" lane="7" entrytime="00:00:27.73" entrycourse="LCM" />
                <RESULT eventid="1251" points="642" swimtime="00:02:25.44" resultid="2404" heatid="5320" lane="5" entrytime="00:02:22.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.27" />
                    <SPLIT distance="100" swimtime="00:01:09.23" />
                    <SPLIT distance="150" swimtime="00:01:48.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="619" swimtime="00:00:30.44" resultid="2405" heatid="5371" lane="5" entrytime="00:00:30.65" entrycourse="LCM" />
                <RESULT eventid="2320" points="640" swimtime="00:01:06.00" resultid="5953" heatid="6414" lane="4" entrytime="00:01:06.07">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2335" points="602" swimtime="00:00:58.54" resultid="6011" heatid="6417" lane="6" entrytime="00:00:58.52">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Silva Telles" birthdate="2011-07-19" gender="M" nation="BRA" license="377311" swrid="5603911" athleteid="2427" externalid="377311">
              <RESULTS>
                <RESULT eventid="1088" points="247" swimtime="00:01:30.57" resultid="2428" heatid="5081" lane="8" entrytime="00:01:29.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="253" swimtime="00:00:33.02" resultid="2429" heatid="5116" lane="6" entrytime="00:00:32.91" entrycourse="LCM" />
                <RESULT eventid="1120" points="238" swimtime="00:02:44.50" resultid="2430" heatid="5148" lane="8">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:19.82" />
                    <SPLIT distance="150" swimtime="00:02:03.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="266" swimtime="00:01:12.78" resultid="2431" heatid="5217" lane="5" />
                <RESULT eventid="1251" points="249" swimtime="00:03:19.21" resultid="2432" heatid="5316" lane="2" entrytime="00:03:23.77" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.40" />
                    <SPLIT distance="100" swimtime="00:01:35.03" />
                    <SPLIT distance="150" swimtime="00:02:28.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="279" swimtime="00:00:39.70" resultid="2433" heatid="5364" lane="7" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Takemura Couto" birthdate="2010-02-08" gender="F" nation="BRA" license="376950" swrid="5603919" athleteid="2420" externalid="376950">
              <RESULTS>
                <RESULT eventid="1096" points="526" swimtime="00:00:29.24" resultid="2421" heatid="5100" lane="6" entrytime="00:00:29.27" entrycourse="LCM" />
                <RESULT eventid="1128" points="299" swimtime="00:01:22.96" resultid="2422" heatid="5159" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="338" swimtime="00:01:22.27" resultid="2423" heatid="5243" lane="2" entrytime="00:01:19.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="479" swimtime="00:01:06.06" resultid="2424" heatid="5205" lane="3" entrytime="00:01:05.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="417" swimtime="00:00:35.95" resultid="2425" heatid="5294" lane="6" entrytime="00:00:36.10" entrycourse="LCM" />
                <RESULT eventid="1259" points="450" swimtime="00:00:31.88" resultid="2426" heatid="5325" lane="4" entrytime="00:00:33.51" entrycourse="LCM" />
                <RESULT eventid="2375" points="521" swimtime="00:00:29.34" resultid="5977" heatid="5978" lane="8" entrytime="00:00:29.24" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Poletti Veiga" birthdate="2010-10-01" gender="F" nation="BRA" license="376951" swrid="5603895" athleteid="2413" externalid="376951">
              <RESULTS>
                <RESULT eventid="1064" points="460" swimtime="00:05:04.77" resultid="2414" heatid="5051" lane="6" entrytime="00:05:02.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.99" />
                    <SPLIT distance="100" swimtime="00:01:12.60" />
                    <SPLIT distance="150" swimtime="00:01:51.37" />
                    <SPLIT distance="200" swimtime="00:02:30.79" />
                    <SPLIT distance="250" swimtime="00:03:09.40" />
                    <SPLIT distance="300" swimtime="00:03:48.52" />
                    <SPLIT distance="350" swimtime="00:04:27.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="500" swimtime="00:02:22.13" resultid="2415" heatid="5141" lane="5" entrytime="00:02:21.46" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.19" />
                    <SPLIT distance="100" swimtime="00:01:09.84" />
                    <SPLIT distance="150" swimtime="00:01:46.78" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="412" swimtime="00:01:17.01" resultid="2416" heatid="5243" lane="5" entrytime="00:01:17.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="501" swimtime="00:01:05.10" resultid="2417" heatid="5205" lane="2" entrytime="00:01:05.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.40" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="439" swimtime="00:00:35.34" resultid="2418" heatid="5293" lane="4" entrytime="00:00:36.93" entrycourse="LCM" />
                <RESULT eventid="1275" points="425" swimtime="00:02:43.75" resultid="2419" heatid="5343" lane="8" entrytime="00:02:44.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                    <SPLIT distance="100" swimtime="00:01:20.91" />
                    <SPLIT distance="150" swimtime="00:02:02.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Bordini Zocco" birthdate="2008-08-04" gender="F" nation="BRA" license="385677" swrid="5332871" athleteid="2406" externalid="385677">
              <RESULTS>
                <RESULT eventid="1080" points="347" swimtime="00:01:31.26" resultid="2407" heatid="5068" lane="7" entrytime="00:01:32.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="388" swimtime="00:00:32.37" resultid="2408" heatid="5101" lane="5" />
                <RESULT eventid="1143" points="381" swimtime="00:02:53.95" resultid="2409" heatid="5189" lane="6" entrytime="00:02:53.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:21.89" />
                    <SPLIT distance="150" swimtime="00:02:13.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="347" swimtime="00:01:21.54" resultid="2410" heatid="5246" lane="2" entrytime="00:01:21.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1243" points="327" swimtime="00:03:19.64" resultid="2411" heatid="5311" lane="2" entrytime="00:03:24.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.99" />
                    <SPLIT distance="100" swimtime="00:01:35.38" />
                    <SPLIT distance="150" swimtime="00:02:27.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="344" swimtime="00:00:41.58" resultid="2412" heatid="5373" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benjamin" lastname="Rinaldi Batistao" birthdate="2010-07-13" gender="M" nation="BRA" license="407035" swrid="5737920" athleteid="2434" externalid="407035">
              <RESULTS>
                <RESULT eventid="1104" points="334" swimtime="00:00:30.12" resultid="2435" heatid="5115" lane="8" />
                <RESULT eventid="1120" points="277" swimtime="00:02:36.30" resultid="2436" heatid="5147" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                    <SPLIT distance="100" swimtime="00:01:13.93" />
                    <SPLIT distance="150" swimtime="00:01:55.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="303" swimtime="00:01:09.75" resultid="2437" heatid="5217" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="229" swimtime="00:00:38.45" resultid="2438" heatid="5282" lane="7" />
                <RESULT eventid="1267" points="302" swimtime="00:00:33.18" resultid="2439" heatid="5329" lane="6" />
                <RESULT eventid="1297" points="219" swimtime="00:00:43.04" resultid="2440" heatid="5363" lane="6" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="3501" nation="BRA" region="PR" clubid="2771" swrid="93752" name="Ortega &amp; De Souza Jesus" shortname="Aquafoz">
          <ATHLETES>
            <ATHLETE firstname="Julio" lastname="Heck" birthdate="1998-02-15" gender="M" nation="BRA" license="185880" swrid="5596906" athleteid="2789" externalid="185880">
              <RESULTS>
                <RESULT eventid="1104" points="624" swimtime="00:00:24.46" resultid="2790" heatid="5130" lane="1" entrytime="00:00:24.28" entrycourse="LCM" />
                <RESULT eventid="1167" points="671" swimtime="00:00:53.50" resultid="2791" heatid="5233" lane="8" entrytime="00:00:53.71" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="403" swimtime="00:00:31.88" resultid="2792" heatid="5286" lane="5" entrytime="00:00:31.55" entrycourse="LCM" />
                <RESULT eventid="1267" status="DNS" swimtime="00:00:00.00" resultid="2793" heatid="5337" lane="8" entrytime="00:00:27.44" entrycourse="LCM" />
                <RESULT eventid="2383" points="628" swimtime="00:00:24.41" resultid="5983" heatid="6425" lane="2" entrytime="00:00:24.46" />
                <RESULT eventid="2351" points="655" swimtime="00:00:53.95" resultid="6120" heatid="6422" lane="2" entrytime="00:00:53.50">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.70" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Gabriel Serighelli" birthdate="1999-03-12" gender="M" nation="BRA" license="121253" swrid="5596899" athleteid="2779" externalid="121253">
              <RESULTS>
                <RESULT eventid="1104" points="557" swimtime="00:00:25.40" resultid="2780" heatid="5129" lane="5" entrytime="00:00:24.84" entrycourse="LCM" />
                <RESULT eventid="1135" points="496" swimtime="00:01:02.44" resultid="2781" heatid="5177" lane="7" entrytime="00:01:03.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="531" swimtime="00:00:29.08" resultid="2782" heatid="5287" lane="4" entrytime="00:00:28.84" entrycourse="LCM" />
                <RESULT eventid="1267" points="563" swimtime="00:00:26.96" resultid="2783" heatid="5337" lane="4" entrytime="00:00:26.84" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leticia" lastname="Marques Lima" birthdate="2010-04-30" gender="F" nation="BRA" license="383051" swrid="5596913" athleteid="2824" externalid="383051">
              <RESULTS>
                <RESULT eventid="1096" points="370" swimtime="00:00:32.86" resultid="2825" heatid="5097" lane="4" entrytime="00:00:34.53" entrycourse="LCM" />
                <RESULT eventid="1128" points="260" swimtime="00:01:26.87" resultid="2826" heatid="5159" lane="4" entrytime="00:01:28.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="337" swimtime="00:01:22.37" resultid="2827" heatid="5243" lane="1" entrytime="00:01:22.01" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="356" swimtime="00:00:37.89" resultid="2828" heatid="5293" lane="3" entrytime="00:00:37.66" entrycourse="LCM" />
                <RESULT eventid="1259" points="363" swimtime="00:00:34.24" resultid="2829" heatid="5324" lane="2" entrytime="00:00:36.41" entrycourse="LCM" />
                <RESULT eventid="1275" points="310" swimtime="00:03:01.76" resultid="2830" heatid="5340" lane="4" entrytime="00:02:57.95" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.15" />
                    <SPLIT distance="100" swimtime="00:01:28.87" />
                    <SPLIT distance="150" swimtime="00:02:16.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yago" lastname="Simon Pires" birthdate="2008-10-29" gender="M" nation="BRA" license="328942" swrid="5596939" athleteid="2800" externalid="328942">
              <RESULTS>
                <RESULT eventid="1104" points="498" swimtime="00:00:26.38" resultid="2801" heatid="5125" lane="2" entrytime="00:00:26.30" entrycourse="LCM" />
                <RESULT eventid="1120" points="394" swimtime="00:02:19.11" resultid="2802" heatid="5155" lane="7" entrytime="00:02:14.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.76" />
                    <SPLIT distance="100" swimtime="00:01:04.33" />
                    <SPLIT distance="150" swimtime="00:01:41.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="511" swimtime="00:00:58.59" resultid="2803" heatid="5228" lane="6" entrytime="00:00:58.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="439" swimtime="00:00:34.12" resultid="2804" heatid="5369" lane="8" entrytime="00:00:35.59" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mateus" lastname="Wirtti" birthdate="2011-01-14" gender="M" nation="BRA" license="383854" swrid="4917570" athleteid="2831" externalid="383854">
              <RESULTS>
                <RESULT eventid="1104" points="350" swimtime="00:00:29.65" resultid="2832" heatid="5118" lane="8" entrytime="00:00:29.86" entrycourse="LCM" />
                <RESULT eventid="1120" points="292" swimtime="00:02:33.72" resultid="2833" heatid="5149" lane="4" entrytime="00:02:32.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                    <SPLIT distance="100" swimtime="00:01:11.49" />
                    <SPLIT distance="150" swimtime="00:01:53.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="369" swimtime="00:01:05.29" resultid="2834" heatid="5220" lane="2" entrytime="00:01:08.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="291" swimtime="00:00:35.53" resultid="2835" heatid="5285" lane="1" entrytime="00:00:35.71" entrycourse="LCM" />
                <RESULT eventid="1267" points="262" swimtime="00:00:34.80" resultid="2836" heatid="5331" lane="3" entrytime="00:00:35.88" entrycourse="LCM" />
                <RESULT eventid="1297" points="215" swimtime="00:00:43.31" resultid="2837" heatid="5363" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Mussi" birthdate="2006-12-31" gender="M" nation="BRA" license="370567" swrid="5596917" athleteid="2812" externalid="370567">
              <RESULTS>
                <RESULT eventid="1088" points="408" swimtime="00:01:16.63" resultid="2813" heatid="5086" lane="4" entrytime="00:01:17.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.11" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="368" swimtime="00:00:32.85" resultid="2814" heatid="5285" lane="6" entrytime="00:00:33.87" entrycourse="LCM" />
                <RESULT comment="SW 7.6 - Não tocou a borda na virada ou na chegada com ambas as mãos; separadamente; simultaneamente.  (Horário: 9:45), Na volta dos 100m." eventid="1251" status="DSQ" swimtime="00:02:58.94" resultid="2815" heatid="5315" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                    <SPLIT distance="100" swimtime="00:01:27.40" />
                    <SPLIT distance="150" swimtime="00:02:13.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="518" swimtime="00:00:32.30" resultid="2816" heatid="5370" lane="6" entrytime="00:00:33.49" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Gustavo Cunha" birthdate="2011-01-31" gender="M" nation="BRA" license="392836" swrid="5641764" athleteid="2845" externalid="392836">
              <RESULTS>
                <RESULT eventid="1088" points="155" swimtime="00:01:45.87" resultid="2846" heatid="5078" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="252" swimtime="00:00:33.08" resultid="2847" heatid="5114" lane="5" />
                <RESULT eventid="1151" points="152" swimtime="00:03:33.32" resultid="2848" heatid="5192" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.40" />
                    <SPLIT distance="150" swimtime="00:02:47.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="262" swimtime="00:01:13.23" resultid="2849" heatid="5217" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="143" swimtime="00:03:59.54" resultid="2850" heatid="5315" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.22" />
                    <SPLIT distance="100" swimtime="00:01:54.95" />
                    <SPLIT distance="150" swimtime="00:02:58.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="179" swimtime="00:00:46.04" resultid="2851" heatid="5363" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="De Souza Tulio" birthdate="2006-06-23" gender="F" nation="BRA" license="342344" swrid="5030980" athleteid="2772" externalid="342344">
              <RESULTS>
                <RESULT eventid="1064" points="514" swimtime="00:04:53.77" resultid="2773" heatid="5055" lane="6" entrytime="00:04:40.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.51" />
                    <SPLIT distance="100" swimtime="00:01:06.84" />
                    <SPLIT distance="150" swimtime="00:01:43.59" />
                    <SPLIT distance="200" swimtime="00:02:21.19" />
                    <SPLIT distance="250" swimtime="00:02:59.44" />
                    <SPLIT distance="300" swimtime="00:03:37.92" />
                    <SPLIT distance="350" swimtime="00:04:16.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="534" swimtime="00:02:19.07" resultid="2774" heatid="5146" lane="3" entrytime="00:02:10.02" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.33" />
                    <SPLIT distance="100" swimtime="00:01:06.67" />
                    <SPLIT distance="150" swimtime="00:01:43.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="509" swimtime="00:01:11.78" resultid="2775" heatid="5248" lane="5" entrytime="00:01:08.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="567" swimtime="00:01:02.45" resultid="2776" heatid="5209" lane="5" entrytime="00:01:00.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="590" swimtime="00:00:32.01" resultid="2777" heatid="5295" lane="3" entrytime="00:00:32.07" entrycourse="LCM" />
                <RESULT eventid="1275" points="437" swimtime="00:02:42.22" resultid="2778" heatid="5343" lane="4" entrytime="00:02:31.00" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.62" />
                    <SPLIT distance="100" swimtime="00:01:16.47" />
                    <SPLIT distance="150" swimtime="00:01:59.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2343" points="562" swimtime="00:01:02.66" resultid="6105" heatid="6421" lane="2" entrytime="00:01:02.45">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2391" points="536" swimtime="00:01:10.54" resultid="6131" heatid="6424" lane="6" entrytime="00:01:11.78">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.68" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauan" lastname="Matheus Cunha" birthdate="2011-01-31" gender="M" nation="BRA" license="392834" swrid="5641770" athleteid="2838" externalid="392834">
              <RESULTS>
                <RESULT eventid="1072" points="172" swimtime="00:06:35.20" resultid="2839" heatid="5056" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.08" />
                    <SPLIT distance="100" swimtime="00:01:29.75" />
                    <SPLIT distance="150" swimtime="00:02:20.43" />
                    <SPLIT distance="200" swimtime="00:03:11.02" />
                    <SPLIT distance="250" swimtime="00:04:01.99" />
                    <SPLIT distance="300" swimtime="00:04:53.47" />
                    <SPLIT distance="350" swimtime="00:05:45.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="273" swimtime="00:00:32.21" resultid="2840" heatid="5114" lane="4" />
                <RESULT eventid="1135" points="126" swimtime="00:01:38.63" resultid="2841" heatid="5169" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="256" swimtime="00:01:13.72" resultid="2842" heatid="5218" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="178" swimtime="00:00:41.82" resultid="2843" heatid="5281" lane="4" />
                <RESULT eventid="1267" points="220" swimtime="00:00:36.88" resultid="2844" heatid="5330" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Xavier" birthdate="2011-10-14" gender="M" nation="BRA" license="370564" swrid="5596949" athleteid="2805" externalid="370564">
              <RESULTS>
                <RESULT eventid="1088" points="255" swimtime="00:01:29.66" resultid="2806" heatid="5080" lane="2" entrytime="00:01:31.68" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="191" swimtime="00:00:36.30" resultid="2807" heatid="5115" lane="3" entrytime="00:00:35.83" entrycourse="LCM" />
                <RESULT eventid="1120" points="194" swimtime="00:02:56.18" resultid="2808" heatid="5148" lane="5" entrytime="00:02:59.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.21" />
                    <SPLIT distance="100" swimtime="00:01:25.64" />
                    <SPLIT distance="150" swimtime="00:02:12.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="218" swimtime="00:01:17.76" resultid="2809" heatid="5218" lane="5" entrytime="00:01:18.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="276" swimtime="00:03:12.57" resultid="2810" heatid="5316" lane="6" entrytime="00:03:20.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.47" />
                    <SPLIT distance="100" swimtime="00:01:34.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="268" swimtime="00:00:40.20" resultid="2811" heatid="5366" lane="2" entrytime="00:00:47.72" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Geórgia" lastname="Adeli Jesus" birthdate="2008-03-27" gender="F" nation="BRA" license="312649" swrid="5596864" athleteid="2794" externalid="312649">
              <RESULTS>
                <RESULT eventid="1064" points="403" swimtime="00:05:18.48" resultid="2795" heatid="5053" lane="1" entrytime="00:05:25.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.98" />
                    <SPLIT distance="100" swimtime="00:01:13.22" />
                    <SPLIT distance="150" swimtime="00:01:53.16" />
                    <SPLIT distance="200" swimtime="00:02:34.61" />
                    <SPLIT distance="250" swimtime="00:03:16.24" />
                    <SPLIT distance="300" swimtime="00:03:57.21" />
                    <SPLIT distance="350" swimtime="00:04:38.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="439" swimtime="00:02:28.40" resultid="2796" heatid="5143" lane="7" entrytime="00:02:31.54" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.41" />
                    <SPLIT distance="100" swimtime="00:01:10.76" />
                    <SPLIT distance="150" swimtime="00:01:49.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="364" swimtime="00:11:18.58" resultid="2797" heatid="5272" lane="2" entrytime="00:11:10.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.07" />
                    <SPLIT distance="100" swimtime="00:01:14.47" />
                    <SPLIT distance="150" swimtime="00:01:54.83" />
                    <SPLIT distance="200" swimtime="00:02:36.70" />
                    <SPLIT distance="250" swimtime="00:03:18.51" />
                    <SPLIT distance="300" swimtime="00:04:00.92" />
                    <SPLIT distance="350" swimtime="00:04:43.63" />
                    <SPLIT distance="400" swimtime="00:05:27.12" />
                    <SPLIT distance="450" swimtime="00:06:10.24" />
                    <SPLIT distance="500" swimtime="00:06:54.20" />
                    <SPLIT distance="550" swimtime="00:07:38.42" />
                    <SPLIT distance="600" swimtime="00:08:23.66" />
                    <SPLIT distance="650" swimtime="00:09:07.75" />
                    <SPLIT distance="700" swimtime="00:09:52.05" />
                    <SPLIT distance="750" swimtime="00:10:36.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="377" swimtime="00:00:37.17" resultid="2798" heatid="5290" lane="1" />
                <RESULT eventid="1279" points="340" swimtime="00:21:58.08" resultid="2799" heatid="5349" lane="3" entrytime="00:21:33.75" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.73" />
                    <SPLIT distance="100" swimtime="00:01:14.86" />
                    <SPLIT distance="150" swimtime="00:01:55.91" />
                    <SPLIT distance="200" swimtime="00:02:38.19" />
                    <SPLIT distance="250" swimtime="00:03:20.64" />
                    <SPLIT distance="300" swimtime="00:04:04.52" />
                    <SPLIT distance="350" swimtime="00:04:47.78" />
                    <SPLIT distance="400" swimtime="00:05:32.37" />
                    <SPLIT distance="450" swimtime="00:06:17.05" />
                    <SPLIT distance="500" swimtime="00:07:01.74" />
                    <SPLIT distance="550" swimtime="00:07:45.14" />
                    <SPLIT distance="600" swimtime="00:08:29.63" />
                    <SPLIT distance="650" swimtime="00:09:14.58" />
                    <SPLIT distance="700" swimtime="00:09:59.64" />
                    <SPLIT distance="750" swimtime="00:10:45.33" />
                    <SPLIT distance="800" swimtime="00:11:30.72" />
                    <SPLIT distance="850" swimtime="00:12:16.13" />
                    <SPLIT distance="900" swimtime="00:13:01.16" />
                    <SPLIT distance="950" swimtime="00:13:47.57" />
                    <SPLIT distance="1000" swimtime="00:14:33.59" />
                    <SPLIT distance="1050" swimtime="00:15:18.73" />
                    <SPLIT distance="1100" swimtime="00:16:04.48" />
                    <SPLIT distance="1150" swimtime="00:16:48.58" />
                    <SPLIT distance="1200" swimtime="00:17:33.39" />
                    <SPLIT distance="1250" swimtime="00:18:17.59" />
                    <SPLIT distance="1300" swimtime="00:19:01.63" />
                    <SPLIT distance="1350" swimtime="00:19:45.13" />
                    <SPLIT distance="1400" swimtime="00:20:29.81" />
                    <SPLIT distance="1450" swimtime="00:21:13.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Dominguez Olivieski" birthdate="2011-04-27" gender="M" nation="BRA" license="405717" swrid="5664737" athleteid="2852" externalid="405717">
              <RESULTS>
                <RESULT eventid="1088" points="185" swimtime="00:01:39.69" resultid="2853" heatid="5079" lane="3" entrytime="00:01:37.09" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="244" swimtime="00:00:33.45" resultid="2854" heatid="5116" lane="2" entrytime="00:00:33.58" entrycourse="LCM" />
                <RESULT eventid="1167" points="262" swimtime="00:01:13.23" resultid="2855" heatid="5218" lane="3" entrytime="00:01:19.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="167" swimtime="00:00:42.70" resultid="2856" heatid="5284" lane="1" entrytime="00:00:42.69" entrycourse="LCM" />
                <RESULT eventid="1251" points="167" swimtime="00:03:47.75" resultid="2857" heatid="5315" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.28" />
                    <SPLIT distance="100" swimtime="00:01:47.63" />
                    <SPLIT distance="150" swimtime="00:02:50.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="193" swimtime="00:00:44.87" resultid="2858" heatid="5364" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Afonso Proteti" birthdate="2002-03-19" gender="M" nation="BRA" license="190464" swrid="5596865" athleteid="2784" externalid="190464">
              <RESULTS>
                <RESULT eventid="1135" points="600" swimtime="00:00:58.60" resultid="2785" heatid="5178" lane="6" entrytime="00:00:57.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="568" swimtime="00:01:02.28" resultid="2786" heatid="5263" lane="6" entrytime="00:01:01.58" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="557" swimtime="00:00:28.62" resultid="2787" heatid="5288" lane="7" entrytime="00:00:28.76" entrycourse="LCM" />
                <RESULT eventid="1267" points="672" swimtime="00:00:25.42" resultid="2788" heatid="5338" lane="5" entrytime="00:00:25.19" entrycourse="LCM" />
                <RESULT eventid="2335" points="603" swimtime="00:00:58.53" resultid="6013" heatid="6417" lane="7" entrytime="00:00:58.60">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2359" points="560" swimtime="00:01:02.57" resultid="6147" heatid="6423" lane="2" entrytime="00:01:02.28">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Victoria Portela" birthdate="2009-12-04" gender="F" nation="BRA" license="383047" swrid="5596945" athleteid="2817" externalid="383047">
              <RESULTS>
                <RESULT eventid="1096" points="533" swimtime="00:00:29.11" resultid="2818" heatid="5104" lane="8" entrytime="00:00:29.56" entrycourse="LCM" />
                <RESULT eventid="1112" points="392" swimtime="00:02:34.14" resultid="2819" heatid="5143" lane="6" entrytime="00:02:30.45" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.02" />
                    <SPLIT distance="100" swimtime="00:01:09.67" />
                    <SPLIT distance="150" swimtime="00:01:50.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" status="DNS" swimtime="00:00:00.00" resultid="2820" heatid="5245" lane="3" />
                <RESULT eventid="1159" points="500" swimtime="00:01:05.15" resultid="2821" heatid="5207" lane="6" entrytime="00:01:06.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="330" swimtime="00:00:38.83" resultid="2822" heatid="5290" lane="6" />
                <RESULT eventid="1305" points="373" swimtime="00:00:40.48" resultid="2823" heatid="5372" lane="3" />
                <RESULT eventid="2375" points="509" swimtime="00:00:29.56" resultid="5976" heatid="5978" lane="1" entrytime="00:00:29.11" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="-1" agemin="20" agetotalmax="-1" agetotalmin="-1" gender="M" name="AQUAFOZ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1241" points="580" swimtime="00:03:45.64" resultid="2859" heatid="5310" lane="6" entrytime="00:03:41.90">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.64" />
                    <SPLIT distance="100" swimtime="00:00:56.67" />
                    <SPLIT distance="150" swimtime="00:01:24.64" />
                    <SPLIT distance="200" swimtime="00:01:57.59" />
                    <SPLIT distance="250" swimtime="00:02:23.71" />
                    <SPLIT distance="300" swimtime="00:02:52.89" />
                    <SPLIT distance="350" swimtime="00:03:17.78" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2779" number="1" />
                    <RELAYPOSITION athleteid="2812" number="2" />
                    <RELAYPOSITION athleteid="2784" number="3" />
                    <RELAYPOSITION athleteid="2789" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1342" points="542" swimtime="00:04:13.60" resultid="2861" heatid="5390" lane="6" entrytime="00:04:13.12">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.28" />
                    <SPLIT distance="100" swimtime="00:01:06.02" />
                    <SPLIT distance="150" swimtime="00:01:40.38" />
                    <SPLIT distance="200" swimtime="00:02:21.04" />
                    <SPLIT distance="250" swimtime="00:02:48.01" />
                    <SPLIT distance="300" swimtime="00:03:19.54" />
                    <SPLIT distance="350" swimtime="00:03:45.09" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2779" number="1" />
                    <RELAYPOSITION athleteid="2812" number="2" />
                    <RELAYPOSITION athleteid="2784" number="3" />
                    <RELAYPOSITION athleteid="2789" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="13" agemin="13" agetotalmax="-1" agetotalmin="-1" gender="M" name="AQUAFOZ &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1231" points="285" swimtime="00:04:45.78" resultid="2860" heatid="5305" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.26" />
                    <SPLIT distance="100" swimtime="00:01:11.93" />
                    <SPLIT distance="150" swimtime="00:01:46.18" />
                    <SPLIT distance="250" swimtime="00:03:00.35" />
                    <SPLIT distance="300" swimtime="00:03:40.15" />
                    <SPLIT distance="350" swimtime="00:04:10.71" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2845" number="1" />
                    <RELAYPOSITION athleteid="2852" number="2" />
                    <RELAYPOSITION athleteid="2838" number="3" />
                    <RELAYPOSITION athleteid="2831" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1332" points="238" swimtime="00:05:33.23" resultid="2862" heatid="5385" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.35" />
                    <SPLIT distance="100" swimtime="00:01:18.78" />
                    <SPLIT distance="150" swimtime="00:02:00.21" />
                    <SPLIT distance="200" swimtime="00:02:48.26" />
                    <SPLIT distance="250" swimtime="00:03:27.45" />
                    <SPLIT distance="300" swimtime="00:04:21.87" />
                    <SPLIT distance="350" swimtime="00:04:54.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="2831" number="1" />
                    <RELAYPOSITION athleteid="2805" number="2" />
                    <RELAYPOSITION athleteid="2838" number="3" />
                    <RELAYPOSITION athleteid="2845" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="CLUB" code="2539" nation="BRA" region="PR" clubid="3177" swrid="93771" name="Círculo Militar Do Paraná" shortname="Círculo Militar">
          <ATHLETES>
            <ATHLETE firstname="Gabriel" lastname="Manocchio" birthdate="2011-07-28" gender="M" nation="BRA" license="384916" swrid="5588573" athleteid="3201" externalid="384916">
              <RESULTS>
                <RESULT eventid="1088" points="258" swimtime="00:01:29.34" resultid="3202" heatid="5080" lane="3" entrytime="00:01:30.56" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="350" swimtime="00:00:29.65" resultid="3203" heatid="5118" lane="6" entrytime="00:00:29.31" entrycourse="LCM" />
                <RESULT eventid="1120" points="376" swimtime="00:02:21.21" resultid="3204" heatid="5150" lane="3" entrytime="00:02:26.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.63" />
                    <SPLIT distance="100" swimtime="00:01:06.90" />
                    <SPLIT distance="150" swimtime="00:01:44.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="411" swimtime="00:01:03.00" resultid="3205" heatid="5221" lane="2" entrytime="00:01:05.31" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="359" swimtime="00:10:35.76" resultid="3206" heatid="5297" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.93" />
                    <SPLIT distance="100" swimtime="00:01:15.80" />
                    <SPLIT distance="150" swimtime="00:01:57.79" />
                    <SPLIT distance="200" swimtime="00:02:39.17" />
                    <SPLIT distance="250" swimtime="00:03:20.87" />
                    <SPLIT distance="300" swimtime="00:04:03.54" />
                    <SPLIT distance="350" swimtime="00:04:45.02" />
                    <SPLIT distance="400" swimtime="00:05:24.66" />
                    <SPLIT distance="450" swimtime="00:06:03.68" />
                    <SPLIT distance="500" swimtime="00:06:45.16" />
                    <SPLIT distance="550" swimtime="00:07:25.02" />
                    <SPLIT distance="600" swimtime="00:08:03.47" />
                    <SPLIT distance="650" swimtime="00:08:41.34" />
                    <SPLIT distance="700" swimtime="00:09:20.89" />
                    <SPLIT distance="750" swimtime="00:09:59.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="342" swimtime="00:20:44.96" resultid="3207" heatid="5379" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.98" />
                    <SPLIT distance="100" swimtime="00:01:16.79" />
                    <SPLIT distance="150" swimtime="00:02:00.21" />
                    <SPLIT distance="200" swimtime="00:02:42.85" />
                    <SPLIT distance="250" swimtime="00:03:25.89" />
                    <SPLIT distance="300" swimtime="00:04:07.81" />
                    <SPLIT distance="350" swimtime="00:04:51.20" />
                    <SPLIT distance="400" swimtime="00:05:33.58" />
                    <SPLIT distance="450" swimtime="00:06:15.81" />
                    <SPLIT distance="500" swimtime="00:06:57.87" />
                    <SPLIT distance="550" swimtime="00:07:40.55" />
                    <SPLIT distance="600" swimtime="00:08:22.50" />
                    <SPLIT distance="650" swimtime="00:09:06.62" />
                    <SPLIT distance="700" swimtime="00:09:50.17" />
                    <SPLIT distance="750" swimtime="00:10:34.20" />
                    <SPLIT distance="800" swimtime="00:11:14.96" />
                    <SPLIT distance="850" swimtime="00:11:57.65" />
                    <SPLIT distance="900" swimtime="00:12:39.68" />
                    <SPLIT distance="950" swimtime="00:13:22.94" />
                    <SPLIT distance="1000" swimtime="00:14:05.13" />
                    <SPLIT distance="1050" swimtime="00:14:47.15" />
                    <SPLIT distance="1100" swimtime="00:15:28.34" />
                    <SPLIT distance="1150" swimtime="00:16:09.36" />
                    <SPLIT distance="1200" swimtime="00:16:49.71" />
                    <SPLIT distance="1250" swimtime="00:17:31.88" />
                    <SPLIT distance="1300" swimtime="00:18:12.23" />
                    <SPLIT distance="1350" swimtime="00:18:52.75" />
                    <SPLIT distance="1400" swimtime="00:19:32.15" />
                    <SPLIT distance="1450" swimtime="00:20:10.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Torres Oliveira" birthdate="2008-04-10" gender="M" nation="BRA" license="400274" swrid="5653303" athleteid="3178" externalid="400274">
              <RESULTS>
                <RESULT eventid="1104" points="361" swimtime="00:00:29.35" resultid="3179" heatid="5123" lane="8" entrytime="00:00:28.38" entrycourse="LCM" />
                <RESULT eventid="1120" points="337" swimtime="00:02:26.44" resultid="3180" heatid="5153" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.43" />
                    <SPLIT distance="100" swimtime="00:01:06.52" />
                    <SPLIT distance="150" swimtime="00:01:46.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="410" swimtime="00:01:03.03" resultid="3181" heatid="5226" lane="7" entrytime="00:01:03.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="292" swimtime="00:11:21.39" resultid="3182" heatid="5296" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.57" />
                    <SPLIT distance="100" swimtime="00:01:14.29" />
                    <SPLIT distance="150" swimtime="00:01:57.97" />
                    <SPLIT distance="200" swimtime="00:02:42.04" />
                    <SPLIT distance="250" swimtime="00:03:26.69" />
                    <SPLIT distance="300" swimtime="00:04:11.46" />
                    <SPLIT distance="350" swimtime="00:04:55.58" />
                    <SPLIT distance="400" swimtime="00:05:39.34" />
                    <SPLIT distance="450" swimtime="00:06:21.85" />
                    <SPLIT distance="500" swimtime="00:07:06.63" />
                    <SPLIT distance="550" swimtime="00:07:49.26" />
                    <SPLIT distance="600" swimtime="00:08:33.52" />
                    <SPLIT distance="650" swimtime="00:09:17.53" />
                    <SPLIT distance="700" swimtime="00:10:03.67" />
                    <SPLIT distance="750" swimtime="00:10:44.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="270" swimtime="00:22:26.45" resultid="3183" heatid="5378" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.78" />
                    <SPLIT distance="100" swimtime="00:01:12.66" />
                    <SPLIT distance="150" swimtime="00:01:57.09" />
                    <SPLIT distance="200" swimtime="00:02:42.50" />
                    <SPLIT distance="250" swimtime="00:03:29.16" />
                    <SPLIT distance="300" swimtime="00:04:16.11" />
                    <SPLIT distance="350" swimtime="00:05:00.70" />
                    <SPLIT distance="400" swimtime="00:05:46.48" />
                    <SPLIT distance="450" swimtime="00:06:31.90" />
                    <SPLIT distance="500" swimtime="00:07:17.70" />
                    <SPLIT distance="550" swimtime="00:08:04.01" />
                    <SPLIT distance="600" swimtime="00:08:50.33" />
                    <SPLIT distance="650" swimtime="00:09:37.58" />
                    <SPLIT distance="700" swimtime="00:10:23.20" />
                    <SPLIT distance="750" swimtime="00:11:07.62" />
                    <SPLIT distance="800" swimtime="00:11:53.80" />
                    <SPLIT distance="850" swimtime="00:12:40.74" />
                    <SPLIT distance="900" swimtime="00:13:26.85" />
                    <SPLIT distance="950" swimtime="00:14:11.99" />
                    <SPLIT distance="1000" swimtime="00:14:59.11" />
                    <SPLIT distance="1050" swimtime="00:15:45.51" />
                    <SPLIT distance="1100" swimtime="00:16:31.35" />
                    <SPLIT distance="1150" swimtime="00:17:16.84" />
                    <SPLIT distance="1200" swimtime="00:18:03.23" />
                    <SPLIT distance="1250" swimtime="00:18:47.96" />
                    <SPLIT distance="1300" swimtime="00:19:33.41" />
                    <SPLIT distance="1350" swimtime="00:20:17.79" />
                    <SPLIT distance="1400" swimtime="00:21:01.35" />
                    <SPLIT distance="1450" swimtime="00:21:45.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Odirlei" lastname="Garcia Nascimento" birthdate="1978-03-03" gender="M" nation="BRA" license="415758" athleteid="3225" externalid="415758">
              <RESULTS>
                <RESULT eventid="1267" points="326" swimtime="00:00:32.33" resultid="3226" heatid="5329" lane="3" />
                <RESULT eventid="1297" status="DNS" swimtime="00:00:00.00" resultid="3227" heatid="5363" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Thomas" lastname="Gomes" birthdate="2009-06-15" gender="M" nation="BRA" license="406948" swrid="5717268" athleteid="3208" externalid="406948">
              <RESULTS>
                <RESULT eventid="1072" points="216" swimtime="00:06:06.33" resultid="3209" heatid="5060" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.13" />
                    <SPLIT distance="100" swimtime="00:01:23.81" />
                    <SPLIT distance="150" swimtime="00:02:10.10" />
                    <SPLIT distance="200" swimtime="00:02:57.88" />
                    <SPLIT distance="250" swimtime="00:03:46.63" />
                    <SPLIT distance="300" swimtime="00:04:34.68" />
                    <SPLIT distance="350" swimtime="00:05:22.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="217" swimtime="00:02:49.72" resultid="3210" heatid="5153" lane="1" entrytime="00:02:47.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.25" />
                    <SPLIT distance="100" swimtime="00:01:20.65" />
                    <SPLIT distance="150" swimtime="00:02:05.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="246" swimtime="00:01:14.77" resultid="3211" heatid="5224" lane="4" entrytime="00:01:16.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruno" lastname="Yamamoto" birthdate="2006-04-22" gender="M" nation="BRA" license="336569" swrid="5717304" athleteid="3184" externalid="336569">
              <RESULTS>
                <RESULT eventid="1267" points="409" swimtime="00:00:29.98" resultid="3185" heatid="5329" lane="8" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernando" lastname="Jun Melo Ogima" birthdate="2006-07-05" gender="M" nation="BRA" license="378332" swrid="5622284" athleteid="3190" externalid="378332">
              <RESULTS>
                <RESULT eventid="1088" points="270" swimtime="00:01:27.93" resultid="3191" heatid="5086" lane="6" entrytime="00:01:27.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="413" swimtime="00:00:28.07" resultid="3192" heatid="5128" lane="8" entrytime="00:00:28.23" entrycourse="LCM" />
                <RESULT eventid="1151" points="289" swimtime="00:02:52.26" resultid="3193" heatid="5199" lane="4" entrytime="00:02:51.74" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.80" />
                    <SPLIT distance="100" swimtime="00:01:20.31" />
                    <SPLIT distance="150" swimtime="00:02:13.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="428" swimtime="00:01:02.18" resultid="3194" heatid="5231" lane="5" entrytime="00:01:02.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.45" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="372" swimtime="00:00:30.96" resultid="3195" heatid="5332" lane="6" entrytime="00:00:32.61" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicole" lastname="Herdy Faria" birthdate="2009-11-10" gender="F" nation="BRA" license="417277" athleteid="3228" externalid="417277">
              <RESULTS>
                <RESULT eventid="1064" points="293" swimtime="00:05:54.33" resultid="3229" heatid="5052" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="100" swimtime="00:01:19.67" />
                    <SPLIT distance="150" swimtime="00:02:04.30" />
                    <SPLIT distance="200" swimtime="00:02:49.79" />
                    <SPLIT distance="250" swimtime="00:03:36.36" />
                    <SPLIT distance="300" swimtime="00:04:22.88" />
                    <SPLIT distance="350" swimtime="00:05:09.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="370" swimtime="00:00:32.87" resultid="3230" heatid="5101" lane="4" />
                <RESULT eventid="1159" points="383" swimtime="00:01:11.18" resultid="3231" heatid="5206" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Henrique" lastname="Karuta" birthdate="2011-10-31" gender="M" nation="BRA" license="414648" swrid="5755375" athleteid="3220" externalid="414648">
              <RESULTS>
                <RESULT eventid="1072" points="250" swimtime="00:05:48.91" resultid="3221" heatid="5057" lane="8" entrytime="00:05:53.27" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.72" />
                    <SPLIT distance="100" swimtime="00:01:23.24" />
                    <SPLIT distance="150" swimtime="00:02:07.84" />
                    <SPLIT distance="200" swimtime="00:02:52.69" />
                    <SPLIT distance="250" swimtime="00:03:37.27" />
                    <SPLIT distance="300" swimtime="00:04:22.53" />
                    <SPLIT distance="350" swimtime="00:05:06.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="236" swimtime="00:02:44.83" resultid="3222" heatid="5147" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                    <SPLIT distance="100" swimtime="00:01:21.20" />
                    <SPLIT distance="150" swimtime="00:02:03.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="262" swimtime="00:11:46.48" resultid="3223" heatid="5297" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.72" />
                    <SPLIT distance="100" swimtime="00:01:21.13" />
                    <SPLIT distance="150" swimtime="00:02:05.24" />
                    <SPLIT distance="200" swimtime="00:02:49.74" />
                    <SPLIT distance="250" swimtime="00:03:34.00" />
                    <SPLIT distance="300" swimtime="00:04:19.18" />
                    <SPLIT distance="350" swimtime="00:05:04.24" />
                    <SPLIT distance="400" swimtime="00:05:49.62" />
                    <SPLIT distance="450" swimtime="00:06:34.55" />
                    <SPLIT distance="500" swimtime="00:07:19.95" />
                    <SPLIT distance="550" swimtime="00:08:04.89" />
                    <SPLIT distance="600" swimtime="00:08:50.40" />
                    <SPLIT distance="650" swimtime="00:09:35.20" />
                    <SPLIT distance="700" swimtime="00:10:19.66" />
                    <SPLIT distance="750" swimtime="00:11:03.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="272" swimtime="00:22:23.62" resultid="3224" heatid="5379" lane="1" entrytime="00:23:35.30" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.79" />
                    <SPLIT distance="100" swimtime="00:01:24.96" />
                    <SPLIT distance="150" swimtime="00:02:10.32" />
                    <SPLIT distance="200" swimtime="00:02:56.33" />
                    <SPLIT distance="250" swimtime="00:03:41.53" />
                    <SPLIT distance="300" swimtime="00:04:27.55" />
                    <SPLIT distance="350" swimtime="00:05:12.49" />
                    <SPLIT distance="400" swimtime="00:05:58.58" />
                    <SPLIT distance="450" swimtime="00:06:43.73" />
                    <SPLIT distance="500" swimtime="00:07:30.06" />
                    <SPLIT distance="550" swimtime="00:08:15.00" />
                    <SPLIT distance="600" swimtime="00:09:00.35" />
                    <SPLIT distance="650" swimtime="00:09:44.86" />
                    <SPLIT distance="700" swimtime="00:10:30.19" />
                    <SPLIT distance="750" swimtime="00:11:14.96" />
                    <SPLIT distance="800" swimtime="00:12:00.16" />
                    <SPLIT distance="850" swimtime="00:12:44.69" />
                    <SPLIT distance="900" swimtime="00:13:29.99" />
                    <SPLIT distance="950" swimtime="00:14:14.72" />
                    <SPLIT distance="1000" swimtime="00:14:59.65" />
                    <SPLIT distance="1050" swimtime="00:15:44.11" />
                    <SPLIT distance="1100" swimtime="00:16:29.01" />
                    <SPLIT distance="1150" swimtime="00:17:13.12" />
                    <SPLIT distance="1200" swimtime="00:17:57.69" />
                    <SPLIT distance="1250" swimtime="00:18:42.38" />
                    <SPLIT distance="1300" swimtime="00:19:27.05" />
                    <SPLIT distance="1350" swimtime="00:20:11.99" />
                    <SPLIT distance="1400" swimtime="00:20:56.64" />
                    <SPLIT distance="1450" swimtime="00:21:40.61" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Oliveira Martini" birthdate="2008-10-31" gender="M" nation="BRA" license="406953" swrid="5717285" athleteid="3218" externalid="406953">
              <RESULTS>
                <RESULT eventid="1120" points="271" swimtime="00:02:37.45" resultid="3219" heatid="5153" lane="2" entrytime="00:02:33.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.40" />
                    <SPLIT distance="100" swimtime="00:01:14.39" />
                    <SPLIT distance="150" swimtime="00:01:56.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Maria Romanelli" birthdate="2011-04-18" gender="F" nation="BRA" license="378335" swrid="5588803" athleteid="3196" externalid="378335">
              <RESULTS>
                <RESULT eventid="1096" points="385" swimtime="00:00:32.43" resultid="3197" heatid="5099" lane="2" entrytime="00:00:31.52" entrycourse="LCM" />
                <RESULT eventid="1159" status="DNS" swimtime="00:00:00.00" resultid="3198" heatid="5203" lane="6" entrytime="00:01:10.02" entrycourse="LCM" />
                <RESULT eventid="1215" status="DNS" swimtime="00:00:00.00" resultid="3199" heatid="5292" lane="3" entrytime="00:00:41.78" entrycourse="LCM" />
                <RESULT eventid="1305" status="DNS" swimtime="00:00:00.00" resultid="3200" heatid="5374" lane="1" entrytime="00:00:47.90" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Flavia" lastname="Scheffler Souza" birthdate="2010-09-14" gender="F" nation="BRA" license="417278" athleteid="3232" externalid="417278">
              <RESULTS>
                <RESULT eventid="1096" points="375" swimtime="00:00:32.72" resultid="3233" heatid="5095" lane="3" />
                <RESULT eventid="1112" status="DNS" swimtime="00:00:00.00" resultid="3234" heatid="5138" lane="8" />
                <RESULT eventid="1159" points="359" swimtime="00:01:12.71" resultid="3235" heatid="5201" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Milena" lastname="Vieira De Macedo Brasil" birthdate="2009-12-19" gender="F" nation="BRA" license="344143" swrid="5622311" athleteid="3186" externalid="344143">
              <RESULTS>
                <RESULT eventid="1096" points="424" swimtime="00:00:31.41" resultid="3187" heatid="5102" lane="2" entrytime="00:00:32.05" entrycourse="LCM" />
                <RESULT eventid="1143" points="280" swimtime="00:03:12.77" resultid="3188" heatid="5189" lane="2" entrytime="00:03:15.06" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.20" />
                    <SPLIT distance="100" swimtime="00:01:35.20" />
                    <SPLIT distance="150" swimtime="00:02:30.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="348" swimtime="00:00:41.42" resultid="3189" heatid="5374" lane="2" entrytime="00:00:45.28" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vicente" lastname="Bileski" birthdate="2011-06-29" gender="M" nation="BRA" license="406950" swrid="5717248" athleteid="3212" externalid="406950">
              <RESULTS>
                <RESULT eventid="1104" points="260" swimtime="00:00:32.76" resultid="3213" heatid="5116" lane="7" entrytime="00:00:33.88" entrycourse="LCM" />
                <RESULT eventid="1120" points="224" swimtime="00:02:47.71" resultid="3214" heatid="5148" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.02" />
                    <SPLIT distance="100" swimtime="00:01:18.96" />
                    <SPLIT distance="150" swimtime="00:02:04.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="209" swimtime="00:03:11.82" resultid="3215" heatid="5193" lane="2" entrytime="00:03:15.62" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.31" />
                    <SPLIT distance="100" swimtime="00:01:30.02" />
                    <SPLIT distance="150" swimtime="00:02:27.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="244" swimtime="00:01:14.97" resultid="3216" heatid="5218" lane="6" entrytime="00:01:22.57" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="242" swimtime="00:00:35.73" resultid="3217" heatid="5331" lane="7" entrytime="00:00:36.48" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="13025" nation="BRA" region="PR" clubid="3035" swrid="93779" name="Instituto Desportos Aquáticos De Foz Do Iguaçu" shortname="Cataratas Natação">
          <ATHLETES>
            <ATHLETE firstname="Ysadora" lastname="Bertoldo" birthdate="2010-04-09" gender="F" nation="BRA" license="376444" swrid="5588553" athleteid="3134" externalid="376444" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1064" points="422" swimtime="00:05:13.59" resultid="3135" heatid="5050" lane="6" entrytime="00:05:10.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.67" />
                    <SPLIT distance="100" swimtime="00:01:14.10" />
                    <SPLIT distance="150" swimtime="00:01:54.32" />
                    <SPLIT distance="200" swimtime="00:02:34.85" />
                    <SPLIT distance="250" swimtime="00:03:15.02" />
                    <SPLIT distance="300" swimtime="00:03:54.89" />
                    <SPLIT distance="350" swimtime="00:04:35.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" points="299" swimtime="00:01:22.95" resultid="3136" heatid="5159" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="423" swimtime="00:02:30.23" resultid="3137" heatid="5140" lane="1" entrytime="00:02:28.99" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.28" />
                    <SPLIT distance="100" swimtime="00:01:12.58" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" status="DNS" swimtime="00:00:00.00" resultid="3138" heatid="5271" lane="6" entrytime="00:10:33.44" entrycourse="LCM" />
                <RESULT eventid="1215" points="380" swimtime="00:00:37.08" resultid="3139" heatid="5291" lane="8" />
                <RESULT eventid="1279" points="416" swimtime="00:20:32.46" resultid="3140" heatid="5350" lane="2" entrytime="00:20:10.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.32" />
                    <SPLIT distance="100" swimtime="00:01:15.76" />
                    <SPLIT distance="150" swimtime="00:01:56.47" />
                    <SPLIT distance="200" swimtime="00:02:37.99" />
                    <SPLIT distance="250" swimtime="00:03:18.89" />
                    <SPLIT distance="300" swimtime="00:04:00.94" />
                    <SPLIT distance="350" swimtime="00:04:41.81" />
                    <SPLIT distance="400" swimtime="00:05:23.38" />
                    <SPLIT distance="450" swimtime="00:06:04.71" />
                    <SPLIT distance="500" swimtime="00:06:46.42" />
                    <SPLIT distance="550" swimtime="00:07:27.17" />
                    <SPLIT distance="600" swimtime="00:08:08.73" />
                    <SPLIT distance="650" swimtime="00:08:50.34" />
                    <SPLIT distance="700" swimtime="00:09:31.77" />
                    <SPLIT distance="750" swimtime="00:10:12.93" />
                    <SPLIT distance="800" swimtime="00:10:54.89" />
                    <SPLIT distance="850" swimtime="00:11:36.79" />
                    <SPLIT distance="900" swimtime="00:12:18.63" />
                    <SPLIT distance="1000" swimtime="00:13:42.41" />
                    <SPLIT distance="1050" swimtime="00:14:24.24" />
                    <SPLIT distance="1150" swimtime="00:15:49.22" />
                    <SPLIT distance="1200" swimtime="00:16:31.16" />
                    <SPLIT distance="1250" swimtime="00:17:13.21" />
                    <SPLIT distance="1300" swimtime="00:17:54.71" />
                    <SPLIT distance="1350" swimtime="00:18:35.01" />
                    <SPLIT distance="1400" swimtime="00:19:15.68" />
                    <SPLIT distance="1450" swimtime="00:19:54.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Gabriel Dreher" birthdate="2011-12-05" gender="M" nation="BRA" license="403148" swrid="5676302" athleteid="3127" externalid="403148" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1104" points="201" swimtime="00:00:35.68" resultid="3128" heatid="5115" lane="6" entrytime="00:00:36.27" entrycourse="LCM" />
                <RESULT eventid="1120" points="196" swimtime="00:02:55.44" resultid="3129" heatid="5148" lane="4" entrytime="00:02:54.91" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                    <SPLIT distance="100" swimtime="00:01:23.20" />
                    <SPLIT distance="150" swimtime="00:02:11.87" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="220" swimtime="00:01:25.36" resultid="3130" heatid="5255" lane="5" entrytime="00:01:30.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="204" swimtime="00:00:39.94" resultid="3131" heatid="5283" lane="6" entrytime="00:00:47.17" entrycourse="LCM" />
                <RESULT eventid="1251" points="182" swimtime="00:03:41.40" resultid="3132" heatid="5315" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.71" />
                    <SPLIT distance="100" swimtime="00:01:46.31" />
                    <SPLIT distance="150" swimtime="00:02:44.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="180" swimtime="00:00:45.90" resultid="3133" heatid="5365" lane="4" entrytime="00:00:53.11" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinicius" lastname="Monteiro Viebrantz" birthdate="2003-01-09" gender="M" nation="BRA" license="291175" swrid="5600219" athleteid="3047" externalid="291175">
              <RESULTS>
                <RESULT eventid="1104" points="596" swimtime="00:00:24.84" resultid="3048" heatid="5130" lane="5" entrytime="00:00:23.44" entrycourse="LCM" />
                <RESULT eventid="1167" status="DNS" swimtime="00:00:00.00" resultid="3049" heatid="5233" lane="5" entrytime="00:00:50.36" entrycourse="LCM" />
                <RESULT eventid="1267" status="DNS" swimtime="00:00:00.00" resultid="3050" heatid="5338" lane="2" entrytime="00:00:26.24" entrycourse="LCM" />
                <RESULT eventid="2383" swimtime="00:00:00.00" resultid="5988" entrytime="00:00:24.84" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Bailke" birthdate="2007-05-04" gender="M" nation="BRA" license="370566" swrid="5596869" athleteid="3093" externalid="370566" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1072" points="349" swimtime="00:05:12.34" resultid="3094" heatid="5064" lane="8" entrytime="00:05:04.65" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.12" />
                    <SPLIT distance="100" swimtime="00:01:07.75" />
                    <SPLIT distance="150" swimtime="00:01:45.40" />
                    <SPLIT distance="200" swimtime="00:02:26.46" />
                    <SPLIT distance="250" swimtime="00:03:07.29" />
                    <SPLIT distance="300" swimtime="00:03:50.44" />
                    <SPLIT distance="350" swimtime="00:04:31.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="335" swimtime="00:01:11.19" resultid="3095" heatid="5176" lane="5" entrytime="00:01:13.61" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="362" swimtime="00:10:34.19" resultid="3096" heatid="5298" lane="2" entrytime="00:10:44.50" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.72" />
                    <SPLIT distance="100" swimtime="00:01:10.93" />
                    <SPLIT distance="150" swimtime="00:01:50.11" />
                    <SPLIT distance="200" swimtime="00:02:30.21" />
                    <SPLIT distance="250" swimtime="00:03:11.03" />
                    <SPLIT distance="300" swimtime="00:03:53.30" />
                    <SPLIT distance="350" swimtime="00:04:34.43" />
                    <SPLIT distance="400" swimtime="00:05:16.02" />
                    <SPLIT distance="450" swimtime="00:05:57.99" />
                    <SPLIT distance="500" swimtime="00:06:39.31" />
                    <SPLIT distance="550" swimtime="00:07:19.82" />
                    <SPLIT distance="600" swimtime="00:08:00.66" />
                    <SPLIT distance="650" swimtime="00:08:39.80" />
                    <SPLIT distance="700" swimtime="00:09:20.12" />
                    <SPLIT distance="750" swimtime="00:09:59.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="356" swimtime="00:00:31.42" resultid="3097" heatid="5328" lane="5" />
                <RESULT eventid="1312" points="343" swimtime="00:20:43.86" resultid="3098" heatid="5379" lane="7" entrytime="00:20:31.34" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.94" />
                    <SPLIT distance="100" swimtime="00:01:14.02" />
                    <SPLIT distance="150" swimtime="00:01:54.50" />
                    <SPLIT distance="200" swimtime="00:02:35.91" />
                    <SPLIT distance="250" swimtime="00:03:16.27" />
                    <SPLIT distance="300" swimtime="00:03:57.58" />
                    <SPLIT distance="350" swimtime="00:04:40.08" />
                    <SPLIT distance="400" swimtime="00:05:21.28" />
                    <SPLIT distance="450" swimtime="00:06:03.52" />
                    <SPLIT distance="500" swimtime="00:06:45.94" />
                    <SPLIT distance="550" swimtime="00:07:29.72" />
                    <SPLIT distance="600" swimtime="00:08:11.54" />
                    <SPLIT distance="650" swimtime="00:08:53.43" />
                    <SPLIT distance="700" swimtime="00:09:35.97" />
                    <SPLIT distance="750" swimtime="00:10:19.45" />
                    <SPLIT distance="800" swimtime="00:11:01.41" />
                    <SPLIT distance="850" swimtime="00:11:44.58" />
                    <SPLIT distance="900" swimtime="00:12:27.62" />
                    <SPLIT distance="950" swimtime="00:13:08.44" />
                    <SPLIT distance="1000" swimtime="00:13:50.38" />
                    <SPLIT distance="1050" swimtime="00:14:32.24" />
                    <SPLIT distance="1100" swimtime="00:15:14.50" />
                    <SPLIT distance="1150" swimtime="00:15:56.28" />
                    <SPLIT distance="1200" swimtime="00:16:37.99" />
                    <SPLIT distance="1250" swimtime="00:17:22.40" />
                    <SPLIT distance="1300" swimtime="00:18:04.18" />
                    <SPLIT distance="1350" swimtime="00:18:46.45" />
                    <SPLIT distance="1400" swimtime="00:19:28.26" />
                    <SPLIT distance="1450" swimtime="00:20:07.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Rogge" birthdate="2008-09-02" gender="M" nation="BRA" license="383387" swrid="4883279" athleteid="3051" externalid="383387" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1104" points="548" swimtime="00:00:25.55" resultid="3052" heatid="5125" lane="6" entrytime="00:00:26.20" entrycourse="LCM" />
                <RESULT eventid="1120" points="418" swimtime="00:02:16.34" resultid="3053" heatid="5154" lane="6" entrytime="00:02:18.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.94" />
                    <SPLIT distance="100" swimtime="00:01:06.71" />
                    <SPLIT distance="150" swimtime="00:01:40.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="347" swimtime="00:02:42.21" resultid="3054" heatid="5196" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.38" />
                    <SPLIT distance="100" swimtime="00:01:15.31" />
                    <SPLIT distance="150" swimtime="00:02:05.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="565" swimtime="00:00:56.66" resultid="3055" heatid="5230" lane="8" entrytime="00:00:56.86" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="412" swimtime="00:00:31.64" resultid="3056" heatid="5286" lane="6" entrytime="00:00:31.79" entrycourse="LCM" />
                <RESULT eventid="1267" points="393" swimtime="00:00:30.40" resultid="3057" heatid="5333" lane="5" entrytime="00:00:30.85" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Mayumi" lastname="Napole" birthdate="2010-02-01" gender="F" nation="BRA" license="376446" swrid="5596918" athleteid="3155" externalid="376446" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1096" points="409" swimtime="00:00:31.80" resultid="3156" heatid="5099" lane="1" entrytime="00:00:31.70" entrycourse="LCM" />
                <RESULT eventid="1143" points="319" swimtime="00:03:04.39" resultid="3157" heatid="5187" lane="8" entrytime="00:03:07.90" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.78" />
                    <SPLIT distance="100" swimtime="00:01:24.34" />
                    <SPLIT distance="150" swimtime="00:02:18.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="325" swimtime="00:01:23.35" resultid="3158" heatid="5243" lane="8" entrytime="00:01:22.49" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="361" swimtime="00:00:37.72" resultid="3159" heatid="5290" lane="3" />
                <RESULT eventid="1275" points="323" swimtime="00:02:59.37" resultid="3160" heatid="5339" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.03" />
                    <SPLIT distance="100" swimtime="00:01:29.90" />
                    <SPLIT distance="150" swimtime="00:02:15.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="316" swimtime="00:00:42.80" resultid="3161" heatid="5372" lane="6" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Marques Petry" birthdate="2008-01-08" gender="M" nation="BRA" license="392351" swrid="4711489" athleteid="3106" externalid="392351" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1072" points="441" swimtime="00:04:48.99" resultid="3107" heatid="5061" lane="2" entrytime="00:04:49.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.07" />
                    <SPLIT distance="100" swimtime="00:01:07.10" />
                    <SPLIT distance="150" swimtime="00:01:43.70" />
                    <SPLIT distance="200" swimtime="00:02:21.41" />
                    <SPLIT distance="250" swimtime="00:02:58.23" />
                    <SPLIT distance="300" swimtime="00:03:36.12" />
                    <SPLIT distance="350" swimtime="00:04:13.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="400" swimtime="00:00:28.37" resultid="3108" heatid="5121" lane="3" entrytime="00:00:30.91" entrycourse="LCM" />
                <RESULT eventid="1135" points="267" swimtime="00:01:16.75" resultid="3109" heatid="5172" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="408" swimtime="00:01:03.13" resultid="3110" heatid="5225" lane="4" entrytime="00:01:04.38" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="391" swimtime="00:10:17.98" resultid="3111" heatid="5299" lane="7" entrytime="00:10:04.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.11" />
                    <SPLIT distance="100" swimtime="00:01:09.62" />
                    <SPLIT distance="150" swimtime="00:01:47.90" />
                    <SPLIT distance="200" swimtime="00:02:26.71" />
                    <SPLIT distance="250" swimtime="00:03:06.35" />
                    <SPLIT distance="300" swimtime="00:03:46.22" />
                    <SPLIT distance="350" swimtime="00:04:25.26" />
                    <SPLIT distance="400" swimtime="00:05:04.20" />
                    <SPLIT distance="450" swimtime="00:05:42.96" />
                    <SPLIT distance="500" swimtime="00:06:22.19" />
                    <SPLIT distance="550" swimtime="00:07:01.62" />
                    <SPLIT distance="600" swimtime="00:07:41.26" />
                    <SPLIT distance="650" swimtime="00:08:20.23" />
                    <SPLIT distance="700" swimtime="00:08:58.72" />
                    <SPLIT distance="750" swimtime="00:09:37.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="407" swimtime="00:19:34.89" resultid="3112" heatid="5379" lane="4" entrytime="00:19:31.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.02" />
                    <SPLIT distance="100" swimtime="00:01:12.34" />
                    <SPLIT distance="150" swimtime="00:01:52.11" />
                    <SPLIT distance="200" swimtime="00:02:32.91" />
                    <SPLIT distance="250" swimtime="00:03:11.83" />
                    <SPLIT distance="300" swimtime="00:03:51.91" />
                    <SPLIT distance="350" swimtime="00:04:31.15" />
                    <SPLIT distance="400" swimtime="00:05:12.27" />
                    <SPLIT distance="450" swimtime="00:05:52.62" />
                    <SPLIT distance="500" swimtime="00:06:33.99" />
                    <SPLIT distance="550" swimtime="00:07:13.41" />
                    <SPLIT distance="600" swimtime="00:07:53.46" />
                    <SPLIT distance="650" swimtime="00:08:32.21" />
                    <SPLIT distance="700" swimtime="00:09:11.61" />
                    <SPLIT distance="750" swimtime="00:09:51.14" />
                    <SPLIT distance="800" swimtime="00:10:31.35" />
                    <SPLIT distance="850" swimtime="00:11:10.30" />
                    <SPLIT distance="900" swimtime="00:11:49.96" />
                    <SPLIT distance="950" swimtime="00:12:29.74" />
                    <SPLIT distance="1000" swimtime="00:13:09.55" />
                    <SPLIT distance="1050" swimtime="00:13:48.91" />
                    <SPLIT distance="1100" swimtime="00:14:29.30" />
                    <SPLIT distance="1150" swimtime="00:15:09.07" />
                    <SPLIT distance="1200" swimtime="00:15:47.90" />
                    <SPLIT distance="1250" swimtime="00:16:27.03" />
                    <SPLIT distance="1300" swimtime="00:17:06.64" />
                    <SPLIT distance="1350" swimtime="00:17:44.13" />
                    <SPLIT distance="1400" swimtime="00:18:22.50" />
                    <SPLIT distance="1450" swimtime="00:18:58.83" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovanna" lastname="Mattiello" birthdate="2009-04-11" gender="F" nation="BRA" license="367011" swrid="5596914" athleteid="3099" externalid="367011" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1096" points="455" swimtime="00:00:30.68" resultid="3100" heatid="5103" lane="8" entrytime="00:00:30.58" entrycourse="LCM" />
                <RESULT eventid="1112" points="422" swimtime="00:02:30.37" resultid="3101" heatid="5143" lane="4" entrytime="00:02:26.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.22" />
                    <SPLIT distance="100" swimtime="00:01:11.51" />
                    <SPLIT distance="150" swimtime="00:01:51.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="352" swimtime="00:01:21.13" resultid="3102" heatid="5245" lane="4" entrytime="00:01:24.47" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="433" swimtime="00:01:08.33" resultid="3103" heatid="5207" lane="7" entrytime="00:01:08.35" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="346" swimtime="00:00:38.26" resultid="3104" heatid="5293" lane="2" entrytime="00:00:38.92" entrycourse="LCM" />
                <RESULT eventid="1275" points="338" swimtime="00:02:56.65" resultid="3105" heatid="5340" lane="5" entrytime="00:02:59.94" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.62" />
                    <SPLIT distance="100" swimtime="00:01:27.29" />
                    <SPLIT distance="150" swimtime="00:02:13.98" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Natalia" lastname="Sermidi" birthdate="2005-06-15" gender="F" nation="BRA" license="283035" swrid="5596938" athleteid="3043" externalid="283035" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1259" points="373" swimtime="00:00:33.93" resultid="3044" heatid="5326" lane="8" entrytime="00:00:33.06" entrycourse="LCM" />
                <RESULT eventid="1275" points="318" swimtime="00:03:00.28" resultid="3045" heatid="5339" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.50" />
                    <SPLIT distance="100" swimtime="00:01:28.46" />
                    <SPLIT distance="150" swimtime="00:02:14.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="223" swimtime="00:00:48.05" resultid="3046" heatid="5372" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Leticia Sbardelatti" birthdate="2011-07-28" gender="F" nation="BRA" license="403147" swrid="5676303" athleteid="3120" externalid="403147" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1064" points="200" swimtime="00:06:41.98" resultid="3121" heatid="5048" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.07" />
                    <SPLIT distance="100" swimtime="00:01:30.86" />
                    <SPLIT distance="150" swimtime="00:02:22.68" />
                    <SPLIT distance="200" swimtime="00:03:13.83" />
                    <SPLIT distance="250" swimtime="00:04:06.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="264" swimtime="00:00:36.77" resultid="3122" heatid="5096" lane="6" entrytime="00:00:37.32" entrycourse="LCM" />
                <RESULT eventid="1112" points="215" swimtime="00:03:08.11" resultid="3123" heatid="5138" lane="1" entrytime="00:03:16.81" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.70" />
                    <SPLIT distance="100" swimtime="00:01:28.78" />
                    <SPLIT distance="150" swimtime="00:02:18.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="250" swimtime="00:01:22.08" resultid="3124" heatid="5201" lane="7" entrytime="00:01:26.04" entrycourse="LCM" />
                <RESULT eventid="1215" points="183" swimtime="00:00:47.29" resultid="3125" heatid="5291" lane="1" entrytime="00:00:53.60" entrycourse="LCM" />
                <RESULT eventid="1305" points="227" swimtime="00:00:47.77" resultid="3126" heatid="5374" lane="8" entrytime="00:00:51.16" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Christopher" lastname="De Araujo" birthdate="2008-08-09" gender="M" nation="BRA" license="366376" swrid="5596884" athleteid="3086" externalid="366376" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1072" points="550" swimtime="00:04:28.47" resultid="3087" heatid="5062" lane="1" entrytime="00:04:33.48" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.22" />
                    <SPLIT distance="100" swimtime="00:01:02.08" />
                    <SPLIT distance="150" swimtime="00:01:35.93" />
                    <SPLIT distance="200" swimtime="00:02:10.74" />
                    <SPLIT distance="250" swimtime="00:02:44.49" />
                    <SPLIT distance="300" swimtime="00:03:19.56" />
                    <SPLIT distance="350" swimtime="00:03:54.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="452" swimtime="00:02:28.52" resultid="3088" heatid="5198" lane="8" entrytime="00:02:25.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.92" />
                    <SPLIT distance="100" swimtime="00:01:09.02" />
                    <SPLIT distance="150" swimtime="00:01:54.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="558" swimtime="00:00:56.91" resultid="3089" heatid="5228" lane="3" entrytime="00:00:58.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="493" swimtime="00:09:32.14" resultid="3090" heatid="5300" lane="2" entrytime="00:09:13.39" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                    <SPLIT distance="100" swimtime="00:01:04.73" />
                    <SPLIT distance="150" swimtime="00:01:39.01" />
                    <SPLIT distance="200" swimtime="00:02:14.21" />
                    <SPLIT distance="250" swimtime="00:02:50.21" />
                    <SPLIT distance="300" swimtime="00:03:26.71" />
                    <SPLIT distance="350" swimtime="00:04:03.70" />
                    <SPLIT distance="400" swimtime="00:04:40.43" />
                    <SPLIT distance="450" swimtime="00:05:17.13" />
                    <SPLIT distance="500" swimtime="00:05:53.76" />
                    <SPLIT distance="550" swimtime="00:06:31.29" />
                    <SPLIT distance="600" swimtime="00:07:07.67" />
                    <SPLIT distance="650" swimtime="00:07:44.69" />
                    <SPLIT distance="700" swimtime="00:08:21.43" />
                    <SPLIT distance="750" swimtime="00:08:57.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="374" swimtime="00:02:54.12" resultid="3091" heatid="5319" lane="6" entrytime="00:02:41.43" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.83" />
                    <SPLIT distance="100" swimtime="00:01:23.07" />
                    <SPLIT distance="150" swimtime="00:02:10.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="487" swimtime="00:18:26.96" resultid="3092" heatid="5380" lane="3" entrytime="00:17:44.18" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.59" />
                    <SPLIT distance="100" swimtime="00:01:04.01" />
                    <SPLIT distance="150" swimtime="00:01:39.52" />
                    <SPLIT distance="200" swimtime="00:02:15.16" />
                    <SPLIT distance="250" swimtime="00:02:51.58" />
                    <SPLIT distance="300" swimtime="00:03:28.53" />
                    <SPLIT distance="350" swimtime="00:04:05.22" />
                    <SPLIT distance="400" swimtime="00:04:42.59" />
                    <SPLIT distance="450" swimtime="00:05:20.63" />
                    <SPLIT distance="500" swimtime="00:05:57.95" />
                    <SPLIT distance="550" swimtime="00:06:34.83" />
                    <SPLIT distance="600" swimtime="00:07:12.38" />
                    <SPLIT distance="650" swimtime="00:07:48.99" />
                    <SPLIT distance="700" swimtime="00:08:26.54" />
                    <SPLIT distance="750" swimtime="00:09:04.39" />
                    <SPLIT distance="800" swimtime="00:09:41.25" />
                    <SPLIT distance="850" swimtime="00:10:18.53" />
                    <SPLIT distance="900" swimtime="00:10:56.63" />
                    <SPLIT distance="950" swimtime="00:11:34.39" />
                    <SPLIT distance="1000" swimtime="00:12:11.74" />
                    <SPLIT distance="1050" swimtime="00:12:49.55" />
                    <SPLIT distance="1100" swimtime="00:13:27.19" />
                    <SPLIT distance="1150" swimtime="00:14:05.06" />
                    <SPLIT distance="1200" swimtime="00:14:42.51" />
                    <SPLIT distance="1250" swimtime="00:15:20.23" />
                    <SPLIT distance="1300" swimtime="00:15:57.61" />
                    <SPLIT distance="1350" swimtime="00:16:35.06" />
                    <SPLIT distance="1400" swimtime="00:17:12.93" />
                    <SPLIT distance="1450" swimtime="00:17:50.48" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Carvalho Carelli" birthdate="2011-10-15" gender="M" nation="BRA" license="403146" swrid="5676300" athleteid="3141" externalid="403146" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1104" points="358" swimtime="00:00:29.43" resultid="3142" heatid="5114" lane="6" />
                <RESULT eventid="1135" points="323" swimtime="00:01:12.07" resultid="3143" heatid="5170" lane="3" entrytime="00:01:16.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="396" swimtime="00:02:18.84" resultid="3144" heatid="5150" lane="4" entrytime="00:02:23.60" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                    <SPLIT distance="100" swimtime="00:01:07.36" />
                    <SPLIT distance="150" swimtime="00:01:43.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="393" swimtime="00:01:03.95" resultid="3145" heatid="5221" lane="8" entrytime="00:01:06.36" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="364" swimtime="00:00:31.18" resultid="3146" heatid="5327" lane="5" />
                <RESULT eventid="1293" status="DNS" swimtime="00:00:00.00" resultid="3147" heatid="5357" lane="4" entrytime="00:03:06.20" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Faisal" lastname="Basem Ghotme" birthdate="2010-12-18" gender="M" nation="BRA" license="390809" swrid="5596871" athleteid="3162" externalid="390809" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1104" points="507" swimtime="00:00:26.22" resultid="3163" heatid="5120" lane="7" entrytime="00:00:27.26" entrycourse="LCM" />
                <RESULT eventid="1120" points="394" swimtime="00:02:19.11" resultid="3164" heatid="5149" lane="1" entrytime="00:02:37.79" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.77" />
                    <SPLIT distance="100" swimtime="00:01:06.04" />
                    <SPLIT distance="150" swimtime="00:01:43.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="429" swimtime="00:01:08.41" resultid="3165" heatid="5258" lane="8" entrytime="00:01:08.37" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="500" swimtime="00:00:59.03" resultid="3166" heatid="5222" lane="5" entrytime="00:01:01.04" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="431" swimtime="00:00:31.16" resultid="3167" heatid="5286" lane="8" entrytime="00:00:32.65" entrycourse="LCM" />
                <RESULT eventid="1277" points="378" swimtime="00:02:34.66" resultid="3168" heatid="5347" lane="7" entrytime="00:02:26.72" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.28" />
                    <SPLIT distance="100" swimtime="00:01:14.20" />
                    <SPLIT distance="150" swimtime="00:01:54.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Luiz Martinazzo" birthdate="2006-05-16" gender="M" nation="BRA" license="345593" swrid="5596910" athleteid="3079" externalid="345593" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1072" points="462" swimtime="00:04:44.66" resultid="3080" heatid="5064" lane="6" entrytime="00:04:33.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.41" />
                    <SPLIT distance="100" swimtime="00:01:02.12" />
                    <SPLIT distance="150" swimtime="00:01:37.16" />
                    <SPLIT distance="200" swimtime="00:02:13.04" />
                    <SPLIT distance="250" swimtime="00:02:50.66" />
                    <SPLIT distance="300" swimtime="00:03:28.66" />
                    <SPLIT distance="350" swimtime="00:04:07.43" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="493" swimtime="00:02:09.07" resultid="3081" heatid="5158" lane="7" entrytime="00:02:06.76" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.00" />
                    <SPLIT distance="100" swimtime="00:01:01.54" />
                    <SPLIT distance="150" swimtime="00:01:35.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="452" swimtime="00:01:07.23" resultid="3082" heatid="5262" lane="4" entrytime="00:01:06.85" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.72" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="459" swimtime="00:09:46.06" resultid="3083" heatid="5299" lane="4" entrytime="00:09:39.07" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.42" />
                    <SPLIT distance="100" swimtime="00:01:04.99" />
                    <SPLIT distance="150" swimtime="00:01:41.18" />
                    <SPLIT distance="200" swimtime="00:02:17.39" />
                    <SPLIT distance="250" swimtime="00:02:54.32" />
                    <SPLIT distance="300" swimtime="00:03:31.45" />
                    <SPLIT distance="350" swimtime="00:04:09.05" />
                    <SPLIT distance="400" swimtime="00:04:46.95" />
                    <SPLIT distance="450" swimtime="00:05:24.82" />
                    <SPLIT distance="500" swimtime="00:06:02.77" />
                    <SPLIT distance="550" swimtime="00:06:40.96" />
                    <SPLIT distance="600" swimtime="00:07:18.90" />
                    <SPLIT distance="650" swimtime="00:07:56.13" />
                    <SPLIT distance="700" swimtime="00:08:33.95" />
                    <SPLIT distance="750" swimtime="00:09:10.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="433" swimtime="00:02:27.91" resultid="3084" heatid="5346" lane="4" entrytime="00:02:30.11" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.81" />
                    <SPLIT distance="100" swimtime="00:01:10.59" />
                    <SPLIT distance="150" swimtime="00:01:49.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1312" points="445" swimtime="00:19:00.88" resultid="3085" heatid="5380" lane="7" entrytime="00:18:43.29" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                    <SPLIT distance="100" swimtime="00:01:06.04" />
                    <SPLIT distance="150" swimtime="00:01:43.17" />
                    <SPLIT distance="200" swimtime="00:02:20.77" />
                    <SPLIT distance="250" swimtime="00:02:58.89" />
                    <SPLIT distance="300" swimtime="00:03:36.93" />
                    <SPLIT distance="350" swimtime="00:04:15.23" />
                    <SPLIT distance="400" swimtime="00:04:53.83" />
                    <SPLIT distance="450" swimtime="00:05:33.06" />
                    <SPLIT distance="500" swimtime="00:06:12.18" />
                    <SPLIT distance="550" swimtime="00:06:51.06" />
                    <SPLIT distance="600" swimtime="00:07:30.37" />
                    <SPLIT distance="650" swimtime="00:08:08.86" />
                    <SPLIT distance="700" swimtime="00:08:47.67" />
                    <SPLIT distance="750" swimtime="00:09:26.41" />
                    <SPLIT distance="800" swimtime="00:10:05.17" />
                    <SPLIT distance="850" swimtime="00:10:43.66" />
                    <SPLIT distance="900" swimtime="00:11:22.90" />
                    <SPLIT distance="950" swimtime="00:12:01.44" />
                    <SPLIT distance="1000" swimtime="00:12:40.10" />
                    <SPLIT distance="1050" swimtime="00:13:18.94" />
                    <SPLIT distance="1100" swimtime="00:13:58.15" />
                    <SPLIT distance="1150" swimtime="00:14:36.72" />
                    <SPLIT distance="1200" swimtime="00:15:14.89" />
                    <SPLIT distance="1250" swimtime="00:15:53.22" />
                    <SPLIT distance="1300" swimtime="00:16:31.11" />
                    <SPLIT distance="1350" swimtime="00:17:08.97" />
                    <SPLIT distance="1400" swimtime="00:17:46.93" />
                    <SPLIT distance="1450" swimtime="00:18:24.25" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Resende Ames" birthdate="2006-02-10" gender="M" nation="BRA" license="365657" swrid="5596931" athleteid="3065" externalid="365657" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1072" points="518" swimtime="00:04:33.88" resultid="3066" heatid="5063" lane="4">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:01.86" />
                    <SPLIT distance="150" swimtime="00:01:35.98" />
                    <SPLIT distance="200" swimtime="00:02:10.38" />
                    <SPLIT distance="250" swimtime="00:02:46.01" />
                    <SPLIT distance="300" swimtime="00:03:21.71" />
                    <SPLIT distance="350" swimtime="00:03:58.44" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1135" points="571" swimtime="00:00:59.60" resultid="3067" heatid="5178" lane="8" entrytime="00:00:59.44" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="422" swimtime="00:01:08.76" resultid="3068" heatid="5262" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.31" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1198" points="464" swimtime="00:05:13.04" resultid="3069" heatid="5275" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.30" />
                    <SPLIT distance="100" swimtime="00:01:03.22" />
                    <SPLIT distance="150" swimtime="00:01:44.18" />
                    <SPLIT distance="200" swimtime="00:02:23.21" />
                    <SPLIT distance="250" swimtime="00:03:13.90" />
                    <SPLIT distance="300" swimtime="00:04:04.29" />
                    <SPLIT distance="350" swimtime="00:04:38.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1277" points="446" swimtime="00:02:26.39" resultid="3070" heatid="5347" lane="5" entrytime="00:02:24.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.57" />
                    <SPLIT distance="100" swimtime="00:01:12.82" />
                    <SPLIT distance="150" swimtime="00:01:50.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1293" points="465" swimtime="00:02:22.33" resultid="3071" heatid="5360" lane="5" entrytime="00:02:13.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.06" />
                    <SPLIT distance="100" swimtime="00:01:04.95" />
                    <SPLIT distance="150" swimtime="00:01:41.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Victor Oliveira" birthdate="2003-07-16" gender="M" nation="BRA" license="295723" swrid="5596944" athleteid="3058" externalid="295723" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1104" points="527" swimtime="00:00:25.88" resultid="3059" heatid="5128" lane="5" entrytime="00:00:26.26" entrycourse="LCM" />
                <RESULT eventid="1135" points="536" swimtime="00:01:00.86" resultid="3060" heatid="5177" lane="4" entrytime="00:00:59.84" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="525" swimtime="00:01:03.95" resultid="3061" heatid="5263" lane="7" entrytime="00:01:02.33" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.75" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="504" swimtime="00:00:29.58" resultid="3062" heatid="5288" lane="1" entrytime="00:00:28.82" entrycourse="LCM" />
                <RESULT eventid="1267" points="528" swimtime="00:00:27.54" resultid="3063" heatid="5337" lane="5" entrytime="00:00:26.85" entrycourse="LCM" />
                <RESULT eventid="1277" points="476" swimtime="00:02:23.26" resultid="3064" heatid="5348" lane="1" entrytime="00:02:20.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.95" />
                    <SPLIT distance="100" swimtime="00:01:09.45" />
                    <SPLIT distance="150" swimtime="00:01:46.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="2359" points="529" swimtime="00:01:03.80" resultid="6448" heatid="6423" lane="8" entrytime="00:01:03.95">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Targat Pinheiro" birthdate="2008-09-04" gender="F" nation="BRA" license="331610" swrid="5596894" athleteid="3036" externalid="331610" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1064" points="437" swimtime="00:05:09.96" resultid="3037" heatid="5053" lane="7" entrytime="00:05:20.52" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                    <SPLIT distance="100" swimtime="00:01:10.72" />
                    <SPLIT distance="150" swimtime="00:01:49.37" />
                    <SPLIT distance="200" swimtime="00:02:30.01" />
                    <SPLIT distance="250" swimtime="00:03:10.23" />
                    <SPLIT distance="300" swimtime="00:03:51.16" />
                    <SPLIT distance="350" swimtime="00:04:30.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1128" points="443" swimtime="00:01:12.77" resultid="3038" heatid="5161" lane="5" entrytime="00:01:12.83" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.14" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="468" swimtime="00:02:25.31" resultid="3039" heatid="5142" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.37" />
                    <SPLIT distance="100" swimtime="00:01:10.65" />
                    <SPLIT distance="150" swimtime="00:01:48.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1190" points="421" swimtime="00:10:46.74" resultid="3040" heatid="5272" lane="3" entrytime="00:10:35.98" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.83" />
                    <SPLIT distance="100" swimtime="00:01:11.19" />
                    <SPLIT distance="150" swimtime="00:01:51.69" />
                    <SPLIT distance="200" swimtime="00:02:31.92" />
                    <SPLIT distance="250" swimtime="00:03:12.97" />
                    <SPLIT distance="300" swimtime="00:03:53.49" />
                    <SPLIT distance="350" swimtime="00:04:34.92" />
                    <SPLIT distance="400" swimtime="00:05:15.75" />
                    <SPLIT distance="450" swimtime="00:05:56.90" />
                    <SPLIT distance="550" swimtime="00:07:21.34" />
                    <SPLIT distance="650" swimtime="00:08:44.77" />
                    <SPLIT distance="750" swimtime="00:10:07.50" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1275" points="411" swimtime="00:02:45.51" resultid="3041" heatid="5342" lane="7" entrytime="00:02:47.67" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.33" />
                    <SPLIT distance="100" swimtime="00:01:19.74" />
                    <SPLIT distance="150" swimtime="00:02:03.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1305" points="339" swimtime="00:00:41.78" resultid="3042" heatid="5372" lane="4" />
                <RESULT eventid="2328" points="443" swimtime="00:01:12.76" resultid="6002" heatid="6418" lane="7" entrytime="00:01:12.77">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.55" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Igor" lastname="De Assis Santos" birthdate="2003-02-21" gender="M" nation="BRA" license="342496" swrid="5596885" athleteid="3072" externalid="342496" level="INTERNE/IT">
              <RESULTS>
                <RESULT eventid="1104" points="479" swimtime="00:00:26.71" resultid="3073" heatid="5128" lane="6" entrytime="00:00:27.24" entrycourse="LCM" />
                <RESULT eventid="1151" points="350" swimtime="00:02:41.73" resultid="3074" heatid="5200" lane="7" entrytime="00:02:36.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.93" />
                    <SPLIT distance="100" swimtime="00:01:10.43" />
                    <SPLIT distance="150" swimtime="00:02:02.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="439" swimtime="00:01:07.89" resultid="3075" heatid="5263" lane="1" entrytime="00:01:05.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="433" swimtime="00:00:31.12" resultid="3076" heatid="5287" lane="1" entrytime="00:00:31.00" entrycourse="LCM" />
                <RESULT eventid="1267" points="453" swimtime="00:00:28.98" resultid="3077" heatid="5330" lane="5" />
                <RESULT eventid="1297" points="367" swimtime="00:00:36.22" resultid="3078" heatid="5365" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Marques Petry" birthdate="2008-01-08" gender="M" nation="BRA" license="392352" swrid="4795316" athleteid="3113" externalid="392352" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1088" points="288" swimtime="00:01:26.10" resultid="3114" heatid="5083" lane="3" entrytime="00:01:29.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1120" points="391" swimtime="00:02:19.40" resultid="3115" heatid="5154" lane="1" entrytime="00:02:19.88" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.05" />
                    <SPLIT distance="150" swimtime="00:01:43.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="360" swimtime="00:02:40.20" resultid="3116" heatid="5196" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.27" />
                    <SPLIT distance="100" swimtime="00:01:17.70" />
                    <SPLIT distance="150" swimtime="00:02:04.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="425" swimtime="00:01:02.30" resultid="3117" heatid="5226" lane="6" entrytime="00:01:02.24" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1217" points="334" swimtime="00:10:51.38" resultid="3118" heatid="5297" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.04" />
                    <SPLIT distance="100" swimtime="00:01:13.46" />
                    <SPLIT distance="150" swimtime="00:01:54.69" />
                    <SPLIT distance="200" swimtime="00:02:36.67" />
                    <SPLIT distance="250" swimtime="00:03:18.85" />
                    <SPLIT distance="300" swimtime="00:04:01.49" />
                    <SPLIT distance="350" swimtime="00:04:43.39" />
                    <SPLIT distance="400" swimtime="00:05:25.40" />
                    <SPLIT distance="450" swimtime="00:06:06.36" />
                    <SPLIT distance="500" swimtime="00:06:47.95" />
                    <SPLIT distance="550" swimtime="00:07:29.54" />
                    <SPLIT distance="600" swimtime="00:08:11.52" />
                    <SPLIT distance="650" swimtime="00:08:52.23" />
                    <SPLIT distance="700" swimtime="00:09:33.39" />
                    <SPLIT distance="750" swimtime="00:10:12.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1251" points="279" swimtime="00:03:11.99" resultid="3119" heatid="5316" lane="5" entrytime="00:03:16.51" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.06" />
                    <SPLIT distance="100" swimtime="00:01:34.61" />
                    <SPLIT distance="150" swimtime="00:02:25.63" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Resende Ames" birthdate="2010-02-02" gender="M" nation="BRA" license="365505" swrid="5588876" athleteid="3148" externalid="365505" level="ITAIPU BIN">
              <RESULTS>
                <RESULT eventid="1104" points="461" swimtime="00:00:27.05" resultid="3149" heatid="5119" lane="8" entrytime="00:00:28.66" entrycourse="LCM" />
                <RESULT eventid="1135" points="407" swimtime="00:01:06.71" resultid="3150" heatid="5171" lane="3" entrytime="00:01:08.21" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="469" swimtime="00:01:06.38" resultid="3151" heatid="5258" lane="5" entrytime="00:01:06.69" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.84" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1213" points="425" swimtime="00:00:31.30" resultid="3152" heatid="5286" lane="3" entrytime="00:00:31.79" entrycourse="LCM" />
                <RESULT eventid="1277" points="428" swimtime="00:02:28.48" resultid="3153" heatid="5347" lane="3" entrytime="00:02:25.32" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.45" />
                    <SPLIT distance="100" swimtime="00:01:10.59" />
                    <SPLIT distance="150" swimtime="00:01:49.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="217" swimtime="00:00:43.18" resultid="3154" heatid="5363" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
          <RELAYS>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="M" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1237" points="491" swimtime="00:03:58.53" resultid="3169" heatid="5308" lane="3" entrytime="00:04:04.70">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.93" />
                    <SPLIT distance="100" swimtime="00:00:56.53" />
                    <SPLIT distance="150" swimtime="00:01:23.53" />
                    <SPLIT distance="200" swimtime="00:01:53.58" />
                    <SPLIT distance="250" swimtime="00:02:23.84" />
                    <SPLIT distance="300" swimtime="00:02:56.00" />
                    <SPLIT distance="350" swimtime="00:03:26.03" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3051" number="1" />
                    <RELAYPOSITION athleteid="3086" number="2" />
                    <RELAYPOSITION athleteid="3113" number="3" />
                    <RELAYPOSITION athleteid="3106" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1338" points="348" swimtime="00:04:53.74" resultid="3174" heatid="5388" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.66" />
                    <SPLIT distance="100" swimtime="00:01:15.28" />
                    <SPLIT distance="150" swimtime="00:01:55.99" />
                    <SPLIT distance="200" swimtime="00:02:39.56" />
                    <SPLIT distance="250" swimtime="00:03:11.57" />
                    <SPLIT distance="300" swimtime="00:03:49.16" />
                    <SPLIT distance="350" swimtime="00:04:19.44" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3051" number="1" />
                    <RELAYPOSITION athleteid="3113" number="2" />
                    <RELAYPOSITION athleteid="3086" number="3" />
                    <RELAYPOSITION athleteid="3106" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="-1" agemin="20" agetotalmax="-1" agetotalmin="-1" gender="M" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1241" points="539" swimtime="00:03:51.29" resultid="3170" heatid="5310" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.26" />
                    <SPLIT distance="100" swimtime="00:00:56.80" />
                    <SPLIT distance="150" swimtime="00:01:23.50" />
                    <SPLIT distance="200" swimtime="00:01:53.63" />
                    <SPLIT distance="250" swimtime="00:02:20.15" />
                    <SPLIT distance="300" swimtime="00:02:51.12" />
                    <SPLIT distance="350" swimtime="00:03:18.50" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3065" number="1" />
                    <RELAYPOSITION athleteid="3079" number="2" />
                    <RELAYPOSITION athleteid="3058" number="3" />
                    <RELAYPOSITION athleteid="3072" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1342" points="466" swimtime="00:04:26.68" resultid="3172" heatid="5390" lane="7">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.05" />
                    <SPLIT distance="100" swimtime="00:01:04.07" />
                    <SPLIT distance="150" swimtime="00:01:43.21" />
                    <SPLIT distance="200" swimtime="00:02:28.80" />
                    <SPLIT distance="250" swimtime="00:02:57.06" />
                    <SPLIT distance="300" swimtime="00:03:29.87" />
                    <SPLIT distance="350" swimtime="00:03:57.00" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3058" number="1" />
                    <RELAYPOSITION athleteid="3072" number="2" />
                    <RELAYPOSITION athleteid="3065" number="3" />
                    <RELAYPOSITION athleteid="3079" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="M" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1233" points="377" swimtime="00:04:20.55" resultid="3171" heatid="5306" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.90" />
                    <SPLIT distance="100" swimtime="00:00:58.65" />
                    <SPLIT distance="150" swimtime="00:01:29.29" />
                    <SPLIT distance="200" swimtime="00:02:02.25" />
                    <SPLIT distance="250" swimtime="00:02:30.58" />
                    <SPLIT distance="300" swimtime="00:03:01.42" />
                    <SPLIT distance="350" swimtime="00:03:38.04" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3148" number="1" />
                    <RELAYPOSITION athleteid="3141" number="2" />
                    <RELAYPOSITION athleteid="3162" number="3" />
                    <RELAYPOSITION athleteid="3127" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
                <RESULT eventid="1334" points="321" swimtime="00:05:01.69" resultid="3173" heatid="5386" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.64" />
                    <SPLIT distance="150" swimtime="00:01:47.36" />
                    <SPLIT distance="250" swimtime="00:03:06.10" />
                    <SPLIT distance="300" swimtime="00:03:42.01" />
                    <SPLIT distance="350" swimtime="00:04:18.40" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3148" number="1" />
                    <RELAYPOSITION athleteid="3162" number="2" />
                    <RELAYPOSITION athleteid="3141" number="3" />
                    <RELAYPOSITION athleteid="3127" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="16" agemin="16" agetotalmax="-1" agetotalmin="-1" gender="X" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1287" points="426" swimtime="00:04:49.09" resultid="3175" heatid="5354" lane="3" entrytime="00:04:42.42">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.90" />
                    <SPLIT distance="100" swimtime="00:01:21.40" />
                    <SPLIT distance="150" swimtime="00:01:56.22" />
                    <SPLIT distance="200" swimtime="00:02:37.03" />
                    <SPLIT distance="250" swimtime="00:03:12.02" />
                    <SPLIT distance="300" swimtime="00:03:52.74" />
                    <SPLIT distance="350" swimtime="00:04:18.83" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3099" number="1" />
                    <RELAYPOSITION athleteid="3086" number="2" />
                    <RELAYPOSITION athleteid="3036" number="3" />
                    <RELAYPOSITION athleteid="3051" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
            <RELAY agemax="14" agemin="14" agetotalmax="-1" agetotalmin="-1" gender="X" name="CATARATAS &quot;A&quot;" number="1">
              <RESULTS>
                <RESULT eventid="1283" points="392" swimtime="00:04:57.10" resultid="3176" heatid="5352" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.66" />
                    <SPLIT distance="150" swimtime="00:01:52.61" />
                    <SPLIT distance="200" swimtime="00:02:42.56" />
                    <SPLIT distance="250" swimtime="00:03:12.45" />
                    <SPLIT distance="300" swimtime="00:03:48.52" />
                    <SPLIT distance="350" swimtime="00:04:21.42" />
                  </SPLITS>
                  <RELAYPOSITIONS>
                    <RELAYPOSITION athleteid="3162" number="1" />
                    <RELAYPOSITION athleteid="3155" number="2" />
                    <RELAYPOSITION athleteid="3148" number="3" />
                    <RELAYPOSITION athleteid="3134" number="4" />
                  </RELAYPOSITIONS>
                </RESULT>
              </RESULTS>
            </RELAY>
          </RELAYS>
        </CLUB>
        <CLUB type="NATION" code="15969" nation="USA" clubid="4088" name="United States of America" shortname="USA">
          <ATHLETES>
            <ATHLETE firstname="Sophia" lastname="Alanis Whitney" birthdate="2007-07-21" gender="F" nation="USA" license="V397028" athleteid="4089" externalid="V397028">
              <RESULTS>
                <RESULT eventid="1096" points="458" status="EXH" swimtime="00:00:30.62" resultid="4090" heatid="5105" lane="5" />
                <RESULT eventid="1128" points="507" status="EXH" swimtime="00:01:09.54" resultid="4091" heatid="5162" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1175" points="414" status="EXH" swimtime="00:01:16.89" resultid="4092" heatid="5248" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1159" points="452" status="EXH" swimtime="00:01:07.33" resultid="4093" heatid="5209" lane="8">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1215" points="425" status="EXH" swimtime="00:00:35.70" resultid="4094" heatid="5290" lane="5" />
                <RESULT eventid="1259" points="482" status="EXH" swimtime="00:00:31.15" resultid="4095" heatid="5322" lane="3" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16044" nation="BRA" region="SC" clubid="4216" swrid="94001" name="Instituto Core">
          <ATHLETES>
            <ATHLETE firstname="Valentino" lastname="Thoth Da Silva" birthdate="2009-08-22" gender="M" nation="BRA" license="378150" swrid="5756256" athleteid="4217" externalid="378150">
              <RESULTS>
                <RESULT eventid="1104" points="496" status="EXH" swimtime="00:00:26.41" resultid="4218" heatid="5125" lane="5" entrytime="00:00:26.06" entrycourse="LCM" />
                <RESULT eventid="1135" points="463" status="EXH" swimtime="00:01:03.92" resultid="4219" heatid="5174" lane="5" entrytime="00:01:02.22" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="489" status="EXH" swimtime="00:00:59.45" resultid="4220" heatid="5228" lane="7" entrytime="00:00:58.93" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="515" status="EXH" swimtime="00:00:27.77" resultid="4221" heatid="5335" lane="5" entrytime="00:00:28.12" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vinícius" lastname="Da Rosa Maia" birthdate="2008-02-12" gender="M" nation="BRA" license="378158" swrid="5756200" athleteid="4222" externalid="378158">
              <RESULTS>
                <RESULT eventid="1104" points="519" status="EXH" swimtime="00:00:26.01" resultid="4223" heatid="5121" lane="2" />
                <RESULT eventid="1135" points="437" status="EXH" swimtime="00:01:05.14" resultid="4224" heatid="5172" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.10" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" points="420" status="EXH" swimtime="00:01:08.86" resultid="4225" heatid="5259" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.90" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Mendes Costa" birthdate="2010-05-27" gender="F" nation="BRA" license="392182" swrid="5756233" athleteid="4226" externalid="392182">
              <RESULTS>
                <RESULT comment="SW 4.4 - Antecipou-se ao sinal de partida.  (Horário: 10:58)" eventid="1275" status="DSQ" swimtime="00:02:48.41" resultid="4227" heatid="5341" lane="5" entrytime="00:02:49.63" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.45" />
                    <SPLIT distance="100" swimtime="00:01:23.94" />
                    <SPLIT distance="150" swimtime="00:02:09.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16131" nation="BRA" region="PR" clubid="4050" swrid="93766" name="Associação Nadar Colombo" shortname="Equipe Nadar">
          <ATHLETES>
            <ATHLETE firstname="Gabriel" lastname="Guarise" birthdate="2008-11-28" gender="M" nation="BRA" license="408881" swrid="5727650" athleteid="4080" externalid="408881">
              <RESULTS>
                <RESULT eventid="1104" points="405" swimtime="00:00:28.24" resultid="4081" heatid="5122" lane="6" entrytime="00:00:28.70" entrycourse="LCM" />
                <RESULT eventid="1167" points="389" swimtime="00:01:04.15" resultid="4082" heatid="5225" lane="1" entrytime="00:01:08.26" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1297" points="338" swimtime="00:00:37.22" resultid="4083" heatid="5368" lane="8" entrytime="00:00:37.99" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Fernanda" lastname="Krik" birthdate="2010-11-24" gender="F" nation="BRA" license="406702" swrid="5717277" athleteid="4077" externalid="406702">
              <RESULTS>
                <RESULT eventid="1080" points="136" swimtime="00:02:04.70" resultid="4078" heatid="5065" lane="7" entrytime="00:02:05.08" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1064" points="179" swimtime="00:06:56.98" resultid="4079" heatid="5048" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.29" />
                    <SPLIT distance="100" swimtime="00:01:36.58" />
                    <SPLIT distance="150" swimtime="00:02:30.98" />
                    <SPLIT distance="200" swimtime="00:03:23.96" />
                    <SPLIT distance="250" swimtime="00:04:16.99" />
                    <SPLIT distance="300" swimtime="00:05:10.94" />
                    <SPLIT distance="350" swimtime="00:06:05.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Carvalho Ezaki" birthdate="2011-10-20" gender="F" nation="BRA" license="399927" swrid="5652882" athleteid="4069" externalid="399927">
              <RESULTS>
                <RESULT eventid="1080" points="282" swimtime="00:01:37.75" resultid="4070" heatid="5065" lane="5" entrytime="00:01:37.59" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="272" swimtime="00:03:14.51" resultid="4071" heatid="5186" lane="5" entrytime="00:03:17.97" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.04" />
                    <SPLIT distance="100" swimtime="00:01:40.55" />
                    <SPLIT distance="150" swimtime="00:02:33.22" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1259" points="196" swimtime="00:00:42.01" resultid="4072" heatid="5323" lane="6" entrytime="00:00:41.70" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="João" lastname="Marcelo Santos Poli" birthdate="2007-09-01" gender="M" nation="BRA" license="388175" swrid="5622292" athleteid="4062" externalid="388175">
              <RESULTS>
                <RESULT eventid="1151" points="262" swimtime="00:02:58.10" resultid="4063" heatid="5199" lane="5" entrytime="00:03:04.42" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.70" />
                    <SPLIT distance="100" swimtime="00:01:23.32" />
                    <SPLIT distance="150" swimtime="00:02:21.32" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1182" status="DNS" swimtime="00:00:00.00" resultid="4064" heatid="5262" lane="2" entrytime="00:01:13.65" entrycourse="LCM" />
                <RESULT eventid="1277" points="282" swimtime="00:02:50.67" resultid="4065" heatid="5345" lane="6" entrytime="00:02:46.73" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.11" />
                    <SPLIT distance="100" swimtime="00:01:23.20" />
                    <SPLIT distance="150" swimtime="00:02:08.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Rafael D Agostin Batistao" birthdate="2008-05-13" gender="M" nation="BRA" license="384738" swrid="5622300" athleteid="4051" externalid="384738">
              <RESULTS>
                <RESULT eventid="1088" status="SICK" swimtime="00:00:00.00" resultid="4052" heatid="5083" lane="4" entrytime="00:01:22.05" entrycourse="LCM" />
                <RESULT eventid="1151" status="SICK" swimtime="00:00:00.00" resultid="4053" heatid="5197" lane="8" entrytime="00:02:56.60" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Santos Poli" birthdate="2010-02-19" gender="M" nation="BRA" license="414563" swrid="5755378" athleteid="4084" externalid="414563">
              <RESULTS>
                <RESULT eventid="1135" points="226" swimtime="00:01:21.07" resultid="4085" heatid="5170" lane="8" entrytime="00:01:26.16" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.62" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="217" swimtime="00:03:09.52" resultid="4086" heatid="5192" lane="5">
                  <SPLITS>
                    <SPLIT distance="100" swimtime="00:01:32.68" />
                    <SPLIT distance="150" swimtime="00:02:28.17" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="303" swimtime="00:00:33.13" resultid="4087" heatid="5331" lane="4" entrytime="00:00:35.17" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Glir" birthdate="2010-07-01" gender="M" nation="BRA" license="406701" swrid="5717266" athleteid="4073" externalid="406701">
              <RESULTS>
                <RESULT eventid="1088" points="231" swimtime="00:01:32.65" resultid="4074" heatid="5079" lane="4" entrytime="00:01:32.80" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1151" points="264" swimtime="00:02:57.57" resultid="4075" heatid="5192" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.00" />
                    <SPLIT distance="150" swimtime="00:02:20.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="334" swimtime="00:01:07.51" resultid="4076" heatid="5219" lane="3" entrytime="00:01:10.12" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Rosa De Souza" birthdate="2009-01-01" gender="F" nation="BRA" license="399926" swrid="5653301" athleteid="4066" externalid="399926">
              <RESULTS>
                <RESULT eventid="1064" points="210" swimtime="00:06:35.78" resultid="4067" heatid="5052" lane="5" entrytime="00:06:27.23" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.47" />
                    <SPLIT distance="100" swimtime="00:01:32.85" />
                    <SPLIT distance="150" swimtime="00:02:23.20" />
                    <SPLIT distance="200" swimtime="00:03:15.71" />
                    <SPLIT distance="250" swimtime="00:04:08.14" />
                    <SPLIT distance="300" swimtime="00:05:01.22" />
                    <SPLIT distance="350" swimtime="00:05:49.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="215" swimtime="00:03:30.39" resultid="4068" heatid="5189" lane="7" entrytime="00:03:25.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.46" />
                    <SPLIT distance="100" swimtime="00:01:39.52" />
                    <SPLIT distance="150" swimtime="00:02:44.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kaylaine" lastname="Sofia Vargas Bueno" birthdate="2006-11-28" gender="F" nation="BRA" license="384739" swrid="5622307" athleteid="4054" externalid="384739">
              <RESULTS>
                <RESULT eventid="1064" points="260" swimtime="00:06:08.70" resultid="4055" heatid="5054" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.82" />
                    <SPLIT distance="100" swimtime="00:01:28.00" />
                    <SPLIT distance="150" swimtime="00:02:15.61" />
                    <SPLIT distance="200" swimtime="00:03:03.73" />
                    <SPLIT distance="250" swimtime="00:03:51.55" />
                    <SPLIT distance="300" swimtime="00:04:38.61" />
                    <SPLIT distance="350" swimtime="00:05:25.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1112" points="301" swimtime="00:02:48.21" resultid="4056" heatid="5145" lane="4" entrytime="00:02:57.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.68" />
                    <SPLIT distance="100" swimtime="00:01:21.44" />
                    <SPLIT distance="150" swimtime="00:02:05.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1143" points="240" swimtime="00:03:22.85" resultid="4057" heatid="5191" lane="7" entrytime="00:03:20.89" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.86" />
                    <SPLIT distance="100" swimtime="00:01:41.81" />
                    <SPLIT distance="150" swimtime="00:02:41.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Luiz Sartori" birthdate="2008-04-07" gender="M" nation="BRA" license="384742" swrid="5622287" athleteid="4058" externalid="384742">
              <RESULTS>
                <RESULT eventid="1120" points="426" swimtime="00:02:15.49" resultid="4059" heatid="5154" lane="4" entrytime="00:02:17.14" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.62" />
                    <SPLIT distance="100" swimtime="00:01:05.83" />
                    <SPLIT distance="150" swimtime="00:01:41.28" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1167" points="483" swimtime="00:00:59.70" resultid="4060" heatid="5227" lane="4" entrytime="00:00:59.28" entrycourse="LCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1267" points="448" swimtime="00:00:29.10" resultid="4061" heatid="5334" lane="6" entrytime="00:00:29.43" entrycourse="LCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
