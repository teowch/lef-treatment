<?xml version="1.0" encoding="UTF-8"?>
<LENEX version="3.0">
  <CONSTRUCTOR name="SPLASH Meet Manager 11" registration="Swim Time Brasil" version="11.79293">
    <CONTACT name="Splash Software GmbH" street="Ahornweg 41" city="Spiegel b. Bern" zip="3095" country="CH" email="sales@swimrankings.net" internet="https://www.swimrankings.net" />
  </CONSTRUCTOR>
  <MEETS>
    <MEET city="Maringá" name="Torneio Regional da 2ª Região (Pré-Mirim/Sênior)" course="SCM" deadline="2024-04-01" entrystartdate="2024-03-26" entrytype="INVITATION" hostclub="Universidade Estadual de Maringá" hostclub.url="http://www.uem.br/" number="38303" organizer="Federação de Desportos Aquáticos do Paraná" organizer.url="https://www.fdap.org.br/" reservecount="2" result.url="https://www.swimtimebrasil.com/evento/natacao/38303" startmethod="1" timing="AUTOMATIC" masters="F" withdrawuntil="2024-04-02" state="PR" nation="BRA">
      <AGEDATE value="2024-04-06" type="YEAR" />
      <POOL name="Universidade Estadual de Maringá" lanemin="1" lanemax="6" />
      <FACILITY city="Maringá" name="Universidade Estadual de Maringá" nation="BRA" state="PR" street="M19" street2="Vila Esperança" zip="87020-900" />
      <POINTTABLE pointtableid="3016" name="FINA Point Scoring" version="2023" />
      <QUALIFY from="2023-04-06" until="2024-04-05" />
      <CONTACT city="Curitiba" email="ti@fdap.org.br" fax="+55 (41) 99206-4448" name="Federação de Desportos Aquáticos do Paraná" phone="+55 (41) 99206-4448" street="Avenida do Batel, 1230" street2="Batel" zip="80420-090" />
      <SESSIONS>
        <SESSION date="2024-04-06" daytime="09:10" endtime="11:52" number="1" officialmeeting="08:30" teamleadermeeting="09:00" warmupfrom="08:00" warmupuntil="09:00">
          <EVENTS>
            <EVENT eventid="1060" daytime="09:10" gender="F" number="1" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1061" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1544" />
                    <RANKING order="2" place="2" resultid="1690" />
                    <RANKING order="3" place="3" resultid="1419" />
                    <RANKING order="4" place="4" resultid="1437" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1062" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1673" />
                    <RANKING order="2" place="2" resultid="1760" />
                    <RANKING order="3" place="3" resultid="1487" />
                    <RANKING order="4" place="4" resultid="1429" />
                    <RANKING order="5" place="5" resultid="1475" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1791" daytime="09:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1792" daytime="09:16" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1063" daytime="09:22" gender="M" number="2" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1064" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1756" />
                    <RANKING order="2" place="2" resultid="1516" />
                    <RANKING order="3" place="3" resultid="1552" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1065" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1669" />
                    <RANKING order="2" place="2" resultid="1706" />
                    <RANKING order="3" place="3" resultid="1661" />
                    <RANKING order="4" place="4" resultid="1415" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1793" daytime="09:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1794" daytime="09:26" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1066" daytime="09:32" gender="F" number="3" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1067" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1492" />
                    <RANKING order="2" place="2" resultid="1410" />
                    <RANKING order="3" place="3" resultid="1421" />
                    <RANKING order="4" place="4" resultid="1732" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1068" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1326" />
                    <RANKING order="2" place="2" resultid="1323" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1069" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1070" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1378" />
                    <RANKING order="2" place="2" resultid="1396" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1071" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1336" />
                    <RANKING order="2" place="2" resultid="1618" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1072" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1368" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1073" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1795" daytime="09:32" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1796" daytime="09:34" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1074" daytime="09:36" gender="M" number="4" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1075" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1404" />
                    <RANKING order="2" place="2" resultid="1717" />
                    <RANKING order="3" place="3" resultid="1676" />
                    <RANKING order="4" place="4" resultid="1623" />
                    <RANKING order="5" place="5" resultid="1693" />
                    <RANKING order="6" place="6" resultid="1333" />
                    <RANKING order="7" place="7" resultid="1489" />
                    <RANKING order="8" place="8" resultid="1770" />
                    <RANKING order="9" place="-1" resultid="1726" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1076" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1527" />
                    <RANKING order="2" place="-1" resultid="1655" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1077" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1393" />
                    <RANKING order="2" place="2" resultid="1424" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1078" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1352" />
                    <RANKING order="2" place="2" resultid="1329" />
                    <RANKING order="3" place="3" resultid="1647" />
                    <RANKING order="4" place="4" resultid="1316" />
                    <RANKING order="5" place="5" resultid="1495" />
                    <RANKING order="6" place="6" resultid="1614" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1079" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1611" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1080" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1340" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1081" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1633" />
                    <RANKING order="2" place="2" resultid="1582" />
                    <RANKING order="3" place="3" resultid="1522" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1797" daytime="09:36" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1798" daytime="09:40" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1799" daytime="09:42" number="3" order="3" status="OFFICIAL" />
                <HEAT heatid="1800" daytime="09:44" number="4" order="4" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1082" daytime="09:48" gender="F" number="5" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1083" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1708" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1084" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1681" />
                    <RANKING order="2" place="2" resultid="1457" />
                    <RANKING order="3" place="3" resultid="1432" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1801" daytime="09:48" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1085" daytime="09:56" gender="M" number="6" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1086" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1444" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1087" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1448" />
                    <RANKING order="2" place="2" resultid="1452" />
                    <RANKING order="3" place="3" resultid="1750" />
                    <RANKING order="4" place="-1" resultid="1440" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1802" daytime="09:56" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1088" daytime="10:04" gender="F" number="7" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1089" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1524" />
                    <RANKING order="2" place="2" resultid="1730" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1090" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1636" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1091" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1092" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1093" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1094" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1095" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1803" daytime="10:04" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1096" daytime="10:10" gender="M" number="8" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1097" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1407" />
                    <RANKING order="2" place="2" resultid="1361" />
                    <RANKING order="3" place="-1" resultid="1332" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1098" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1654" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1099" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1100" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1390" />
                    <RANKING order="2" place="2" resultid="1358" />
                    <RANKING order="3" place="3" resultid="1642" />
                    <RANKING order="4" place="4" resultid="1503" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1101" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1311" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1102" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1103" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1343" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1804" daytime="10:10" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1805" daytime="10:14" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1104" daytime="10:18" gender="F" number="9" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1105" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1543" />
                    <RANKING order="2" place="2" resultid="1689" />
                    <RANKING order="3" place="3" resultid="1709" />
                    <RANKING order="4" place="4" resultid="1417" />
                    <RANKING order="5" place="5" resultid="1460" />
                    <RANKING order="6" place="6" resultid="1651" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1106" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1665" />
                    <RANKING order="2" place="2" resultid="1671" />
                    <RANKING order="3" place="3" resultid="1433" />
                    <RANKING order="4" place="4" resultid="1758" />
                    <RANKING order="5" place="5" resultid="1473" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1806" daytime="10:18" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1807" daytime="10:20" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1107" daytime="10:22" gender="M" number="10" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1108" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1519" />
                    <RANKING order="2" place="2" resultid="1754" />
                    <RANKING order="3" place="3" resultid="1511" />
                    <RANKING order="4" place="4" resultid="1514" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1109" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1449" />
                    <RANKING order="2" place="2" resultid="1668" />
                    <RANKING order="3" place="3" resultid="1507" />
                    <RANKING order="4" place="4" resultid="1559" />
                    <RANKING order="5" place="-1" resultid="1751" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1808" daytime="10:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1809" daytime="10:24" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1110" daytime="10:28" gender="F" number="11" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1111" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1112" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1637" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1113" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1114" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1115" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1319" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1116" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1117" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1810" daytime="10:28" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1118" daytime="10:38" gender="M" number="12" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="800" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1119" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1120" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1121" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1355" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1122" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1123" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1124" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1125" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1632" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1811" daytime="10:38" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1126" daytime="11:04" gender="F" number="13" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1127" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1688" />
                    <RANKING order="2" place="2" resultid="1685" />
                    <RANKING order="3" place="3" resultid="1628" />
                    <RANKING order="4" place="4" resultid="1435" />
                    <RANKING order="5" place="5" resultid="1722" />
                    <RANKING order="6" place="6" resultid="1650" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1128" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1664" />
                    <RANKING order="2" place="2" resultid="1456" />
                    <RANKING order="3" place="3" resultid="1485" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1812" daytime="11:04" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1813" daytime="11:08" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1129" daytime="11:12" gender="M" number="14" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1130" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1443" />
                    <RANKING order="2" place="2" resultid="1518" />
                    <RANKING order="3" place="-1" resultid="1701" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1131" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1447" />
                    <RANKING order="2" place="2" resultid="1667" />
                    <RANKING order="3" place="3" resultid="1659" />
                    <RANKING order="4" place="4" resultid="1451" />
                    <RANKING order="5" place="5" resultid="1506" />
                    <RANKING order="6" place="-1" resultid="1439" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1814" daytime="11:12" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1815" daytime="11:14" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1132" daytime="11:18" gender="F" number="15" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1133" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1134" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1467" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1135" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1381" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1136" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1137" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1617" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1138" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1367" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1139" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1816" daytime="11:18" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1140" daytime="11:22" gender="M" number="16" order="17" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1141" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1716" />
                    <RANKING order="2" place="2" resultid="1675" />
                    <RANKING order="3" place="3" resultid="1622" />
                    <RANKING order="4" place="-1" resultid="1725" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1142" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1399" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1143" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1144" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="-1" resultid="1641" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1145" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1146" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1147" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1631" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1817" daytime="11:22" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1818" daytime="11:26" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1148" daytime="11:30" gender="F" number="17" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1149" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1542" />
                    <RANKING order="2" place="2" resultid="1743" />
                    <RANKING order="3" place="3" resultid="1721" />
                    <RANKING order="4" place="4" resultid="1684" />
                    <RANKING order="5" place="5" resultid="1627" />
                    <RANKING order="6" place="6" resultid="1459" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1150" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1663" />
                    <RANKING order="2" place="2" resultid="1455" />
                    <RANKING order="3" place="3" resultid="1431" />
                    <RANKING order="4" place="4" resultid="1680" />
                    <RANKING order="5" place="5" resultid="1427" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1819" daytime="11:30" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1820" daytime="11:32" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1151" daytime="11:36" gender="M" number="18" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1152" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1510" />
                    <RANKING order="2" place="2" resultid="1550" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1153" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1704" />
                    <RANKING order="2" place="2" resultid="1413" />
                    <RANKING order="3" place="3" resultid="1558" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1821" daytime="11:36" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1154" daytime="11:38" gender="F" number="19" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1155" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1731" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1156" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1470" />
                    <RANKING order="2" place="2" resultid="1325" />
                    <RANKING order="3" place="3" resultid="1322" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1157" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1384" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1158" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1387" />
                    <RANKING order="2" place="2" resultid="1372" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1159" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1335" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1160" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1161" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1822" daytime="11:38" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1823" daytime="11:42" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1162" daytime="11:44" gender="M" number="20" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1163" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1403" />
                    <RANKING order="2" place="2" resultid="1692" />
                    <RANKING order="3" place="3" resultid="1769" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1164" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1349" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1165" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1346" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1166" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1646" />
                    <RANKING order="2" place="2" resultid="1328" />
                    <RANKING order="3" place="3" resultid="1315" />
                    <RANKING order="4" place="4" resultid="1502" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1167" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1168" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1375" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1169" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1364" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1824" daytime="11:44" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1825" daytime="11:46" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1170" daytime="11:50" gender="F" number="21" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1171" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1686" />
                    <RANKING order="2" place="2" resultid="1710" />
                    <RANKING order="3" place="3" resultid="1744" />
                    <RANKING order="4" place="4" resultid="1418" />
                    <RANKING order="5" place="5" resultid="1629" />
                    <RANKING order="6" place="6" resultid="1461" />
                    <RANKING order="7" place="7" resultid="1723" />
                    <RANKING order="8" place="8" resultid="1436" />
                    <RANKING order="9" place="9" resultid="1652" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1172" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1672" />
                    <RANKING order="2" place="2" resultid="1682" />
                    <RANKING order="3" place="3" resultid="1759" />
                    <RANKING order="4" place="4" resultid="1474" />
                    <RANKING order="5" place="5" resultid="1486" />
                    <RANKING order="6" place="6" resultid="1428" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1826" daytime="11:50" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1827" daytime="11:52" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1828" daytime="11:56" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1173" daytime="11:58" gender="M" number="22" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1174" agemax="11" agemin="11">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1445" />
                    <RANKING order="2" place="2" resultid="1755" />
                    <RANKING order="3" place="3" resultid="1512" />
                    <RANKING order="4" place="4" resultid="1520" />
                    <RANKING order="5" place="5" resultid="1515" />
                    <RANKING order="6" place="6" resultid="1551" />
                    <RANKING order="7" place="-1" resultid="1702" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1175" agemax="12" agemin="12">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1660" />
                    <RANKING order="2" place="2" resultid="1705" />
                    <RANKING order="3" place="3" resultid="1453" />
                    <RANKING order="4" place="4" resultid="1752" />
                    <RANKING order="5" place="5" resultid="1508" />
                    <RANKING order="6" place="6" resultid="1560" />
                    <RANKING order="7" place="7" resultid="1414" />
                    <RANKING order="8" place="-1" resultid="1441" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1829" daytime="11:58" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1830" daytime="12:02" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1831" daytime="12:04" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
        <SESSION date="2024-04-06" daytime="15:40" endtime="17:44" number="2" officialmeeting="15:00" warmupfrom="14:30" warmupuntil="15:30">
          <EVENTS>
            <EVENT eventid="1176" daytime="15:40" gender="F" number="23" order="1" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1177" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1178" daytime="15:40" gender="M" number="24" order="2" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1179" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1778" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1832" daytime="15:40" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1180" daytime="15:42" gender="F" number="25" order="3" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1181" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1534" />
                    <RANKING order="2" place="2" resultid="1575" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1182" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1698" />
                    <RANKING order="2" place="2" resultid="1580" />
                    <RANKING order="3" place="3" resultid="1464" />
                    <RANKING order="4" place="4" resultid="1584" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1833" daytime="15:42" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1183" daytime="15:46" gender="M" number="26" order="4" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1184" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1714" />
                    <RANKING order="2" place="2" resultid="1555" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1185" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1478" />
                    <RANKING order="2" place="2" resultid="1548" />
                    <RANKING order="3" place="3" resultid="1747" />
                    <RANKING order="4" place="4" resultid="1482" />
                    <RANKING order="5" place="5" resultid="1568" />
                    <RANKING order="6" place="6" resultid="1530" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1834" daytime="15:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1835" daytime="15:48" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1186" daytime="15:52" gender="F" number="27" order="5" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1187" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1188" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1189" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1190" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1191" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1192" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1193" agemax="-1" agemin="20" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1194" daytime="15:52" gender="M" number="28" order="6" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="400" relaycount="1" stroke="MEDLEY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1195" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1196" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1197" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1356" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1198" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1199" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1200" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1376" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1201" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1836" daytime="15:52" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1202" daytime="16:00" gender="F" number="29" order="7" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1203" agemax="9" agemin="9" />
                <AGEGROUP agegroupid="1204" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1572" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1837" daytime="16:00" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1205" daytime="16:04" gender="M" number="30" order="8" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1206" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1500" />
                    <RANKING order="2" place="2" resultid="1540" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1207" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1767" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1838" daytime="16:04" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1208" daytime="16:06" gender="F" number="31" order="9" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1209" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1210" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1471" />
                    <RANKING order="2" place="2" resultid="1639" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1211" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1212" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1373" />
                    <RANKING order="2" place="2" resultid="1397" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1213" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1320" />
                    <RANKING order="2" place="2" resultid="1620" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1214" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1370" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1215" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1839" daytime="16:06" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1840" daytime="16:10" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1216" daytime="16:14" gender="M" number="32" order="10" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1217" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1405" />
                    <RANKING order="2" place="2" resultid="1719" />
                    <RANKING order="3" place="3" resultid="1678" />
                    <RANKING order="4" place="4" resultid="1625" />
                    <RANKING order="5" place="5" resultid="1772" />
                    <RANKING order="6" place="-1" resultid="1728" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1218" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1528" />
                    <RANKING order="2" place="-1" resultid="1657" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1219" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1220" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1644" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1221" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1313" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1222" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1341" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1223" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1841" daytime="16:14" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1842" daytime="16:18" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1224" daytime="16:22" gender="F" number="33" order="11" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1225" agemax="8" agemin="8" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1226" daytime="16:22" gender="M" number="34" order="12" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1227" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1593" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1843" daytime="16:22" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1228" daytime="16:26" gender="F" number="35" order="13" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1229" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1535" />
                    <RANKING order="2" place="2" resultid="1576" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1230" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1585" />
                    <RANKING order="2" place="2" resultid="1740" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1844" daytime="16:26" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1231" daytime="16:28" gender="M" number="36" order="14" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1232" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1498" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1233" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1479" />
                    <RANKING order="2" place="2" resultid="1483" />
                    <RANKING order="3" place="3" resultid="1531" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1845" daytime="16:28" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1234" daytime="16:30" gender="F" number="37" order="15" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1235" agemax="13" agemin="13" />
                <AGEGROUP agegroupid="1236" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1237" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1238" agemax="16" agemin="16" />
                <AGEGROUP agegroupid="1239" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1240" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1241" agemax="-1" agemin="20" />
              </AGEGROUPS>
            </EVENT>
            <EVENT eventid="1242" daytime="16:30" gender="M" number="38" order="16" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="200" relaycount="1" stroke="FLY" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1243" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1695" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1244" agemax="14" agemin="14" />
                <AGEGROUP agegroupid="1245" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1394" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1246" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1648" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1247" agemax="17" agemin="17" />
                <AGEGROUP agegroupid="1248" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1249" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1846" daytime="16:30" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1250" daytime="16:50" gender="F" number="39" order="18" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1251" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1781" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1847" daytime="16:50" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1252" daytime="16:52" gender="M" number="40" order="19" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1253" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1594" />
                    <RANKING order="2" place="2" resultid="1786" />
                    <RANKING order="3" place="-1" resultid="1788" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1848" daytime="16:52" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1254" daytime="16:54" gender="F" number="41" order="20" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1255" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1737" />
                    <RANKING order="2" place="2" resultid="1608" />
                    <RANKING order="3" place="3" resultid="1563" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1256" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1579" />
                    <RANKING order="2" place="2" resultid="1697" />
                    <RANKING order="3" place="3" resultid="1571" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1849" daytime="16:54" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1257" daytime="16:56" gender="M" number="42" order="21" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1258" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1713" />
                    <RANKING order="2" place="2" resultid="1554" />
                    <RANKING order="3" place="3" resultid="1604" />
                    <RANKING order="4" place="4" resultid="1597" />
                    <RANKING order="5" place="-1" resultid="1589" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1259" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1547" />
                    <RANKING order="2" place="2" resultid="1481" />
                    <RANKING order="3" place="3" resultid="1567" />
                    <RANKING order="4" place="4" resultid="1600" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1850" daytime="16:56" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1851" daytime="17:00" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1260" daytime="17:02" gender="F" number="43" order="22" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1261" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1493" />
                    <RANKING order="2" place="2" resultid="1411" />
                    <RANKING order="3" place="3" resultid="1422" />
                    <RANKING order="4" place="4" resultid="1734" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1262" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1468" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1263" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1382" />
                    <RANKING order="2" place="2" resultid="1385" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1264" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1388" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1265" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1619" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1266" agemax="19" agemin="18">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1369" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1267" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1852" daytime="17:02" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1853" daytime="17:06" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1268" daytime="17:08" gender="M" number="44" order="23" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BACK" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1269" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1718" />
                    <RANKING order="2" place="2" resultid="1624" />
                    <RANKING order="3" place="3" resultid="1677" />
                    <RANKING order="4" place="4" resultid="1490" />
                    <RANKING order="5" place="-1" resultid="1727" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1270" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1401" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1271" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1272" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1353" />
                    <RANKING order="2" place="2" resultid="1317" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1273" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1612" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1274" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1275" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1365" />
                    <RANKING order="2" place="2" resultid="1634" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1854" daytime="17:08" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1855" daytime="17:12" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1276" daytime="17:16" gender="F" number="45" order="24" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1277" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1536" />
                    <RANKING order="2" place="2" resultid="1609" />
                    <RANKING order="3" place="3" resultid="1564" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1278" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1465" />
                    <RANKING order="2" place="2" resultid="1699" />
                    <RANKING order="3" place="3" resultid="1586" />
                    <RANKING order="4" place="4" resultid="1741" />
                    <RANKING order="5" place="-1" resultid="1763" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1856" daytime="17:16" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1857" daytime="17:18" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1279" daytime="17:20" gender="M" number="46" order="25" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1280" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1556" />
                    <RANKING order="2" place="2" resultid="1499" />
                    <RANKING order="3" place="3" resultid="1539" />
                    <RANKING order="4" place="4" resultid="1605" />
                    <RANKING order="5" place="-1" resultid="1590" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1281" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1748" />
                    <RANKING order="2" place="2" resultid="1775" />
                    <RANKING order="3" place="3" resultid="1532" />
                    <RANKING order="4" place="4" resultid="1766" />
                    <RANKING order="5" place="5" resultid="1601" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1858" daytime="17:20" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1859" daytime="17:22" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1282" daytime="17:24" gender="F" number="47" order="26" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1283" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1525" />
                    <RANKING order="2" place="2" resultid="1733" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1284" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1638" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1285" agemax="15" agemin="15" />
                <AGEGROUP agegroupid="1286" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1379" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1287" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1337" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1288" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1289" agemax="-1" agemin="20" />
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1860" daytime="17:24" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1290" daytime="17:28" gender="M" number="48" order="27" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="100" relaycount="1" stroke="BREAST" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1291" agemax="13" agemin="13">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1408" />
                    <RANKING order="2" place="2" resultid="1362" />
                    <RANKING order="3" place="3" resultid="1694" />
                    <RANKING order="4" place="4" resultid="1771" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1292" agemax="14" agemin="14">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1350" />
                    <RANKING order="2" place="2" resultid="1656" />
                    <RANKING order="3" place="3" resultid="1400" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1293" agemax="15" agemin="15">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1347" />
                    <RANKING order="2" place="2" resultid="1425" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1294" agemax="16" agemin="16">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1391" />
                    <RANKING order="2" place="2" resultid="1359" />
                    <RANKING order="3" place="3" resultid="1330" />
                    <RANKING order="4" place="4" resultid="1643" />
                    <RANKING order="5" place="5" resultid="1496" />
                    <RANKING order="6" place="6" resultid="1504" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1295" agemax="17" agemin="17">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1312" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1296" agemax="19" agemin="18" />
                <AGEGROUP agegroupid="1297" agemax="-1" agemin="20">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1344" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1861" daytime="17:28" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1862" daytime="17:30" number="2" order="2" status="OFFICIAL" />
                <HEAT heatid="1863" daytime="17:34" number="3" order="3" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1298" daytime="17:36" gender="F" number="49" order="28" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1299" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1783" />
                    <RANKING order="2" place="2" resultid="1780" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1864" daytime="17:36" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1300" daytime="17:38" gender="M" number="50" order="29" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1301" agemax="8" agemin="8">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1777" />
                    <RANKING order="2" place="2" resultid="1592" />
                    <RANKING order="3" place="3" resultid="1785" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1865" daytime="17:38" number="1" order="1" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1302" daytime="17:40" gender="F" number="51" order="30" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1303" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1736" />
                    <RANKING order="2" place="2" resultid="1574" />
                    <RANKING order="3" place="3" resultid="1607" />
                    <RANKING order="4" place="4" resultid="1562" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1304" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1578" />
                    <RANKING order="2" place="2" resultid="1463" />
                    <RANKING order="3" place="3" resultid="1570" />
                    <RANKING order="4" place="4" resultid="1739" />
                    <RANKING order="5" place="-1" resultid="1762" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1866" daytime="17:40" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1867" daytime="17:42" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
            <EVENT eventid="1305" daytime="17:46" gender="M" number="52" order="31" round="TIM" preveventid="-1">
              <SWIMSTYLE distance="50" relaycount="1" stroke="FREE" />
              <FEE currency="BRL" value="2600" />
              <AGEGROUPS>
                <AGEGROUP agegroupid="1306" agemax="9" agemin="9">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1712" />
                    <RANKING order="2" place="2" resultid="1538" />
                    <RANKING order="3" place="3" resultid="1603" />
                    <RANKING order="4" place="4" resultid="1596" />
                    <RANKING order="5" place="-1" resultid="1588" />
                  </RANKINGS>
                </AGEGROUP>
                <AGEGROUP agegroupid="1307" agemax="10" agemin="10">
                  <RANKINGS>
                    <RANKING order="1" place="1" resultid="1477" />
                    <RANKING order="2" place="2" resultid="1546" />
                    <RANKING order="3" place="3" resultid="1746" />
                    <RANKING order="4" place="4" resultid="1566" />
                    <RANKING order="5" place="5" resultid="1765" />
                    <RANKING order="6" place="6" resultid="1774" />
                    <RANKING order="7" place="7" resultid="1599" />
                  </RANKINGS>
                </AGEGROUP>
              </AGEGROUPS>
              <HEATS>
                <HEAT heatid="1868" daytime="17:46" number="1" order="1" status="OFFICIAL" />
                <HEAT heatid="1869" daytime="17:48" number="2" order="2" status="OFFICIAL" />
              </HEATS>
            </EVENT>
          </EVENTS>
        </SESSION>
      </SESSIONS>
      <CLUBS>
        <CLUB type="CLUB" code="15981" nation="BRA" region="PR" clubid="1309" swrid="93783" name="Quinto Nado" shortname="5º Nado">
          <ATHLETES>
            <ATHLETE firstname="Maria" lastname="Fernanda Romero" birthdate="2007-04-18" gender="F" nation="BRA" license="404750" athleteid="1334" externalid="404750">
              <RESULTS>
                <RESULT eventid="1154" points="455" swimtime="00:01:10.26" resultid="1335" heatid="1822" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.88" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="513" swimtime="00:01:02.75" resultid="1336" heatid="1795" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="481" swimtime="00:01:19.55" resultid="1337" heatid="1860" lane="4" entrytime="00:01:21.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.10" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Takemura Couto" birthdate="2010-02-08" gender="F" nation="BRA" license="376950" swrid="5603919" athleteid="1324" externalid="376950">
              <RESULTS>
                <RESULT eventid="1154" points="325" swimtime="00:01:18.58" resultid="1325" heatid="1823" lane="5" entrytime="00:01:19.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="458" swimtime="00:01:05.18" resultid="1326" heatid="1796" lane="4" entrytime="00:01:05.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Guilherme" lastname="Kikuchi Fujii" birthdate="2007-01-04" gender="M" nation="BRA" license="297805" swrid="5603863" athleteid="1310" externalid="297805" level="G-OLIMPICA">
              <RESULTS>
                <RESULT eventid="1096" points="578" swimtime="00:02:24.24" resultid="1311" heatid="1805" lane="4" entrytime="00:02:23.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.18" />
                    <SPLIT distance="100" swimtime="00:01:10.19" />
                    <SPLIT distance="150" swimtime="00:01:47.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="606" swimtime="00:01:05.29" resultid="1312" heatid="1863" lane="4" entrytime="00:01:05.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="543" swimtime="00:02:01.80" resultid="1313" heatid="1841" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.32" />
                    <SPLIT distance="100" swimtime="00:00:59.32" />
                    <SPLIT distance="150" swimtime="00:01:30.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Sorace Spironelli" birthdate="2008-05-14" gender="M" nation="BRA" license="371318" swrid="5622308" athleteid="1327" externalid="371318">
              <RESULTS>
                <RESULT eventid="1162" points="357" swimtime="00:01:07.30" resultid="1328" heatid="1825" lane="6" entrytime="00:01:07.42" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="423" swimtime="00:00:59.70" resultid="1329" heatid="1800" lane="5" entrytime="00:01:01.30" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.91" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="391" swimtime="00:01:15.55" resultid="1330" heatid="1861" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriela" lastname="Poletti Veiga" birthdate="2010-10-01" gender="F" nation="BRA" license="376951" swrid="5603895" athleteid="1321" externalid="376951">
              <RESULTS>
                <RESULT eventid="1154" points="270" swimtime="00:01:23.55" resultid="1322" heatid="1823" lane="1" entrytime="00:01:19.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="433" swimtime="00:01:06.42" resultid="1323" heatid="1796" lane="2" entrytime="00:01:05.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.08" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Francisco" lastname="Silva Telles" birthdate="2011-07-19" gender="M" nation="BRA" license="377311" swrid="5603911" athleteid="1331" externalid="377311">
              <RESULTS>
                <RESULT eventid="1096" status="DSQ" swimtime="00:03:31.11" resultid="1332" heatid="1804" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.55" />
                    <SPLIT distance="100" swimtime="00:01:41.28" />
                    <SPLIT distance="150" swimtime="00:02:37.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="192" swimtime="00:01:17.69" resultid="1333" heatid="1798" lane="3" entrytime="00:01:15.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Vieira Daudt" birthdate="2008-08-14" gender="M" nation="BRA" license="350467" swrid="5603926" athleteid="1314" externalid="350467" level="VIBE">
              <RESULTS>
                <RESULT eventid="1162" points="262" swimtime="00:01:14.66" resultid="1315" heatid="1824" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.66" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="356" swimtime="00:01:03.21" resultid="1316" heatid="1797" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="285" swimtime="00:01:13.44" resultid="1317" heatid="1855" lane="5" entrytime="00:01:15.12" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.52" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Betina" lastname="Tramontini Queiroz" birthdate="2007-09-11" gender="F" nation="BRA" license="357155" swrid="5658063" athleteid="1318" externalid="357155" level="VIBE">
              <RESULTS>
                <RESULT eventid="1110" points="459" swimtime="00:10:18.75" resultid="1319" heatid="1810" lane="3" entrytime="00:09:51.57" entrycourse="SCM" />
                <RESULT eventid="1208" points="484" swimtime="00:02:20.47" resultid="1320" heatid="1840" lane="4" entrytime="00:02:22.67" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="2416" nation="BRA" region="PR" clubid="1338" swrid="93758" name="Apan/Maringá">
          <ATHLETES>
            <ATHLETE firstname="Carina" lastname="Costa Profeta" birthdate="2008-03-20" gender="F" nation="BRA" license="366964" swrid="5591584" athleteid="1377" externalid="366964">
              <RESULTS>
                <RESULT eventid="1066" points="442" swimtime="00:01:05.95" resultid="1378" heatid="1796" lane="5" entrytime="00:01:06.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="472" swimtime="00:01:20.08" resultid="1379" heatid="1860" lane="3" entrytime="00:01:17.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Marques" birthdate="2015-10-15" gender="F" nation="BRA" license="399738" swrid="5651346" athleteid="1561" externalid="399738">
              <RESULTS>
                <RESULT eventid="1302" points="26" swimtime="00:01:16.99" resultid="1562" heatid="1867" lane="1" entrytime="00:01:22.02" entrycourse="SCM" />
                <RESULT eventid="1254" points="35" swimtime="00:01:16.66" resultid="1563" heatid="1849" lane="2" entrytime="00:01:15.08" entrycourse="SCM" />
                <RESULT eventid="1276" points="21" swimtime="00:01:41.83" resultid="1564" heatid="1856" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Batista Sanchez" birthdate="2009-05-22" gender="M" nation="BRA" license="370668" swrid="5255779" athleteid="1354" externalid="370668">
              <RESULTS>
                <RESULT eventid="1118" points="336" swimtime="00:10:37.45" resultid="1355" heatid="1811" lane="3" />
                <RESULT eventid="1194" points="306" swimtime="00:05:48.08" resultid="1356" heatid="1836" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.85" />
                    <SPLIT distance="100" swimtime="00:01:20.48" />
                    <SPLIT distance="150" swimtime="00:02:09.27" />
                    <SPLIT distance="200" swimtime="00:02:53.94" />
                    <SPLIT distance="250" swimtime="00:03:39.45" />
                    <SPLIT distance="300" swimtime="00:04:26.29" />
                    <SPLIT distance="350" swimtime="00:05:07.75" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiz" lastname="Otavio Costa" birthdate="2009-01-28" gender="M" nation="BRA" license="370666" swrid="5603881" athleteid="1423" externalid="370666">
              <RESULTS>
                <RESULT eventid="1074" points="258" swimtime="00:01:10.37" resultid="1424" heatid="1797" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="272" swimtime="00:01:25.22" resultid="1425" heatid="1862" lane="6" entrytime="00:01:31.70" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.15" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Carlos" lastname="Eduardo Ebiner" birthdate="2013-07-29" gender="M" nation="BRA" license="397371" swrid="5641763" athleteid="1549" externalid="397371">
              <RESULTS>
                <RESULT eventid="1151" points="102" swimtime="00:00:53.39" resultid="1550" heatid="1821" lane="5" entrytime="00:00:56.52" entrycourse="SCM" />
                <RESULT eventid="1173" points="117" swimtime="00:01:31.58" resultid="1551" heatid="1829" lane="3" entrytime="00:01:53.15" entrycourse="SCM" />
                <RESULT eventid="1063" points="106" swimtime="00:03:50.94" resultid="1552" heatid="1793" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.18" />
                    <SPLIT distance="100" swimtime="00:01:55.22" />
                    <SPLIT distance="150" swimtime="00:02:58.53" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bernardo" lastname="Tomazeli" birthdate="2013-02-05" gender="M" nation="BRA" license="392109" swrid="5614097" athleteid="1513" externalid="392109">
              <RESULTS>
                <RESULT eventid="1107" points="104" swimtime="00:00:46.24" resultid="1514" heatid="1809" lane="5" entrytime="00:00:54.90" entrycourse="SCM" />
                <RESULT eventid="1173" points="136" swimtime="00:01:27.01" resultid="1515" heatid="1830" lane="4" entrytime="00:01:28.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.46" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="138" swimtime="00:03:31.97" resultid="1516" heatid="1794" lane="5" entrytime="00:03:40.01" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.12" />
                    <SPLIT distance="100" swimtime="00:01:42.66" />
                    <SPLIT distance="150" swimtime="00:02:44.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Furuchi Martins" birthdate="2011-10-05" gender="F" nation="BRA" license="367001" swrid="5602616" athleteid="1523" externalid="367001">
              <RESULTS>
                <RESULT eventid="1088" points="277" swimtime="00:03:26.35" resultid="1524" heatid="1803" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.56" />
                    <SPLIT distance="100" swimtime="00:01:41.35" />
                    <SPLIT distance="150" swimtime="00:02:35.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="290" swimtime="00:01:34.16" resultid="1525" heatid="1860" lane="1" entrytime="00:01:49.86" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.69" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Henrique Goes" birthdate="2008-10-26" gender="M" nation="BRA" license="392105" swrid="5603853" athleteid="1501" externalid="392105">
              <RESULTS>
                <RESULT eventid="1162" points="162" swimtime="00:01:27.63" resultid="1502" heatid="1824" lane="4" entrytime="00:01:22.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.54" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="202" swimtime="00:03:24.75" resultid="1503" heatid="1804" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.38" />
                    <SPLIT distance="100" swimtime="00:01:40.16" />
                    <SPLIT distance="150" swimtime="00:02:33.36" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="206" swimtime="00:01:33.59" resultid="1504" heatid="1861" lane="3" entrytime="00:01:37.15" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isabella" lastname="Pastre" birthdate="2014-03-10" gender="F" nation="BRA" license="403760" swrid="5684593" athleteid="1577" externalid="403760">
              <RESULTS>
                <RESULT eventid="1302" points="154" swimtime="00:00:42.70" resultid="1578" heatid="1867" lane="4" entrytime="00:00:46.81" entrycourse="SCM" />
                <RESULT eventid="1254" points="179" swimtime="00:00:44.79" resultid="1579" heatid="1849" lane="3" entrytime="00:00:48.08" entrycourse="SCM" />
                <RESULT eventid="1180" points="142" swimtime="00:01:48.08" resultid="1580" heatid="1833" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joaquim" lastname="De Correa" birthdate="2014-12-03" gender="M" nation="BRA" license="403387" swrid="5676286" athleteid="1565" externalid="403387">
              <RESULTS>
                <RESULT eventid="1305" points="96" swimtime="00:00:44.00" resultid="1566" heatid="1869" lane="5" entrytime="00:00:44.02" entrycourse="SCM" />
                <RESULT eventid="1257" points="79" swimtime="00:00:51.46" resultid="1567" heatid="1850" lane="3" />
                <RESULT eventid="1183" points="88" swimtime="00:01:50.59" resultid="1568" heatid="1835" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicolas" lastname="Baldo De França" birthdate="2014-04-21" gender="M" nation="BRA" license="393773" swrid="5507467" athleteid="1529" externalid="393773">
              <RESULTS>
                <RESULT eventid="1183" points="80" swimtime="00:01:54.15" resultid="1530" heatid="1835" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.99" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1231" points="74" swimtime="00:00:51.80" resultid="1531" heatid="1845" lane="2" entrytime="00:00:48.49" entrycourse="SCM" />
                <RESULT eventid="1279" points="70" swimtime="00:01:00.32" resultid="1532" heatid="1859" lane="2" entrytime="00:00:58.84" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Otavio Luz" birthdate="2013-07-27" gender="M" nation="BRA" license="392111" swrid="5603882" athleteid="1517" externalid="392111">
              <RESULTS>
                <RESULT eventid="1129" points="112" swimtime="00:01:39.97" resultid="1518" heatid="1814" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="147" swimtime="00:00:41.12" resultid="1519" heatid="1809" lane="2" entrytime="00:00:52.73" entrycourse="SCM" />
                <RESULT eventid="1173" points="171" swimtime="00:01:20.73" resultid="1520" heatid="1830" lane="3" entrytime="00:01:28.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.11" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Quental De Meireles" birthdate="2008-11-20" gender="M" nation="BRA" license="392103" swrid="5603898" athleteid="1494" externalid="392103">
              <RESULTS>
                <RESULT eventid="1074" points="329" swimtime="00:01:04.95" resultid="1495" heatid="1799" lane="4" entrytime="00:01:04.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.83" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="336" swimtime="00:01:19.46" resultid="1496" heatid="1862" lane="2" entrytime="00:01:20.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.19" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laura" lastname="Sanches Ghelere" birthdate="2008-08-06" gender="F" nation="BRA" license="372024" swrid="5603905" athleteid="1386" externalid="372024">
              <RESULTS>
                <RESULT eventid="1154" points="412" swimtime="00:01:12.58" resultid="1387" heatid="1823" lane="3" entrytime="00:01:12.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="395" swimtime="00:01:14.77" resultid="1388" heatid="1853" lane="1" entrytime="00:01:17.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:09.51" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Leonardo" lastname="Pauloski Murante" birthdate="1997-06-06" gender="M" nation="BRA" license="367086" swrid="5603887" athleteid="1581" externalid="367086">
              <RESULTS>
                <RESULT eventid="1074" points="253" swimtime="00:01:10.82" resultid="1582" heatid="1797" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.97" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Pacheco" birthdate="2006-12-20" gender="M" nation="BRA" license="336850" swrid="5603854" athleteid="1374" externalid="336850">
              <RESULTS>
                <RESULT eventid="1162" points="443" swimtime="00:01:02.67" resultid="1375" heatid="1825" lane="5" entrytime="00:01:02.39" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.52" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1194" points="434" swimtime="00:05:09.95" resultid="1376" heatid="1836" lane="3" entrytime="00:05:32.02" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.41" />
                    <SPLIT distance="100" swimtime="00:01:06.99" />
                    <SPLIT distance="150" swimtime="00:01:48.53" />
                    <SPLIT distance="200" swimtime="00:02:29.64" />
                    <SPLIT distance="250" swimtime="00:03:15.65" />
                    <SPLIT distance="300" swimtime="00:04:01.36" />
                    <SPLIT distance="350" swimtime="00:04:36.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Fernandes Rivadavia" birthdate="2015-11-15" gender="F" nation="BRA" license="393774" swrid="5651342" athleteid="1533" externalid="393774">
              <RESULTS>
                <RESULT eventid="1180" points="157" swimtime="00:01:44.55" resultid="1534" heatid="1833" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="106" swimtime="00:00:51.40" resultid="1535" heatid="1844" lane="3" entrytime="00:00:53.26" entrycourse="SCM" />
                <RESULT eventid="1276" points="145" swimtime="00:00:53.96" resultid="1536" heatid="1857" lane="3" entrytime="00:00:57.20" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Diogo" lastname="Sanchez" birthdate="2012-11-29" gender="M" nation="BRA" license="370658" swrid="5603906" athleteid="1412" externalid="370658">
              <RESULTS>
                <RESULT eventid="1151" points="145" swimtime="00:00:47.43" resultid="1413" heatid="1821" lane="2" entrytime="00:00:55.38" entrycourse="SCM" />
                <RESULT eventid="1173" points="113" swimtime="00:01:32.66" resultid="1414" heatid="1830" lane="1" entrytime="00:01:38.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="120" swimtime="00:03:41.74" resultid="1415" heatid="1793" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.20" />
                    <SPLIT distance="100" swimtime="00:01:49.78" />
                    <SPLIT distance="150" swimtime="00:02:49.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Henrique Campelo" birthdate="2011-09-12" gender="M" nation="BRA" license="366963" swrid="5588742" athleteid="1402" externalid="366963">
              <RESULTS>
                <RESULT eventid="1162" points="249" swimtime="00:01:15.87" resultid="1403" heatid="1824" lane="3" entrytime="00:01:14.85" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.65" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="369" swimtime="00:01:02.50" resultid="1404" heatid="1799" lane="3" entrytime="00:01:03.59" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.05" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="344" swimtime="00:02:21.69" resultid="1405" heatid="1842" lane="5" entrytime="00:02:31.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.48" />
                    <SPLIT distance="100" swimtime="00:01:07.70" />
                    <SPLIT distance="150" swimtime="00:01:45.35" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enzo" lastname="Marques Picolo Vinha" birthdate="2010-07-01" gender="M" nation="BRA" license="366990" swrid="5603869" athleteid="1526" externalid="366990">
              <RESULTS>
                <RESULT eventid="1074" points="342" swimtime="00:01:04.09" resultid="1527" heatid="1799" lane="2" entrytime="00:01:05.40" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="342" swimtime="00:02:22.00" resultid="1528" heatid="1842" lane="4" entrytime="00:02:30.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.60" />
                    <SPLIT distance="100" swimtime="00:01:09.15" />
                    <SPLIT distance="150" swimtime="00:01:47.39" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pietro" lastname="Nabas De Assis" birthdate="2011-07-09" gender="M" nation="BRA" license="366968" swrid="5603878" athleteid="1406" externalid="366968">
              <RESULTS>
                <RESULT eventid="1096" points="327" swimtime="00:02:54.37" resultid="1407" heatid="1804" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.04" />
                    <SPLIT distance="100" swimtime="00:01:23.76" />
                    <SPLIT distance="150" swimtime="00:02:09.59" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="336" swimtime="00:01:19.51" resultid="1408" heatid="1862" lane="4" entrytime="00:01:19.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nicole" lastname="De Meira" birthdate="2012-01-21" gender="F" nation="BRA" license="377257" swrid="5615583" athleteid="1426" externalid="377257">
              <RESULTS>
                <RESULT eventid="1148" points="112" swimtime="00:00:58.75" resultid="1427" heatid="1819" lane="5" />
                <RESULT eventid="1170" points="111" swimtime="00:01:44.54" resultid="1428" heatid="1827" lane="6" entrytime="00:01:48.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="122" swimtime="00:04:05.47" resultid="1429" heatid="1792" lane="6" entrytime="00:04:18.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:59.99" />
                    <SPLIT distance="100" swimtime="00:01:59.52" />
                    <SPLIT distance="150" swimtime="00:03:09.20" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Laion" lastname="Miguel Simoes" birthdate="2016-04-02" gender="M" nation="BRA" license="407179" swrid="5718695" athleteid="1591" externalid="407179">
              <RESULTS>
                <RESULT eventid="1300" points="29" swimtime="00:01:05.23" resultid="1592" heatid="1865" lane="3" />
                <RESULT eventid="1226" points="40" swimtime="00:01:12.56" resultid="1593" heatid="1843" lane="3" />
                <RESULT eventid="1252" points="32" swimtime="00:01:09.55" resultid="1594" heatid="1848" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Otavio" lastname="Sossai Altoe" birthdate="2006-09-04" gender="M" nation="BRA" license="296488" swrid="5603915" athleteid="1339" externalid="296488">
              <RESULTS>
                <RESULT eventid="1074" points="602" swimtime="00:00:53.08" resultid="1340" heatid="1800" lane="3" entrytime="00:00:52.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:25.26" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="596" swimtime="00:01:58.04" resultid="1341" heatid="1842" lane="3" entrytime="00:01:55.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.76" />
                    <SPLIT distance="100" swimtime="00:00:56.26" />
                    <SPLIT distance="150" swimtime="00:01:26.85" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Campos" birthdate="2013-02-17" gender="M" nation="BRA" license="377262" swrid="5641756" athleteid="1442" externalid="377262">
              <RESULTS>
                <RESULT eventid="1129" points="132" swimtime="00:01:34.76" resultid="1443" heatid="1814" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="157" swimtime="00:06:33.24" resultid="1444" heatid="1802" lane="5" />
                <RESULT eventid="1173" points="190" swimtime="00:01:17.95" resultid="1445" heatid="1831" lane="6" entrytime="00:01:26.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.31" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Izzo Breschiliare" birthdate="2015-09-23" gender="M" nation="BRA" license="407182" swrid="5718669" athleteid="1602" externalid="407182">
              <RESULTS>
                <RESULT eventid="1305" points="32" swimtime="00:01:03.30" resultid="1603" heatid="1868" lane="4" entrytime="00:01:00.12" entrycourse="SCM" />
                <RESULT eventid="1257" points="36" swimtime="00:01:06.57" resultid="1604" heatid="1851" lane="5" entrytime="00:01:04.74" entrycourse="SCM" />
                <RESULT eventid="1279" points="21" swimtime="00:01:29.73" resultid="1605" heatid="1858" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Pavão" birthdate="2012-04-04" gender="F" nation="BRA" license="377259" swrid="5603888" athleteid="1430" externalid="377259">
              <RESULTS>
                <RESULT eventid="1148" points="194" swimtime="00:00:48.99" resultid="1431" heatid="1819" lane="2" />
                <RESULT eventid="1082" points="192" swimtime="00:06:40.81" resultid="1432" heatid="1801" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.69" />
                    <SPLIT distance="100" swimtime="00:01:35.68" />
                    <SPLIT distance="150" swimtime="00:02:26.79" />
                    <SPLIT distance="200" swimtime="00:03:17.84" />
                    <SPLIT distance="250" swimtime="00:04:08.61" />
                    <SPLIT distance="300" swimtime="00:04:59.57" />
                    <SPLIT distance="350" swimtime="00:05:51.69" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="154" swimtime="00:00:45.40" resultid="1433" heatid="1806" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Santos Carraro" birthdate="2014-06-04" gender="M" nation="BRA" license="392097" swrid="5603908" athleteid="1480" externalid="392097">
              <RESULTS>
                <RESULT eventid="1257" points="101" swimtime="00:00:47.33" resultid="1481" heatid="1851" lane="3" entrytime="00:00:50.69" entrycourse="SCM" />
                <RESULT eventid="1183" points="108" swimtime="00:01:43.38" resultid="1482" heatid="1835" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1231" points="87" swimtime="00:00:48.92" resultid="1483" heatid="1845" lane="4" entrytime="00:00:47.47" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Kauan" lastname="Gabriel Pereira" birthdate="2014-05-14" gender="M" nation="BRA" license="407181" swrid="5718625" athleteid="1598" externalid="407181">
              <RESULTS>
                <RESULT eventid="1305" points="51" swimtime="00:00:54.02" resultid="1599" heatid="1868" lane="3" entrytime="00:00:52.03" entrycourse="SCM" />
                <RESULT eventid="1257" points="48" swimtime="00:01:00.71" resultid="1600" heatid="1851" lane="1" entrytime="00:01:05.08" entrycourse="SCM" />
                <RESULT eventid="1279" points="19" swimtime="00:01:32.58" resultid="1601" heatid="1858" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Antônio Boeing" birthdate="2004-06-04" gender="M" nation="BRA" license="317474" swrid="5184340" athleteid="1363" externalid="317474">
              <RESULTS>
                <RESULT eventid="1162" points="639" swimtime="00:00:55.47" resultid="1364" heatid="1825" lane="3" entrytime="00:00:54.21" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:26.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="522" swimtime="00:00:59.99" resultid="1365" heatid="1854" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Garcia Cavalcante" birthdate="2011-11-21" gender="M" nation="BRA" license="378200" swrid="5603840" athleteid="1360" externalid="378200">
              <RESULTS>
                <RESULT eventid="1096" points="225" swimtime="00:03:17.30" resultid="1361" heatid="1804" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.78" />
                    <SPLIT distance="100" swimtime="00:01:33.58" />
                    <SPLIT distance="150" swimtime="00:02:25.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="250" swimtime="00:01:27.65" resultid="1362" heatid="1862" lane="5" entrytime="00:01:31.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Luiza Rampasi" birthdate="2013-10-16" gender="F" nation="BRA" license="382209" swrid="5603866" athleteid="1458" externalid="382209">
              <RESULTS>
                <RESULT eventid="1148" points="134" swimtime="00:00:55.36" resultid="1459" heatid="1820" lane="6" entrytime="00:01:01.19" entrycourse="SCM" />
                <RESULT eventid="1104" points="130" swimtime="00:00:48.10" resultid="1460" heatid="1807" lane="6" entrytime="00:00:54.50" entrycourse="SCM" />
                <RESULT eventid="1170" points="173" swimtime="00:01:30.08" resultid="1461" heatid="1827" lane="2" entrytime="00:01:39.28" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mochiutti Carneiro" birthdate="2010-04-22" gender="F" nation="BRA" license="370670" swrid="5588817" athleteid="1469" externalid="370670">
              <RESULTS>
                <RESULT eventid="1154" points="391" swimtime="00:01:13.88" resultid="1470" heatid="1823" lane="4" entrytime="00:01:16.89" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.18" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="442" swimtime="00:02:24.77" resultid="1471" heatid="1840" lane="2" entrytime="00:02:24.59" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Tiago" lastname="Ficher Delmont Pais" birthdate="2010-07-15" gender="M" nation="BRA" license="338533" swrid="5588701" athleteid="1348" externalid="338533">
              <RESULTS>
                <RESULT eventid="1162" points="432" swimtime="00:01:03.16" resultid="1349" heatid="1825" lane="1" entrytime="00:01:03.74" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="409" swimtime="00:01:14.43" resultid="1350" heatid="1863" lane="6" entrytime="00:01:16.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Pedro" lastname="Antonio Pratti" birthdate="2015-10-14" gender="M" nation="BRA" license="407180" athleteid="1595" externalid="407180">
              <RESULTS>
                <RESULT eventid="1305" points="24" swimtime="00:01:09.67" resultid="1596" heatid="1868" lane="2" />
                <RESULT eventid="1257" points="21" swimtime="00:01:19.69" resultid="1597" heatid="1850" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="De Araujo" birthdate="2015-08-09" gender="F" nation="BRA" license="407185" athleteid="1606" externalid="407185">
              <RESULTS>
                <RESULT eventid="1302" points="55" swimtime="00:01:00.25" resultid="1607" heatid="1867" lane="6" />
                <RESULT eventid="1254" points="44" swimtime="00:01:11.46" resultid="1608" heatid="1849" lane="6" />
                <RESULT eventid="1276" points="61" swimtime="00:01:11.85" resultid="1609" heatid="1856" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Ayres" birthdate="2012-05-05" gender="M" nation="BRA" license="378035" swrid="5208079" athleteid="1446" externalid="378035">
              <RESULTS>
                <RESULT eventid="1129" points="270" swimtime="00:01:14.76" resultid="1447" heatid="1815" lane="3" entrytime="00:01:22.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="284" swimtime="00:05:22.54" resultid="1448" heatid="1802" lane="3" entrytime="00:05:50.54" entrycourse="SCM" />
                <RESULT eventid="1107" points="246" swimtime="00:00:34.70" resultid="1449" heatid="1809" lane="3" entrytime="00:00:33.20" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heitor" lastname="Bello Paula" birthdate="2015-06-14" gender="M" nation="BRA" license="393776" swrid="5507529" athleteid="1537" externalid="393776">
              <RESULTS>
                <RESULT eventid="1305" points="97" swimtime="00:00:43.87" resultid="1538" heatid="1869" lane="1" entrytime="00:00:45.12" entrycourse="SCM" />
                <RESULT eventid="1279" points="63" swimtime="00:01:02.70" resultid="1539" heatid="1858" lane="5" />
                <RESULT eventid="1205" points="88" swimtime="00:03:42.84" resultid="1540" heatid="1838" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.34" />
                    <SPLIT distance="100" swimtime="00:01:45.90" />
                    <SPLIT distance="150" swimtime="00:02:47.27" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Vitoria Moreira Ferreira" birthdate="2012-08-04" gender="F" nation="BRA" license="392098" swrid="5603928" athleteid="1484" externalid="392098">
              <RESULTS>
                <RESULT eventid="1126" points="126" swimtime="00:01:49.33" resultid="1485" heatid="1813" lane="4" entrytime="00:01:53.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:55.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="124" swimtime="00:01:40.74" resultid="1486" heatid="1826" lane="3" entrytime="00:02:12.81" entrycourse="SCM" />
                <RESULT eventid="1060" points="140" swimtime="00:03:54.32" resultid="1487" heatid="1791" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:58.35" />
                    <SPLIT distance="100" swimtime="00:01:56.94" />
                    <SPLIT distance="150" swimtime="00:03:02.89" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Arthur Da Silva Ortiz" birthdate="2015-04-20" gender="M" nation="BRA" license="399733" swrid="5676285" athleteid="1553" externalid="399733">
              <RESULTS>
                <RESULT eventid="1257" points="60" swimtime="00:00:56.40" resultid="1554" heatid="1850" lane="4" />
                <RESULT eventid="1183" points="81" swimtime="00:01:53.85" resultid="1555" heatid="1834" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.76" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1279" points="86" swimtime="00:00:56.39" resultid="1556" heatid="1859" lane="4" entrytime="00:00:56.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Garcia Cavalcante" birthdate="2008-08-11" gender="M" nation="BRA" license="369676" swrid="5603841" athleteid="1357" externalid="369676">
              <RESULTS>
                <RESULT eventid="1096" points="413" swimtime="00:02:41.27" resultid="1358" heatid="1805" lane="2" entrytime="00:02:45.31" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.80" />
                    <SPLIT distance="100" swimtime="00:01:16.07" />
                    <SPLIT distance="150" swimtime="00:01:57.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="413" swimtime="00:01:14.21" resultid="1359" heatid="1863" lane="5" entrytime="00:01:13.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Catarina" lastname="Wendt Jesus" birthdate="2013-07-09" gender="F" nation="BRA" license="393778" swrid="5641780" athleteid="1541" externalid="393778">
              <RESULTS>
                <RESULT eventid="1148" points="276" swimtime="00:00:43.54" resultid="1542" heatid="1820" lane="4" entrytime="00:00:45.79" entrycourse="SCM" />
                <RESULT eventid="1104" points="259" swimtime="00:00:38.23" resultid="1543" heatid="1807" lane="2" entrytime="00:00:41.93" entrycourse="SCM" />
                <RESULT eventid="1060" points="291" swimtime="00:03:03.72" resultid="1544" heatid="1792" lane="4" entrytime="00:03:17.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.79" />
                    <SPLIT distance="100" swimtime="00:01:29.88" />
                    <SPLIT distance="150" swimtime="00:02:22.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Murilo" lastname="Muniz" birthdate="2012-09-03" gender="M" nation="BRA" license="392106" swrid="5603877" athleteid="1505" externalid="392106">
              <RESULTS>
                <RESULT eventid="1129" points="82" swimtime="00:01:50.85" resultid="1506" heatid="1815" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.57" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="78" swimtime="00:00:50.79" resultid="1507" heatid="1809" lane="6" />
                <RESULT eventid="1173" points="125" swimtime="00:01:29.52" resultid="1508" heatid="1830" lane="2" entrytime="00:01:31.17" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.18" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabrielle" lastname="Borba" birthdate="2014-06-15" gender="F" nation="BRA" license="385705" swrid="5323267" athleteid="1462" externalid="385705">
              <RESULTS>
                <RESULT eventid="1302" points="139" swimtime="00:00:44.25" resultid="1463" heatid="1867" lane="3" entrytime="00:00:45.19" entrycourse="SCM" />
                <RESULT eventid="1180" points="123" swimtime="00:01:53.49" resultid="1464" heatid="1833" lane="3" entrytime="00:02:05.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:53.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1276" points="109" swimtime="00:00:59.33" resultid="1465" heatid="1857" lane="4" entrytime="00:00:57.94" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gustavo" lastname="Bessa" birthdate="2003-06-19" gender="M" nation="BRA" license="317841" swrid="5312237" athleteid="1342" externalid="317841">
              <RESULTS>
                <RESULT eventid="1096" points="563" swimtime="00:02:25.51" resultid="1343" heatid="1805" lane="3" entrytime="00:02:21.91" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.92" />
                    <SPLIT distance="100" swimtime="00:01:08.56" />
                    <SPLIT distance="150" swimtime="00:01:46.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="620" swimtime="00:01:04.80" resultid="1344" heatid="1863" lane="3" entrytime="00:01:03.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Daniela" lastname="Inoue" birthdate="2008-10-31" gender="F" nation="BRA" license="378348" swrid="5603856" athleteid="1395" externalid="378348">
              <RESULTS>
                <RESULT eventid="1066" points="364" swimtime="00:01:10.35" resultid="1396" heatid="1796" lane="6" entrytime="00:01:12.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="333" swimtime="00:02:38.99" resultid="1397" heatid="1839" lane="4" entrytime="00:02:47.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.00" />
                    <SPLIT distance="100" swimtime="00:01:15.45" />
                    <SPLIT distance="150" swimtime="00:01:58.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eduardo" lastname="Biason Santana" birthdate="2009-01-21" gender="M" nation="BRA" license="366969" swrid="5317765" athleteid="1392" externalid="366969">
              <RESULTS>
                <RESULT eventid="1074" points="403" swimtime="00:01:00.69" resultid="1393" heatid="1800" lane="2" entrytime="00:01:00.51" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.92" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="359" swimtime="00:02:30.30" resultid="1394" heatid="1846" lane="4" entrytime="00:02:32.97" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.36" />
                    <SPLIT distance="100" swimtime="00:01:10.33" />
                    <SPLIT distance="150" swimtime="00:01:49.76" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Agnes" lastname="Sophie Amadei" birthdate="2014-01-10" gender="F" nation="BRA" license="403388" swrid="5676293" athleteid="1569" externalid="403388">
              <RESULTS>
                <RESULT eventid="1302" points="91" swimtime="00:00:50.80" resultid="1570" heatid="1866" lane="2" />
                <RESULT eventid="1254" points="61" swimtime="00:01:04.08" resultid="1571" heatid="1849" lane="5" />
                <RESULT eventid="1202" points="101" swimtime="00:03:56.14" resultid="1572" heatid="1837" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:51.54" />
                    <SPLIT distance="100" swimtime="00:01:52.95" />
                    <SPLIT distance="150" swimtime="00:02:56.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Donato De Morais" birthdate="2009-03-28" gender="F" nation="BRA" license="345588" swrid="5485198" athleteid="1380" externalid="345588">
              <RESULTS>
                <RESULT eventid="1132" points="396" swimtime="00:02:41.96" resultid="1381" heatid="1816" lane="2" entrytime="00:02:44.43" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.47" />
                    <SPLIT distance="100" swimtime="00:01:18.68" />
                    <SPLIT distance="150" swimtime="00:02:00.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="373" swimtime="00:01:16.23" resultid="1382" heatid="1853" lane="5" entrytime="00:01:16.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Matheus" lastname="Junio Brambilla" birthdate="2002-04-08" gender="M" nation="BRA" license="392112" swrid="5603859" athleteid="1521" externalid="392112">
              <RESULTS>
                <RESULT eventid="1074" points="212" swimtime="00:01:15.12" resultid="1522" heatid="1797" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.01" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Danilo" lastname="Seganfredo Boscolo" birthdate="2012-09-15" gender="M" nation="BRA" license="399737" swrid="5651351" athleteid="1557" externalid="399737">
              <RESULTS>
                <RESULT eventid="1151" points="99" swimtime="00:00:53.79" resultid="1558" heatid="1821" lane="1" />
                <RESULT eventid="1107" points="49" swimtime="00:00:59.07" resultid="1559" heatid="1809" lane="1" />
                <RESULT eventid="1173" points="113" swimtime="00:01:32.62" resultid="1560" heatid="1829" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Juan" lastname="Bernardo Padua" birthdate="2013-07-15" gender="M" nation="BRA" license="392108" swrid="5305422" athleteid="1509" externalid="392108">
              <RESULTS>
                <RESULT eventid="1151" points="148" swimtime="00:00:47.13" resultid="1510" heatid="1821" lane="4" entrytime="00:00:50.60" entrycourse="SCM" />
                <RESULT eventid="1107" points="114" swimtime="00:00:44.82" resultid="1511" heatid="1808" lane="2" />
                <RESULT eventid="1173" points="175" swimtime="00:01:20.04" resultid="1512" heatid="1830" lane="5" entrytime="00:01:33.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Antonio Mendes" birthdate="2008-12-04" gender="M" nation="BRA" license="366962" swrid="5196287" athleteid="1389" externalid="366962">
              <RESULTS>
                <RESULT eventid="1096" points="472" swimtime="00:02:34.23" resultid="1390" heatid="1805" lane="5" entrytime="00:02:48.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.13" />
                    <SPLIT distance="100" swimtime="00:01:12.72" />
                    <SPLIT distance="150" swimtime="00:01:52.86" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="521" swimtime="00:01:08.68" resultid="1391" heatid="1863" lane="2" entrytime="00:01:13.04" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.22" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Manuela" lastname="Martins Pedro" birthdate="2015-01-19" gender="F" nation="BRA" license="403390" swrid="5676290" athleteid="1573" externalid="403390">
              <RESULTS>
                <RESULT eventid="1302" points="93" swimtime="00:00:50.54" resultid="1574" heatid="1866" lane="4" />
                <RESULT eventid="1180" points="52" swimtime="00:02:30.81" resultid="1575" heatid="1833" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.79" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="58" swimtime="00:01:02.78" resultid="1576" heatid="1844" lane="5" entrytime="00:01:12.55" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Yasmin" lastname="Ghelere" birthdate="2011-04-03" gender="F" nation="BRA" license="368146" swrid="5603843" athleteid="1409" externalid="368146">
              <RESULTS>
                <RESULT eventid="1066" points="326" swimtime="00:01:12.96" resultid="1410" heatid="1795" lane="3" entrytime="00:01:13.71" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="276" swimtime="00:01:24.29" resultid="1411" heatid="1852" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.50" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Camila Cuenca" birthdate="2005-10-06" gender="F" nation="BRA" license="308081" swrid="5357445" athleteid="1366" externalid="308081">
              <RESULTS>
                <RESULT eventid="1132" points="362" swimtime="00:02:46.77" resultid="1367" heatid="1816" lane="3" entrytime="00:02:36.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.08" />
                    <SPLIT distance="100" swimtime="00:01:21.92" />
                    <SPLIT distance="150" swimtime="00:02:04.35" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="413" swimtime="00:01:07.47" resultid="1368" heatid="1796" lane="3" entrytime="00:01:03.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.48" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="371" swimtime="00:01:16.35" resultid="1369" heatid="1853" lane="2" entrytime="00:01:16.14" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.41" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="425" swimtime="00:02:26.69" resultid="1370" heatid="1840" lane="3" entrytime="00:02:22.34" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Heloisa" lastname="Peroni Passafaro" birthdate="2013-09-17" gender="F" nation="BRA" license="370659" swrid="5603893" athleteid="1416" externalid="370659">
              <RESULTS>
                <RESULT eventid="1104" points="144" swimtime="00:00:46.48" resultid="1417" heatid="1806" lane="2" />
                <RESULT eventid="1170" points="186" swimtime="00:01:28.00" resultid="1418" heatid="1828" lane="4" entrytime="00:01:27.16" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="171" swimtime="00:03:39.26" resultid="1419" heatid="1792" lane="1" entrytime="00:03:52.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.78" />
                    <SPLIT distance="100" swimtime="00:01:40.76" />
                    <SPLIT distance="150" swimtime="00:02:49.71" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sarah" lastname="Chaim" birthdate="2011-05-29" gender="F" nation="BRA" license="370662" swrid="5409721" athleteid="1420" externalid="370662">
              <RESULTS>
                <RESULT eventid="1066" points="268" swimtime="00:01:17.89" resultid="1421" heatid="1795" lane="2" entrytime="00:01:19.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="204" swimtime="00:01:33.20" resultid="1422" heatid="1852" lane="3" entrytime="00:01:35.34" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.74" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Wellington" lastname="De Lima" birthdate="2008-03-01" gender="M" nation="BRA" license="370024" swrid="5470912" athleteid="1351" externalid="370024">
              <RESULTS>
                <RESULT eventid="1074" points="490" swimtime="00:00:56.86" resultid="1352" heatid="1800" lane="4" entrytime="00:00:56.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:27.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="377" swimtime="00:01:06.89" resultid="1353" heatid="1855" lane="3" entrytime="00:01:07.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.43" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Schuch Pimpao" birthdate="2010-12-31" gender="M" nation="BRA" license="355586" swrid="5588908" athleteid="1398" externalid="355586">
              <RESULTS>
                <RESULT eventid="1140" points="323" swimtime="00:02:33.84" resultid="1399" heatid="1818" lane="4" entrytime="00:02:47.23" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.56" />
                    <SPLIT distance="100" swimtime="00:01:13.76" />
                    <SPLIT distance="150" swimtime="00:01:53.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="312" swimtime="00:01:21.43" resultid="1400" heatid="1861" lane="2" />
                <RESULT eventid="1268" points="322" swimtime="00:01:10.45" resultid="1401" heatid="1855" lane="2" entrytime="00:01:13.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.62" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Isadora" lastname="Mendes Costa" birthdate="2014-04-03" gender="F" nation="BRA" license="378341" swrid="5603873" athleteid="1583" externalid="378341">
              <RESULTS>
                <RESULT eventid="1180" points="107" swimtime="00:01:58.99" resultid="1584" heatid="1833" lane="4" entrytime="00:02:08.48" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.94" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1228" points="88" swimtime="00:00:54.62" resultid="1585" heatid="1844" lane="4" entrytime="00:00:56.06" entrycourse="SCM" />
                <RESULT eventid="1276" points="102" swimtime="00:01:00.69" resultid="1586" heatid="1857" lane="2" entrytime="00:00:58.27" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Hammon" lastname="Henrique Costa" birthdate="2008-09-19" gender="M" nation="BRA" license="408703" athleteid="1613" externalid="408703">
              <RESULTS>
                <RESULT eventid="1074" points="322" swimtime="00:01:05.42" resultid="1614" heatid="1797" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lavinia" lastname="Bossoni" birthdate="2013-11-03" gender="F" nation="BRA" license="377260" swrid="5343093" athleteid="1434" externalid="377260">
              <RESULTS>
                <RESULT eventid="1126" points="134" swimtime="00:01:47.18" resultid="1435" heatid="1813" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="136" swimtime="00:01:37.62" resultid="1436" heatid="1827" lane="5" entrytime="00:01:42.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.29" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="146" swimtime="00:03:50.99" resultid="1437" heatid="1792" lane="5" entrytime="00:03:50.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.23" />
                    <SPLIT distance="100" swimtime="00:01:52.76" />
                    <SPLIT distance="150" swimtime="00:02:58.41" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Amanda" lastname="Beatriz Meira" birthdate="2012-04-11" gender="F" nation="BRA" license="392094" swrid="5305414" athleteid="1472" externalid="392094">
              <RESULTS>
                <RESULT eventid="1104" points="83" swimtime="00:00:55.71" resultid="1473" heatid="1806" lane="1" />
                <RESULT eventid="1170" points="159" swimtime="00:01:32.70" resultid="1474" heatid="1827" lane="1" entrytime="00:01:45.53" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.03" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="117" swimtime="00:04:08.78" resultid="1475" heatid="1791" lane="3" entrytime="00:04:30.80" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:54.85" />
                    <SPLIT distance="100" swimtime="00:01:55.71" />
                    <SPLIT distance="150" swimtime="00:03:12.40" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Beatriz" lastname="Passafaro" birthdate="2009-02-01" gender="F" nation="BRA" license="370673" swrid="5603885" athleteid="1383" externalid="370673">
              <RESULTS>
                <RESULT eventid="1154" points="266" swimtime="00:01:24.00" resultid="1384" heatid="1822" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.67" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="233" swimtime="00:01:29.20" resultid="1385" heatid="1852" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.21" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Gabriel" lastname="Casavechia Carraro" birthdate="2009-07-28" gender="M" nation="BRA" license="368150" swrid="5384752" athleteid="1345" externalid="368150">
              <RESULTS>
                <RESULT eventid="1162" points="485" swimtime="00:01:00.78" resultid="1346" heatid="1825" lane="4" entrytime="00:01:00.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:28.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="390" swimtime="00:01:15.62" resultid="1347" heatid="1861" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Nathan" lastname="Novak Pinho" birthdate="2012-11-14" gender="M" nation="BRA" license="378199" swrid="5603879" athleteid="1450" externalid="378199">
              <RESULTS>
                <RESULT eventid="1129" points="155" swimtime="00:01:29.83" resultid="1451" heatid="1815" lane="1" entrytime="00:01:34.95" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1085" points="197" swimtime="00:06:04.55" resultid="1452" heatid="1802" lane="4" entrytime="00:06:14.68" entrycourse="SCM" />
                <RESULT eventid="1173" points="198" swimtime="00:01:16.86" resultid="1453" heatid="1831" lane="2" entrytime="00:01:20.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.56" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Felipe Sakaguti" birthdate="2007-06-22" gender="M" nation="BRA" license="407187" swrid="5688778" athleteid="1610" externalid="407187">
              <RESULTS>
                <RESULT eventid="1074" points="69" swimtime="00:01:49.09" resultid="1611" heatid="1798" lane="6" entrytime="00:01:46.46" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.47" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="52" swimtime="00:02:09.07" resultid="1612" heatid="1854" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:57.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Bassil" birthdate="2015-07-02" gender="M" nation="BRA" license="407178" swrid="5718890" athleteid="1587" externalid="407178">
              <RESULTS>
                <RESULT eventid="1305" status="DNS" swimtime="00:00:00.00" resultid="1588" heatid="1869" lane="6" entrytime="00:00:49.14" entrycourse="SCM" />
                <RESULT eventid="1257" status="DNS" swimtime="00:00:00.00" resultid="1589" heatid="1851" lane="6" />
                <RESULT eventid="1279" status="DNS" swimtime="00:00:00.00" resultid="1590" heatid="1859" lane="5" entrytime="00:00:59.32" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Raphael" lastname="Piai Pellegrini" birthdate="2012-03-24" gender="M" nation="BRA" license="377261" swrid="5603894" athleteid="1438" externalid="377261">
              <RESULTS>
                <RESULT eventid="1129" status="DNS" swimtime="00:00:00.00" resultid="1439" heatid="1815" lane="2" entrytime="00:01:26.85" entrycourse="SCM" />
                <RESULT eventid="1085" status="DNS" swimtime="00:00:00.00" resultid="1440" heatid="1802" lane="2" />
                <RESULT eventid="1173" status="DNS" swimtime="00:00:00.00" resultid="1441" heatid="1831" lane="3" entrytime="00:01:09.19" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felype" lastname="Gongora Zago" birthdate="2011-09-14" gender="M" nation="BRA" license="392099" swrid="5603848" athleteid="1488" externalid="392099">
              <RESULTS>
                <RESULT eventid="1074" points="187" swimtime="00:01:18.34" resultid="1489" heatid="1798" lane="1" entrytime="00:01:29.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="137" swimtime="00:01:33.61" resultid="1490" heatid="1854" lane="4" entrytime="00:01:45.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.12" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Luiza" lastname="Sol Reolon Gomes" birthdate="2011-02-28" gender="F" nation="BRA" license="392100" swrid="5603914" athleteid="1491" externalid="392100">
              <RESULTS>
                <RESULT eventid="1066" points="343" swimtime="00:01:11.72" resultid="1492" heatid="1795" lane="4" entrytime="00:01:14.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="297" swimtime="00:01:22.19" resultid="1493" heatid="1853" lane="6" entrytime="00:01:32.65" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.86" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Miguel" lastname="Dos Reis Monteiro" birthdate="2014-08-05" gender="M" nation="BRA" license="392095" swrid="5697226" athleteid="1476" externalid="392095">
              <RESULTS>
                <RESULT eventid="1305" points="189" swimtime="00:00:35.10" resultid="1477" heatid="1869" lane="3" entrytime="00:00:34.32" entrycourse="SCM" />
                <RESULT eventid="1183" points="166" swimtime="00:01:29.53" resultid="1478" heatid="1834" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1231" points="152" swimtime="00:00:40.67" resultid="1479" heatid="1845" lane="3" entrytime="00:00:38.62" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Julia" lastname="Paiva Boeing" birthdate="2008-01-22" gender="F" nation="BRA" license="318185" swrid="5603884" athleteid="1371" externalid="318185">
              <RESULTS>
                <RESULT eventid="1154" points="350" swimtime="00:01:16.63" resultid="1372" heatid="1823" lane="2" entrytime="00:01:17.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="400" swimtime="00:02:29.59" resultid="1373" heatid="1839" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:32.77" />
                    <SPLIT distance="100" swimtime="00:01:09.99" />
                    <SPLIT distance="150" swimtime="00:01:50.23" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Antonio" lastname="Rafael Padial" birthdate="2014-03-07" gender="M" nation="BRA" license="397331" swrid="5641774" athleteid="1545" externalid="397331">
              <RESULTS>
                <RESULT eventid="1305" points="155" swimtime="00:00:37.46" resultid="1546" heatid="1868" lane="6" />
                <RESULT eventid="1257" points="131" swimtime="00:00:43.53" resultid="1547" heatid="1851" lane="2" entrytime="00:00:54.03" entrycourse="SCM" />
                <RESULT eventid="1183" points="117" swimtime="00:01:40.50" resultid="1548" heatid="1834" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.03" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bianca" lastname="Corsine Ferreira" birthdate="2010-03-10" gender="F" nation="BRA" license="353591" swrid="5588608" athleteid="1466" externalid="353591">
              <RESULTS>
                <RESULT eventid="1132" points="397" swimtime="00:02:41.74" resultid="1467" heatid="1816" lane="5" entrytime="00:02:46.03" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.96" />
                    <SPLIT distance="100" swimtime="00:01:18.28" />
                    <SPLIT distance="150" swimtime="00:01:59.85" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="364" swimtime="00:01:16.87" resultid="1468" heatid="1853" lane="3" entrytime="00:01:13.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.95" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Vitor" lastname="Forti Francisco" birthdate="2015-07-08" gender="M" nation="BRA" license="392104" swrid="5534395" athleteid="1497" externalid="392104">
              <RESULTS>
                <RESULT eventid="1231" points="54" swimtime="00:00:57.51" resultid="1498" heatid="1845" lane="5" entrytime="00:00:57.51" entrycourse="SCM" />
                <RESULT eventid="1279" points="83" swimtime="00:00:57.13" resultid="1499" heatid="1859" lane="6" entrytime="00:01:00.48" entrycourse="SCM" />
                <RESULT eventid="1205" points="94" swimtime="00:03:38.17" resultid="1500" heatid="1838" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.34" />
                    <SPLIT distance="100" swimtime="00:01:44.55" />
                    <SPLIT distance="150" swimtime="00:02:42.14" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lara" lastname="Constantino" birthdate="2012-06-02" gender="F" nation="BRA" license="382208" swrid="5420069" athleteid="1454" externalid="382208">
              <RESULTS>
                <RESULT eventid="1148" points="224" swimtime="00:00:46.71" resultid="1455" heatid="1820" lane="2" entrytime="00:00:46.73" entrycourse="SCM" />
                <RESULT eventid="1126" points="169" swimtime="00:01:39.20" resultid="1456" heatid="1812" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1082" points="232" swimtime="00:06:16.14" resultid="1457" heatid="1801" lane="4" entrytime="00:07:19.75" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.56" />
                    <SPLIT distance="100" swimtime="00:01:27.55" />
                    <SPLIT distance="150" swimtime="00:02:15.44" />
                    <SPLIT distance="200" swimtime="00:03:03.37" />
                    <SPLIT distance="250" swimtime="00:03:50.88" />
                    <SPLIT distance="300" swimtime="00:04:39.62" />
                    <SPLIT distance="350" swimtime="00:05:28.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
        <CLUB type="CLUB" code="16053" nation="BRA" region="PR" clubid="1615" swrid="93777" name="Fábrica De Nadadores" shortname="Fábrica">
          <ATHLETES>
            <ATHLETE firstname="Alex" lastname="Junior" birthdate="2013-03-11" gender="M" nation="BRA" license="385710" swrid="5603860" athleteid="1700" externalid="385710">
              <RESULTS>
                <RESULT eventid="1129" status="WDR" swimtime="00:00:00.00" resultid="1701" heatid="1814" lane="2" />
                <RESULT eventid="1173" status="WDR" swimtime="00:00:00.00" resultid="1702" heatid="1829" lane="4" entrytime="00:02:05.87" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Guilherme Ortega" birthdate="1999-08-05" gender="M" nation="BRA" license="383118" swrid="5603852" athleteid="1630" externalid="383118">
              <RESULTS>
                <RESULT eventid="1140" points="351" swimtime="00:02:29.61" resultid="1631" heatid="1818" lane="3" entrytime="00:02:45.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.84" />
                    <SPLIT distance="100" swimtime="00:01:11.52" />
                    <SPLIT distance="150" swimtime="00:01:51.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1118" points="301" swimtime="00:11:01.57" resultid="1632" heatid="1811" lane="4" />
                <RESULT eventid="1074" points="390" swimtime="00:01:01.37" resultid="1633" heatid="1800" lane="6" entrytime="00:01:02.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.24" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="380" swimtime="00:01:06.71" resultid="1634" heatid="1855" lane="4" entrytime="00:01:09.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.82" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Theo" lastname="Rossi" birthdate="2012-05-21" gender="M" nation="BRA" license="378346" swrid="5603901" athleteid="1658" externalid="378346">
              <RESULTS>
                <RESULT eventid="1129" points="197" swimtime="00:01:23.00" resultid="1659" heatid="1815" lane="5" entrytime="00:01:30.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1173" points="235" swimtime="00:01:12.60" resultid="1660" heatid="1831" lane="4" entrytime="00:01:16.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.15" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="200" swimtime="00:03:07.45" resultid="1661" heatid="1794" lane="2" entrytime="00:03:19.25" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.36" />
                    <SPLIT distance="100" swimtime="00:01:26.90" />
                    <SPLIT distance="150" swimtime="00:02:25.73" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Rafael" lastname="Britto" birthdate="2012-10-04" gender="M" nation="BRA" license="378350" swrid="5588566" athleteid="1666" externalid="378350">
              <RESULTS>
                <RESULT eventid="1129" points="260" swimtime="00:01:15.63" resultid="1667" heatid="1815" lane="4" entrytime="00:01:22.67" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.51" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1107" points="229" swimtime="00:00:35.52" resultid="1668" heatid="1808" lane="3" />
                <RESULT eventid="1063" points="219" swimtime="00:03:01.68" resultid="1669" heatid="1794" lane="3" entrytime="00:03:13.22" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.45" />
                    <SPLIT distance="100" swimtime="00:01:21.95" />
                    <SPLIT distance="150" swimtime="00:02:19.02" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andressa" lastname="Zamarian Gouvea" birthdate="2007-09-18" gender="F" nation="BRA" license="318503" swrid="5603929" athleteid="1616" externalid="318503">
              <RESULTS>
                <RESULT eventid="1132" points="388" swimtime="00:02:43.03" resultid="1617" heatid="1816" lane="4" entrytime="00:02:42.20" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.97" />
                    <SPLIT distance="100" swimtime="00:01:19.73" />
                    <SPLIT distance="150" swimtime="00:02:01.68" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="387" swimtime="00:01:08.94" resultid="1618" heatid="1796" lane="1" entrytime="00:01:07.32" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:19.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="362" swimtime="00:01:16.95" resultid="1619" heatid="1853" lane="4" entrytime="00:01:15.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="389" swimtime="00:02:31.01" resultid="1620" heatid="1840" lane="5" entrytime="00:02:29.36" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Dias Rezende" birthdate="2016-03-04" gender="F" nation="BRA" license="406930" swrid="5685657" athleteid="1782" externalid="406930">
              <RESULTS>
                <RESULT eventid="1298" points="30" swimtime="00:01:13.75" resultid="1783" heatid="1864" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Rezende" birthdate="2012-01-23" gender="F" nation="BRA" license="370669" swrid="5603899" athleteid="1679" externalid="370669">
              <RESULTS>
                <RESULT eventid="1148" points="173" swimtime="00:00:50.89" resultid="1680" heatid="1820" lane="1" entrytime="00:00:55.50" entrycourse="SCM" />
                <RESULT eventid="1082" points="244" swimtime="00:06:09.65" resultid="1681" heatid="1801" lane="3" entrytime="00:06:53.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.37" />
                    <SPLIT distance="100" swimtime="00:01:27.63" />
                    <SPLIT distance="150" swimtime="00:02:15.27" />
                    <SPLIT distance="200" swimtime="00:03:03.20" />
                    <SPLIT distance="250" swimtime="00:03:49.77" />
                    <SPLIT distance="300" swimtime="00:04:37.04" />
                    <SPLIT distance="350" swimtime="00:05:23.55" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="199" swimtime="00:01:25.93" resultid="1682" heatid="1826" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Bruna" lastname="Scalise Drapzichinski" birthdate="2012-03-07" gender="F" nation="BRA" license="378349" swrid="5603909" athleteid="1662" externalid="378349">
              <RESULTS>
                <RESULT eventid="1148" points="403" swimtime="00:00:38.38" resultid="1663" heatid="1820" lane="3" entrytime="00:00:39.30" entrycourse="SCM" />
                <RESULT eventid="1126" points="293" swimtime="00:01:22.57" resultid="1664" heatid="1813" lane="3" entrytime="00:01:35.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.27" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="328" swimtime="00:00:35.33" resultid="1665" heatid="1806" lane="5" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Clara" lastname="Dias Rezende" birthdate="2016-03-04" gender="F" nation="BRA" license="406929" swrid="5631410" athleteid="1779" externalid="406929">
              <RESULTS>
                <RESULT eventid="1298" points="20" swimtime="00:01:24.31" resultid="1780" heatid="1864" lane="3" />
                <RESULT eventid="1250" points="22" swimtime="00:01:29.96" resultid="1781" heatid="1847" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Monique" lastname="Istake" birthdate="2012-04-03" gender="F" nation="BRA" license="372023" swrid="5603857" athleteid="1670" externalid="372023">
              <RESULTS>
                <RESULT eventid="1104" points="298" swimtime="00:00:36.50" resultid="1671" heatid="1807" lane="3" entrytime="00:00:36.43" entrycourse="SCM" />
                <RESULT eventid="1170" points="282" swimtime="00:01:16.55" resultid="1672" heatid="1828" lane="3" entrytime="00:01:16.27" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.19" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="271" swimtime="00:03:08.24" resultid="1673" heatid="1792" lane="3" entrytime="00:03:08.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.60" />
                    <SPLIT distance="100" swimtime="00:01:28.27" />
                    <SPLIT distance="150" swimtime="00:02:22.47" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Andre" lastname="Bilemjian Leszczynski" birthdate="2011-08-06" gender="M" nation="BRA" license="406925" swrid="5587326" athleteid="1768" externalid="406925">
              <RESULTS>
                <RESULT eventid="1162" points="105" swimtime="00:01:41.13" resultid="1769" heatid="1824" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.37" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="135" swimtime="00:01:27.27" resultid="1770" heatid="1798" lane="5" entrytime="00:01:27.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.30" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="112" swimtime="00:01:54.52" resultid="1771" heatid="1861" lane="1" />
                <RESULT eventid="1216" points="157" swimtime="00:03:04.03" resultid="1772" heatid="1841" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.39" />
                    <SPLIT distance="100" swimtime="00:01:24.81" />
                    <SPLIT distance="150" swimtime="00:02:15.66" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Souza" birthdate="2013-09-11" gender="M" nation="BRA" license="382211" swrid="5603916" athleteid="1753" externalid="382211">
              <RESULTS>
                <RESULT eventid="1107" points="133" swimtime="00:00:42.52" resultid="1754" heatid="1809" lane="4" entrytime="00:00:45.96" entrycourse="SCM" />
                <RESULT eventid="1173" points="190" swimtime="00:01:17.97" resultid="1755" heatid="1831" lane="5" entrytime="00:01:22.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.39" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="148" swimtime="00:03:26.81" resultid="1756" heatid="1793" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.25" />
                    <SPLIT distance="100" swimtime="00:01:40.01" />
                    <SPLIT distance="150" swimtime="00:02:44.13" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Joao" lastname="Pedro Drapzichinski" birthdate="2015-08-21" gender="M" nation="BRA" license="391848" swrid="5603890" athleteid="1711" externalid="391848">
              <RESULTS>
                <RESULT eventid="1305" points="102" swimtime="00:00:43.03" resultid="1712" heatid="1869" lane="2" entrytime="00:00:42.94" entrycourse="SCM" />
                <RESULT eventid="1257" points="77" swimtime="00:00:51.97" resultid="1713" heatid="1851" lane="4" entrytime="00:00:53.31" entrycourse="SCM" />
                <RESULT eventid="1183" points="85" swimtime="00:01:51.82" resultid="1714" heatid="1835" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:10.49" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Fernandes Dantas" birthdate="2016-12-14" gender="M" nation="BRA" license="406932" swrid="5700463" athleteid="1784" externalid="406932">
              <RESULTS>
                <RESULT eventid="1300" points="21" swimtime="00:01:12.80" resultid="1785" heatid="1865" lane="4" />
                <RESULT eventid="1252" points="31" swimtime="00:01:10.31" resultid="1786" heatid="1848" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Gevaerd Verssutti Garcia" birthdate="2013-10-15" gender="F" nation="BRA" license="378404" swrid="5588723" athleteid="1683" externalid="378404">
              <RESULTS>
                <RESULT eventid="1148" points="153" swimtime="00:00:53.03" resultid="1684" heatid="1819" lane="1" />
                <RESULT eventid="1126" points="210" swimtime="00:01:32.21" resultid="1685" heatid="1812" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.95" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="215" swimtime="00:01:23.77" resultid="1686" heatid="1828" lane="5" entrytime="00:01:27.96" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.88" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Benicio" lastname="Garcia" birthdate="2011-09-09" gender="M" nation="BRA" license="378347" swrid="5603842" athleteid="1621" externalid="378347">
              <RESULTS>
                <RESULT eventid="1140" points="215" swimtime="00:02:56.13" resultid="1622" heatid="1818" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.35" />
                    <SPLIT distance="100" swimtime="00:01:24.93" />
                    <SPLIT distance="150" swimtime="00:02:11.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="257" swimtime="00:01:10.49" resultid="1623" heatid="1798" lane="4" entrytime="00:01:16.35" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.77" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="242" swimtime="00:01:17.55" resultid="1624" heatid="1855" lane="6" entrytime="00:01:20.44" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.93" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="237" swimtime="00:02:40.43" resultid="1625" heatid="1842" lane="6" entrytime="00:02:45.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.23" />
                    <SPLIT distance="100" swimtime="00:01:17.21" />
                    <SPLIT distance="150" swimtime="00:01:58.92" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Stephany" birthdate="2012-07-27" gender="F" nation="BRA" license="382210" swrid="5603917" athleteid="1757" externalid="382210">
              <RESULTS>
                <RESULT eventid="1104" points="140" swimtime="00:00:46.92" resultid="1758" heatid="1807" lane="1" entrytime="00:00:51.08" entrycourse="SCM" />
                <RESULT eventid="1170" points="194" swimtime="00:01:26.71" resultid="1759" heatid="1828" lane="2" entrytime="00:01:27.69" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.96" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1060" points="174" swimtime="00:03:38.27" resultid="1760" heatid="1791" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.43" />
                    <SPLIT distance="100" swimtime="00:01:42.60" />
                    <SPLIT distance="150" swimtime="00:02:52.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Valentina" lastname="Posser" birthdate="2013-02-07" gender="F" nation="BRA" license="378343" swrid="5603896" athleteid="1649" externalid="378343">
              <RESULTS>
                <RESULT eventid="1126" points="96" swimtime="00:01:59.67" resultid="1650" heatid="1813" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:56.00" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="115" swimtime="00:00:50.03" resultid="1651" heatid="1806" lane="3" entrytime="00:00:54.68" entrycourse="SCM" />
                <RESULT eventid="1170" points="116" swimtime="00:01:42.88" resultid="1652" heatid="1827" lane="4" entrytime="00:01:38.92" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:46.36" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eva" lastname="Fernandes" birthdate="2015-09-19" gender="F" nation="BRA" license="396848" swrid="5651343" athleteid="1735" externalid="396848">
              <RESULTS>
                <RESULT eventid="1302" points="94" swimtime="00:00:50.36" resultid="1736" heatid="1866" lane="3" />
                <RESULT eventid="1254" points="82" swimtime="00:00:57.99" resultid="1737" heatid="1849" lane="1" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Azevedo Martins" birthdate="2014-07-05" gender="F" nation="BRA" license="401859" swrid="5661340" athleteid="1738" externalid="401859">
              <RESULTS>
                <RESULT eventid="1302" points="68" swimtime="00:00:56.14" resultid="1739" heatid="1867" lane="5" entrytime="00:00:57.20" entrycourse="SCM" />
                <RESULT eventid="1228" points="50" swimtime="00:01:06.12" resultid="1740" heatid="1844" lane="2" entrytime="00:01:06.21" entrycourse="SCM" />
                <RESULT eventid="1276" points="86" swimtime="00:01:04.27" resultid="1741" heatid="1857" lane="5" entrytime="00:01:03.64" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Traci Rodrigues" birthdate="2014-10-27" gender="M" nation="BRA" license="406926" athleteid="1773" externalid="406926">
              <RESULTS>
                <RESULT eventid="1305" points="65" swimtime="00:00:50.03" resultid="1774" heatid="1868" lane="1" />
                <RESULT eventid="1279" points="80" swimtime="00:00:57.84" resultid="1775" heatid="1858" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caio" lastname="Braga" birthdate="2010-05-07" gender="M" nation="BRA" license="378345" swrid="5343953" athleteid="1653" externalid="378345">
              <RESULTS>
                <RESULT eventid="1096" points="360" swimtime="00:02:48.88" resultid="1654" heatid="1805" lane="6" entrytime="00:03:06.58" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.01" />
                    <SPLIT distance="100" swimtime="00:01:20.74" />
                    <SPLIT distance="150" swimtime="00:02:04.64" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" status="DNS" swimtime="00:00:00.00" resultid="1655" heatid="1799" lane="5" entrytime="00:01:06.54" entrycourse="SCM" />
                <RESULT eventid="1290" points="384" swimtime="00:01:16.02" resultid="1656" heatid="1863" lane="1" entrytime="00:01:15.11" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.61" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" status="DNS" swimtime="00:00:00.00" resultid="1657" heatid="1841" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lorenzo" lastname="Jacobsen Donati" birthdate="2011-07-14" gender="M" nation="BRA" license="391851" swrid="5615735" athleteid="1715" externalid="391851">
              <RESULTS>
                <RESULT eventid="1140" points="267" swimtime="00:02:43.95" resultid="1716" heatid="1817" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.87" />
                    <SPLIT distance="100" swimtime="00:01:18.38" />
                    <SPLIT distance="150" swimtime="00:02:02.34" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="354" swimtime="00:01:03.33" resultid="1717" heatid="1799" lane="1" entrytime="00:01:06.76" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.98" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="283" swimtime="00:01:13.54" resultid="1718" heatid="1854" lane="3" entrytime="00:01:24.87" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.08" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="305" swimtime="00:02:27.59" resultid="1719" heatid="1842" lane="1" entrytime="00:02:32.60" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.23" />
                    <SPLIT distance="100" swimtime="00:01:12.26" />
                    <SPLIT distance="150" swimtime="00:01:51.17" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sophia" lastname="Schmeiske Ruivo" birthdate="2013-10-21" gender="F" nation="BRA" license="402006" swrid="5661354" athleteid="1742" externalid="402006">
              <RESULTS>
                <RESULT eventid="1148" points="189" swimtime="00:00:49.38" resultid="1743" heatid="1819" lane="3" entrytime="00:01:01.67" entrycourse="SCM" />
                <RESULT eventid="1170" points="200" swimtime="00:01:25.91" resultid="1744" heatid="1826" lane="4" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Eduarda Guinoza" birthdate="2013-01-06" gender="F" nation="BRA" license="392012" swrid="5510698" athleteid="1720" externalid="392012">
              <RESULTS>
                <RESULT eventid="1148" points="175" swimtime="00:00:50.72" resultid="1721" heatid="1820" lane="5" entrytime="00:00:54.86" entrycourse="SCM" />
                <RESULT eventid="1126" points="119" swimtime="00:01:51.30" resultid="1722" heatid="1813" lane="6">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:52.80" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="152" swimtime="00:01:34.15" resultid="1723" heatid="1827" lane="3" entrytime="00:01:38.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.80" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Helena" lastname="Magalhães Rezende" birthdate="2010-05-29" gender="F" nation="BRA" license="366960" swrid="5588793" athleteid="1635" externalid="366960">
              <RESULTS>
                <RESULT eventid="1088" points="332" swimtime="00:03:14.27" resultid="1636" heatid="1803" lane="3" entrytime="00:03:17.29" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:43.36" />
                    <SPLIT distance="100" swimtime="00:01:31.77" />
                    <SPLIT distance="150" swimtime="00:02:22.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1110" points="309" swimtime="00:11:46.02" resultid="1637" heatid="1810" lane="4" />
                <RESULT eventid="1282" points="314" swimtime="00:01:31.73" resultid="1638" heatid="1860" lane="2" entrytime="00:01:27.93" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.13" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1208" points="344" swimtime="00:02:37.29" resultid="1639" heatid="1839" lane="3" entrytime="00:02:34.19" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:34.78" />
                    <SPLIT distance="100" swimtime="00:01:13.69" />
                    <SPLIT distance="150" swimtime="00:01:54.99" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Davi" lastname="Silverio Duarte" birthdate="2011-08-08" gender="M" nation="BRA" license="392138" swrid="5603913" athleteid="1724" externalid="392138">
              <RESULTS>
                <RESULT eventid="1140" status="WDR" swimtime="00:00:00.00" resultid="1725" heatid="1817" lane="3" />
                <RESULT eventid="1074" status="WDR" swimtime="00:00:00.00" resultid="1726" heatid="1797" lane="3" entrytime="00:01:49.84" entrycourse="SCM" />
                <RESULT eventid="1268" status="WDR" swimtime="00:00:00.00" resultid="1727" heatid="1854" lane="5" />
                <RESULT eventid="1216" status="WDR" swimtime="00:00:00.00" resultid="1728" heatid="1841" lane="2" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Caua" lastname="Pazinato" birthdate="2011-01-05" gender="M" nation="BRA" license="368149" swrid="5603889" athleteid="1674" externalid="368149">
              <RESULTS>
                <RESULT eventid="1140" points="225" swimtime="00:02:53.60" resultid="1675" heatid="1817" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.25" />
                    <SPLIT distance="100" swimtime="00:01:24.16" />
                    <SPLIT distance="150" swimtime="00:02:09.81" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="311" swimtime="00:01:06.14" resultid="1676" heatid="1799" lane="6" entrytime="00:01:08.33" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:31.53" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1268" points="229" swimtime="00:01:18.99" resultid="1677" heatid="1855" lane="1" entrytime="00:01:18.84" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:38.38" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="289" swimtime="00:02:30.27" resultid="1678" heatid="1842" lane="2" entrytime="00:02:31.08" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:35.04" />
                    <SPLIT distance="100" swimtime="00:01:13.87" />
                    <SPLIT distance="150" swimtime="00:01:53.33" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eloah" lastname="Juvedi Trindade" birthdate="2011-03-05" gender="F" nation="BRA" license="396829" swrid="5641768" athleteid="1729" externalid="396829">
              <RESULTS>
                <RESULT eventid="1088" points="232" swimtime="00:03:38.80" resultid="1730" heatid="1803" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.64" />
                    <SPLIT distance="100" swimtime="00:01:45.57" />
                    <SPLIT distance="150" swimtime="00:02:43.42" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1154" points="115" swimtime="00:01:50.84" resultid="1731" heatid="1822" lane="3" entrytime="00:02:01.15" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:50.02" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1066" points="225" swimtime="00:01:22.52" resultid="1732" heatid="1795" lane="5" entrytime="00:01:28.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.49" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1282" points="213" swimtime="00:01:44.37" resultid="1733" heatid="1860" lane="5" entrytime="00:01:46.73" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.74" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1260" points="196" swimtime="00:01:34.48" resultid="1734" heatid="1852" lane="4" entrytime="00:01:36.68" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.64" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Alice" lastname="Tiemi Yamaguchi" birthdate="2013-02-28" gender="F" nation="BRA" license="385707" swrid="5603920" athleteid="1687" externalid="385707">
              <RESULTS>
                <RESULT eventid="1126" points="213" swimtime="00:01:31.90" resultid="1688" heatid="1812" lane="3">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:45.97" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="251" swimtime="00:00:38.63" resultid="1689" heatid="1807" lane="4" entrytime="00:00:41.20" entrycourse="SCM" />
                <RESULT eventid="1060" points="264" swimtime="00:03:09.74" resultid="1690" heatid="1792" lane="2" entrytime="00:03:25.38" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.28" />
                    <SPLIT distance="100" swimtime="00:01:29.85" />
                    <SPLIT distance="150" swimtime="00:02:22.72" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Enrico" lastname="Santin Rezende" birthdate="2016-02-15" gender="M" nation="BRA" license="407196" swrid="5718892" athleteid="1787" externalid="407196">
              <RESULTS>
                <RESULT eventid="1252" status="WDR" swimtime="00:00:00.00" resultid="1788" heatid="1848" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Berto" birthdate="2008-10-22" gender="M" nation="BRA" license="378342" swrid="5312223" athleteid="1640" externalid="378342">
              <RESULTS>
                <RESULT eventid="1140" status="DSQ" swimtime="00:03:04.72" resultid="1641" heatid="1818" lane="5">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:41.70" />
                    <SPLIT distance="100" swimtime="00:01:29.01" />
                    <SPLIT distance="150" swimtime="00:02:16.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1096" points="366" swimtime="00:02:47.96" resultid="1642" heatid="1805" lane="1" entrytime="00:03:03.63" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.55" />
                    <SPLIT distance="100" swimtime="00:01:18.17" />
                    <SPLIT distance="150" swimtime="00:02:02.12" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="345" swimtime="00:01:18.81" resultid="1643" heatid="1862" lane="3" entrytime="00:01:17.98" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:37.23" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1216" points="278" swimtime="00:02:32.10" resultid="1644" heatid="1841" lane="4">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.74" />
                    <SPLIT distance="100" swimtime="00:01:13.52" />
                    <SPLIT distance="150" swimtime="00:01:52.24" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Robsson" lastname="Tows Oliveira" birthdate="2014-03-05" gender="M" nation="BRA" license="392107" swrid="5603922" athleteid="1745" externalid="392107">
              <RESULTS>
                <RESULT eventid="1305" points="110" swimtime="00:00:41.98" resultid="1746" heatid="1869" lane="4" entrytime="00:00:38.87" entrycourse="SCM" />
                <RESULT eventid="1183" points="117" swimtime="00:01:40.61" resultid="1747" heatid="1835" lane="3" entrytime="00:01:43.62" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.20" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1279" points="115" swimtime="00:00:51.16" resultid="1748" heatid="1859" lane="3" entrytime="00:00:49.66" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Eric" lastname="Moreschi" birthdate="2012-08-09" gender="M" nation="BRA" license="385715" swrid="5603876" athleteid="1703" externalid="385715">
              <RESULTS>
                <RESULT eventid="1151" points="185" swimtime="00:00:43.76" resultid="1704" heatid="1821" lane="3" entrytime="00:00:43.57" entrycourse="SCM" />
                <RESULT eventid="1173" points="205" swimtime="00:01:16.04" resultid="1705" heatid="1831" lane="1" entrytime="00:01:25.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.73" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1063" points="208" swimtime="00:03:04.88" resultid="1706" heatid="1794" lane="4" entrytime="00:03:13.83" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.12" />
                    <SPLIT distance="100" swimtime="00:01:31.04" />
                    <SPLIT distance="150" swimtime="00:02:23.44" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Dante" lastname="Gabriel Rossi" birthdate="2016-01-19" gender="M" nation="BRA" license="406928" swrid="5718627" athleteid="1776" externalid="406928">
              <RESULTS>
                <RESULT eventid="1300" points="40" swimtime="00:00:58.50" resultid="1777" heatid="1865" lane="2" />
                <RESULT eventid="1178" points="34" swimtime="00:01:06.92" resultid="1778" heatid="1832" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Arthur" lastname="Bilemjian Leszczynski" birthdate="2014-02-22" gender="M" nation="BRA" license="406924" swrid="5631285" athleteid="1764" externalid="406924">
              <RESULTS>
                <RESULT eventid="1305" points="73" swimtime="00:00:48.21" resultid="1765" heatid="1868" lane="5" />
                <RESULT eventid="1279" points="61" swimtime="00:01:03.31" resultid="1766" heatid="1859" lane="1" entrytime="00:00:59.86" entrycourse="SCM" />
                <RESULT eventid="1205" points="87" swimtime="00:03:44.03" resultid="1767" heatid="1838" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:47.61" />
                    <SPLIT distance="100" swimtime="00:01:47.03" />
                    <SPLIT distance="150" swimtime="00:02:46.46" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Sofia" lastname="Ognibeni Paupitz" birthdate="2014-08-08" gender="F" nation="BRA" license="406923" swrid="5718889" athleteid="1761" externalid="406923">
              <RESULTS>
                <RESULT eventid="1302" status="DNS" swimtime="00:00:00.00" resultid="1762" heatid="1867" lane="2" entrytime="00:00:47.38" entrycourse="SCM" />
                <RESULT eventid="1276" status="DNS" swimtime="00:00:00.00" resultid="1763" heatid="1857" lane="1" entrytime="00:01:04.07" entrycourse="SCM" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Felipe" lastname="Lima Coelho" birthdate="2012-12-12" gender="M" nation="BRA" license="393775" swrid="5615959" athleteid="1749" externalid="393775">
              <RESULTS>
                <RESULT eventid="1085" points="138" swimtime="00:06:50.29" resultid="1750" heatid="1802" lane="1" />
                <RESULT eventid="1107" status="DSQ" swimtime="00:00:45.18" resultid="1751" heatid="1808" lane="4" />
                <RESULT eventid="1173" points="141" swimtime="00:01:26.02" resultid="1752" heatid="1830" lane="6" entrytime="00:01:42.00" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.93" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Victor" lastname="Kenji Yamaguchi" birthdate="2011-08-25" gender="M" nation="BRA" license="385708" swrid="5603862" athleteid="1691" externalid="385708">
              <RESULTS>
                <RESULT eventid="1162" points="217" swimtime="00:01:19.45" resultid="1692" heatid="1824" lane="2" entrytime="00:01:25.55" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:36.60" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="245" swimtime="00:01:11.61" resultid="1693" heatid="1798" lane="2" entrytime="00:01:22.36" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:33.63" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1290" points="221" swimtime="00:01:31.42" resultid="1694" heatid="1862" lane="1" entrytime="00:01:31.56" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:44.06" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="194" swimtime="00:03:04.53" resultid="1695" heatid="1846" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:39.08" />
                    <SPLIT distance="100" swimtime="00:01:26.22" />
                    <SPLIT distance="150" swimtime="00:02:15.07" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Giovana" lastname="Jupi Takaki" birthdate="2013-03-26" gender="F" nation="BRA" license="391845" swrid="5603861" athleteid="1707" externalid="391845">
              <RESULTS>
                <RESULT eventid="1082" points="222" swimtime="00:06:21.53" resultid="1708" heatid="1801" lane="2">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.46" />
                    <SPLIT distance="100" swimtime="00:01:28.76" />
                    <SPLIT distance="150" swimtime="00:02:17.38" />
                    <SPLIT distance="200" swimtime="00:03:05.80" />
                    <SPLIT distance="250" swimtime="00:03:54.00" />
                    <SPLIT distance="300" swimtime="00:04:43.15" />
                    <SPLIT distance="350" swimtime="00:05:32.89" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1104" points="207" swimtime="00:00:41.17" resultid="1709" heatid="1807" lane="5" entrytime="00:00:47.68" entrycourse="SCM" />
                <RESULT eventid="1170" points="207" swimtime="00:01:24.87" resultid="1710" heatid="1828" lane="1" entrytime="00:01:35.90" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:40.28" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Lucas" lastname="Silveira De Almeida" birthdate="2008-07-08" gender="M" nation="BRA" license="368152" swrid="5603912" athleteid="1645" externalid="368152">
              <RESULTS>
                <RESULT eventid="1162" points="441" swimtime="00:01:02.76" resultid="1646" heatid="1825" lane="2" entrytime="00:01:01.06" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.21" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1074" points="388" swimtime="00:01:01.44" resultid="1647" heatid="1800" lane="1" entrytime="00:01:02.05" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:29.09" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1242" points="459" swimtime="00:02:18.46" resultid="1648" heatid="1846" lane="3" entrytime="00:02:26.07" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:30.80" />
                    <SPLIT distance="100" swimtime="00:01:05.98" />
                    <SPLIT distance="150" swimtime="00:01:41.65" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Maria" lastname="Valentina Gozaga" birthdate="2014-06-28" gender="F" nation="BRA" license="385709" swrid="5603924" athleteid="1696" externalid="385709">
              <RESULTS>
                <RESULT eventid="1254" points="150" swimtime="00:00:47.42" resultid="1697" heatid="1849" lane="4" entrytime="00:00:49.59" entrycourse="SCM" />
                <RESULT eventid="1180" points="151" swimtime="00:01:45.93" resultid="1698" heatid="1833" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:49.70" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1276" points="105" swimtime="00:00:59.95" resultid="1699" heatid="1856" lane="3" />
              </RESULTS>
            </ATHLETE>
            <ATHLETE firstname="Izabel" lastname="Rezende" birthdate="2013-12-13" gender="F" nation="BRA" license="370657" swrid="5603900" athleteid="1626" externalid="370657">
              <RESULTS>
                <RESULT eventid="1148" points="152" swimtime="00:00:53.10" resultid="1627" heatid="1819" lane="4" entrytime="00:01:01.94" entrycourse="SCM" />
                <RESULT eventid="1126" points="165" swimtime="00:01:40.01" resultid="1628" heatid="1813" lane="1">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:48.04" />
                  </SPLITS>
                </RESULT>
                <RESULT eventid="1170" points="185" swimtime="00:01:28.11" resultid="1629" heatid="1828" lane="6" entrytime="00:01:37.52" entrycourse="SCM">
                  <SPLITS>
                    <SPLIT distance="50" swimtime="00:00:42.00" />
                  </SPLITS>
                </RESULT>
              </RESULTS>
            </ATHLETE>
          </ATHLETES>
        </CLUB>
      </CLUBS>
    </MEET>
  </MEETS>
</LENEX>
